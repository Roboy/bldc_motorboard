// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Sep 18 21:05:11 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    inout PIN_1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    inout PIN_2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    input PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    input PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    input PIN_12 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    input PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    input PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    input PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire GND_net, VCC_net, LED_c, tx_o, tx2_o, tx_enable, tx2_enable, 
        rx_i;
    wire [25:0]blink_counter;   // verilog/TinyFPGA_B.v(64[14:27])
    
    wire n8191;
    wire [31:0]rand_data;   // verilog/TinyFPGA_B.v(77[14:23])
    wire [31:0]rand_setpoint;   // verilog/TinyFPGA_B.v(78[14:27])
    wire [7:0]byte_transmit_counter;   // coms.v(19[11:32])
    
    wire n63;
    wire [7:0]\data_out[10] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[9] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[8] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[5] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[3] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[2] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[1] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[0] ;   // coms.v(21[11:19])
    wire [7:0]\UART_TRANSMITTER.state ;   // coms.v(277[13:18])
    
    wire rx_data_ready;
    wire [7:0]rx_data;   // coms.v(374[13:20])
    wire [7:0]\data_in[3] ;   // coms.v(378[12:19])
    wire [7:0]\data_in[2] ;   // coms.v(378[12:19])
    wire [7:0]\data_in[1] ;   // coms.v(378[12:19])
    wire [7:0]\data_in[0] ;   // coms.v(378[12:19])
    wire [7:0]\data_in_frame[6] ;   // coms.v(379[12:25])
    wire [7:0]\data_out_frame2[18] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[17] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[16] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[15] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[14] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[13] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[12] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[11] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[10] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[9] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[8] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[7] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[6] ;   // coms.v(380[12:27])
    wire [7:0]\data_out_frame2[5] ;   // coms.v(380[12:27])
    
    wire tx2_active;
    wire [31:0]\FRAME_MATCHER.state ;   // coms.v(409[11:16])
    wire [7:0]tx_transmit_N_1947;
    
    wire n5266, n5244, n4, n17349, n17327, n17090, data_out_9__2__N_367, 
        n6, n17664, n18073, n18070, data_out_10__7__N_110, n160, 
        n159, n158, n157, n156, n155, n154, n153, n2699, n110, 
        n11260, n11259, n11258, n11257, n11256, n11255, n11254, 
        n11253, n11252, n11251, n11250, n11249, n11248, n11247, 
        n11246, n11245, n11244, n11243, n11242, n11241, n11240, 
        n152, n151, n150, n149, n148, n147, n146, n145, n11239, 
        n11238, n18, n11237, n9999, n11236, n11235, n11234, n11233, 
        n11232, n11231, n11230, n11229, n11228;
    wire [31:0]\FRAME_MATCHER.state_31__N_1406 ;
    
    wire n11227, n11226, n10596, n8, n2061, n11225, n11224, n10, 
        n13116, n16902, n17361, n16056, n16055, n16054, n16053, 
        n16052, n16051, n16050, n16049, n16048, n16006, n16047, 
        n18287, n16046, n16005, n5, n9, n44, n16045, n16004, 
        n16044, n16043, n16003, n16042, n16002, n16001, n5_adj_2407, 
        n16041, n16040, n16000, n16039, n16038, n15999, n16037, 
        n15998, n15994, n16036, n16035, n15997, n16034, n15996, 
        n10_adj_2408, n10_adj_2409, n6_adj_2410, n18286, n10914, n10913, 
        n11223, n11222, n10_adj_2411, n16033, n11221, n11220, n11219, 
        n11218, n11217, n10912, n11216, n16032, n10911, n11215, 
        n11214, n11213, n16031, n8_adj_2412, n11212, n16030, n11211, 
        n11210, n17412, n11209, n13744, n11208, n16029, n11207, 
        n11206, n11205, n11204, n16028, n11203, n10_adj_2413, n16027, 
        n11202, n18271, n11201, n16026, n31, n28, n11200, n11199, 
        n11198, n11197, n11196, n11195, n11194, n11193, n11192, 
        n11191, n11190, n10907, n16025, n16024, n11189, n11188, 
        n11187, n4_adj_2414, n11186, n22, n10906, n11185, n11184, 
        n10905, n11183, n11182, n10904, n31_adj_2415, n11181, n16023, 
        n4_adj_2416, n16022, n11180, n11179, n16021, n11178, n16020, 
        n10902, n11177, n15993, n15987, n16019, n11176, n11175, 
        n11174, n165, n11173, n16018, n15992, n15986, n2594, n11172, 
        n16017, n15991, n10901, n11171, n16016, n11170, n11169, 
        n16015, n16014, n11168, n16065, n16013, n11167, n11166, 
        n16064, n11165, n16012, n15990, n15985, n15983, n15982, 
        n4_adj_2417, n15980, n15979, n11164, n11163, n11162, n11161, 
        n16011, n11160, n11159, n164, n16063, n16010, n15989, 
        n11158, n15984, n15981, n15988, n63_adj_2418, n11157, n25, 
        n10900, n11156, n3779, n11155, n11154, n16062, n11153, 
        n16061, n11152, n32, n29, n11151, n4_adj_2419, n11150, 
        n11149, n23, n17, n16, n15, n14, n13, n12, n11, n10_adj_2420, 
        n9_adj_2421, n16009, n16008, n163, n18223, n10_adj_2422, 
        n26, n16060, n10899, n16924, n10898, n26_adj_2423, n25_adj_2424, 
        n24, n23_adj_2425, n22_adj_2426, n10897, n4_adj_2427, n10088, 
        n488, n63_adj_2428, n162, n7, n6_adj_2429, n10895, n4408, 
        n450, n444, \FRAME_MATCHER.i_31__N_1272 , \FRAME_MATCHER.i_31__N_1273 , 
        \FRAME_MATCHER.i_31__N_1275 , n11139, n11136, n11135, n11132, 
        n11131, n11130, n11129, n11128, n11127, n11126, n11125, 
        n11124, n11123, n11121, n11120, n11119, n11118, n11117, 
        n11116, n11115, n11114, n11113, n11112, n11111, n11110, 
        n11109, n11108, n11107, n11106, n11105, n11104, n11103, 
        n11102, n11101, n11100, n11099, n11098, n11097, n11096, 
        n11095, n11094, n11093, n11092, n11091, n11090, n11089, 
        n16620, n16618, n11039, n11038, n11037, n11034, n11033, 
        n11032, n11031, n144, n143, n142, n141, n140, n139, 
        n138, n137, n136, n135, n134, n9257, n11028, n11027, 
        n11026, n11025, n11024, n11023, n16912, n10_adj_2430, n18199, 
        n11019, n11018, n11016, n18196, n10_adj_2431, n10_adj_2432, 
        n18187, n135_adj_2433, n134_adj_2434, n133, n132, n131, 
        n130, n129, n16622, n16624, n16626, n17427, n16628, n16914, 
        n161, n16059, n18175, n16058, n10996, n10994, n17416, 
        n17765;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n16057, n16926, n128, n127, n126, n125, n124, n123, 
        n122, n121, n120, n10987, n10983, r_Rx_Data;
    wire [2:0]r_Bit_Index_adj_2499;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_adj_2500;   // verilog/uart_rx.v(36[17:26])
    
    wire n16630, n13_adj_2437, n10725, n10977, n10976, n119, n118, 
        n117, n116, n115, n114, n113, n112, n10974, n10972, 
        n10971, n18169, n10969, n10968, n10966;
    wire [2:0]r_SM_Main_adj_2503;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_2505;   // verilog/uart_tx.v(33[16:27])
    
    wire n10965;
    wire [2:0]r_SM_Main_2__N_2031_adj_2510;
    
    wire n17759, n10963, n10962, n10960, n111, n5142, n10959, 
        n10957, n10956, n10954, n10953, n10951, n10705, n16928, 
        n17089, n10_adj_2443, n16930, n16932, n16614, n16007, n10674, 
        n16632, n3, n16634, n10_adj_2444, n1, n8_adj_2445, n6_adj_2446, 
        n2, n8_adj_2447, n18280, n5_adj_2448, n1_adj_2449, n10_adj_2450, 
        n15995, n21, n20, n10923, n19, n18091, n134_adj_2451, 
        n135_adj_2452, n136_adj_2453, n137_adj_2454, n138_adj_2455, 
        n139_adj_2456, n140_adj_2457, n141_adj_2458, n142_adj_2459, 
        n143_adj_2460, n144_adj_2461, n145_adj_2462, n146_adj_2463, 
        n147_adj_2464, n148_adj_2465, n149_adj_2466, n150_adj_2467, 
        n151_adj_2468, n152_adj_2469, n153_adj_2470, n154_adj_2471, 
        n155_adj_2472, n156_adj_2473, n157_adj_2474, n158_adj_2475, 
        n159_adj_2476, n160_adj_2477, n161_adj_2478, n162_adj_2479, 
        n163_adj_2480, n164_adj_2481, n165_adj_2482, n17428, n10_adj_2483, 
        n17075, n17086, n17708, n10140, n17707, n17392, n10010, 
        n4_adj_2484, n3_adj_2485, n1_adj_2486, n21_adj_2487, n17063, 
        n13692, n9524, n6_adj_2488, n16662, n10920, n9378;
    
    VCC i2 (.Y(VCC_net));
    SB_IO tx2_output (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx2_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx2_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx2_output.PIN_TYPE = 6'b101001;
    defparam tx2_output.PULLUP = 1'b1;
    defparam tx2_output.NEG_TRIGGER = 1'b0;
    defparam tx2_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO rx_input (.PACKAGE_PIN(PIN_2), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net), .D_IN_0(rx_i)) /* synthesis lattice_noprune=1, syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam rx_input.PIN_TYPE = 6'b000001;
    defparam rx_input.PULLUP = 1'b1;
    defparam rx_input.NEG_TRIGGER = 1'b0;
    defparam rx_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_1), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i8566_3_lut (.I0(\data_out_frame2[17] [7]), .I1(rand_data[15]), 
            .I2(n10725), .I3(GND_net), .O(n11252));   // coms.v(416[12] 543[6])
    defparam i8566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8567_3_lut (.I0(\data_out_frame2[18] [0]), .I1(rand_data[0]), 
            .I2(n10725), .I3(GND_net), .O(n11253));   // coms.v(416[12] 543[6])
    defparam i8567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8568_3_lut (.I0(\data_out_frame2[18] [1]), .I1(rand_data[1]), 
            .I2(n10725), .I3(GND_net), .O(n11254));   // coms.v(416[12] 543[6])
    defparam i8568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8569_3_lut (.I0(\data_out_frame2[18] [2]), .I1(rand_data[2]), 
            .I2(n10725), .I3(GND_net), .O(n11255));   // coms.v(416[12] 543[6])
    defparam i8569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8570_3_lut (.I0(\data_out_frame2[18] [3]), .I1(rand_data[3]), 
            .I2(n10725), .I3(GND_net), .O(n11256));   // coms.v(416[12] 543[6])
    defparam i8570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8571_3_lut (.I0(\data_out_frame2[18] [4]), .I1(rand_data[4]), 
            .I2(n10725), .I3(GND_net), .O(n11257));   // coms.v(416[12] 543[6])
    defparam i8571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8572_3_lut (.I0(\data_out_frame2[18] [5]), .I1(rand_data[5]), 
            .I2(n10725), .I3(GND_net), .O(n11258));   // coms.v(416[12] 543[6])
    defparam i8572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8573_3_lut (.I0(\data_out_frame2[18] [6]), .I1(rand_data[6]), 
            .I2(n10725), .I3(GND_net), .O(n11259));   // coms.v(416[12] 543[6])
    defparam i8573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8574_3_lut (.I0(\data_out_frame2[18] [7]), .I1(rand_data[7]), 
            .I2(n10725), .I3(GND_net), .O(n11260));   // coms.v(416[12] 543[6])
    defparam i8574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8345_4_lut (.I0(n11018), .I1(r_Bit_Index_adj_2499[1]), .I2(r_Bit_Index_adj_2499[0]), 
            .I3(n17361), .O(n11031));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8345_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main_adj_2503[1]), .I1(r_SM_Main_2__N_2031_adj_2510[1]), 
            .I2(r_SM_Main_adj_2503[0]), .I3(r_SM_Main_adj_2503[2]), .O(n18280));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i8333_4_lut (.I0(n11018), .I1(r_Bit_Index_adj_2499[2]), .I2(n5244), 
            .I3(n17361), .O(n11019));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8333_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 i23_4_lut (.I0(byte_transmit_counter[1]), .I1(tx_transmit_N_1947[1]), 
            .I2(n10705), .I3(n10_adj_2444), .O(n16620));   // coms.v(280[12] 370[6])
    defparam i23_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i23_4_lut_adj_769 (.I0(byte_transmit_counter[2]), .I1(tx_transmit_N_1947[2]), 
            .I2(n10705), .I3(n10_adj_2444), .O(n16622));   // coms.v(280[12] 370[6])
    defparam i23_4_lut_adj_769.LUT_INIT = 16'hca0a;
    SB_LUT4 i23_4_lut_adj_770 (.I0(byte_transmit_counter[3]), .I1(tx_transmit_N_1947[3]), 
            .I2(n10705), .I3(n10_adj_2444), .O(n16624));   // coms.v(280[12] 370[6])
    defparam i23_4_lut_adj_770.LUT_INIT = 16'hca0a;
    SB_LUT4 i23_4_lut_adj_771 (.I0(byte_transmit_counter[4]), .I1(tx_transmit_N_1947[4]), 
            .I2(n10705), .I3(n10_adj_2444), .O(n16626));   // coms.v(280[12] 370[6])
    defparam i23_4_lut_adj_771.LUT_INIT = 16'hca0a;
    SB_LUT4 i8310_2_lut (.I0(n5142), .I1(n10994), .I2(GND_net), .I3(GND_net), 
            .O(n10996));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8310_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i24_4_lut (.I0(n18223), .I1(n10_adj_2413), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut_adj_772 (.I0(r_Tx_Data[7]), .I1(n10), .I2(n9257), 
            .I3(byte_transmit_counter[4]), .O(n16902));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i23_4_lut_adj_772.LUT_INIT = 16'h0aca;
    SB_DFF rand_data_2358__i0 (.Q(rand_data[0]), .C(CLK_c), .D(n165_adj_2482));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i53_4_lut (.I0(\data_out[0] [0]), .I1(n2), .I2(byte_transmit_counter[1]), 
            .I3(byte_transmit_counter[0]), .O(n23));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_DFF rand_setpoint_2359__i0 (.Q(rand_setpoint[0]), .C(CLK_c), .D(n165));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 i51_4_lut (.I0(n8_adj_2445), .I1(\data_out[10] [0]), .I2(byte_transmit_counter[1]), 
            .I3(byte_transmit_counter[0]), .O(n32));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i51_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i52_3_lut (.I0(n23), .I1(n6_adj_2446), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n29));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i52_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49_4_lut (.I0(n29), .I1(n32), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n26));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i49_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i50_4_lut (.I0(r_Tx_Data[0]), .I1(n26), .I2(n9257), .I3(byte_transmit_counter[4]), 
            .O(n16924));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i50_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF blink_counter_2360__i0 (.Q(n26_adj_2423), .C(CLK_c), .D(n135_adj_2433));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i24_4_lut_adj_773 (.I0(n18187), .I1(n10_adj_2422), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10_adj_2443));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_4_lut_adj_773.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut_adj_774 (.I0(r_Tx_Data[6]), .I1(n10_adj_2443), .I2(n9257), 
            .I3(byte_transmit_counter[4]), .O(n16914));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i23_4_lut_adj_774.LUT_INIT = 16'h0aca;
    SB_LUT4 i8463_3_lut (.I0(\data_out_frame2[5] [0]), .I1(rand_data[24]), 
            .I2(n10725), .I3(GND_net), .O(n11149));   // coms.v(416[12] 543[6])
    defparam i8463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8464_3_lut (.I0(\data_out_frame2[5] [1]), .I1(rand_data[25]), 
            .I2(n10725), .I3(GND_net), .O(n11150));   // coms.v(416[12] 543[6])
    defparam i8464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8465_3_lut (.I0(\data_out_frame2[5] [2]), .I1(rand_data[26]), 
            .I2(n10725), .I3(GND_net), .O(n11151));   // coms.v(416[12] 543[6])
    defparam i8465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[6]), .I3(r_Bit_Index[1]), .O(n18196));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i8466_3_lut (.I0(\data_out_frame2[5] [3]), .I1(rand_data[27]), 
            .I2(n10725), .I3(GND_net), .O(n11152));   // coms.v(416[12] 543[6])
    defparam i8466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n18196_bdd_4_lut (.I0(n18196), .I1(r_Tx_Data[4]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n18199));
    defparam n18196_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8297_3_lut (.I0(n11018), .I1(r_Bit_Index_adj_2499[0]), .I2(n17361), 
            .I3(GND_net), .O(n10983));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8297_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i8467_3_lut (.I0(\data_out_frame2[5] [4]), .I1(rand_data[28]), 
            .I2(n10725), .I3(GND_net), .O(n11153));   // coms.v(416[12] 543[6])
    defparam i8467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23_4_lut_adj_775 (.I0(byte_transmit_counter[0]), .I1(tx_transmit_N_1947[0]), 
            .I2(n10705), .I3(n10_adj_2444), .O(n16628));   // coms.v(280[12] 370[6])
    defparam i23_4_lut_adj_775.LUT_INIT = 16'hca0a;
    SB_LUT4 i8291_3_lut (.I0(n10976), .I1(r_Bit_Index_adj_2505[0]), .I2(n17412), 
            .I3(GND_net), .O(n10977));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8291_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i8468_3_lut (.I0(\data_out_frame2[5] [5]), .I1(rand_data[29]), 
            .I2(n10725), .I3(GND_net), .O(n11154));   // coms.v(416[12] 543[6])
    defparam i8468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8469_3_lut (.I0(\data_out_frame2[5] [6]), .I1(rand_data[30]), 
            .I2(n10725), .I3(GND_net), .O(n11155));   // coms.v(416[12] 543[6])
    defparam i8469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8288_2_lut (.I0(n5142), .I1(n10972), .I2(GND_net), .I3(GND_net), 
            .O(n10974));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8288_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8470_3_lut (.I0(\data_out_frame2[5] [7]), .I1(rand_data[31]), 
            .I2(n10725), .I3(GND_net), .O(n11156));   // coms.v(416[12] 543[6])
    defparam i8470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8471_3_lut (.I0(\data_out_frame2[6] [0]), .I1(rand_data[16]), 
            .I2(n10725), .I3(GND_net), .O(n11157));   // coms.v(416[12] 543[6])
    defparam i8471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8472_3_lut (.I0(\data_out_frame2[6] [1]), .I1(rand_data[17]), 
            .I2(n10725), .I3(GND_net), .O(n11158));   // coms.v(416[12] 543[6])
    defparam i8472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8285_2_lut (.I0(n5142), .I1(n10969), .I2(GND_net), .I3(GND_net), 
            .O(n10971));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8285_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8473_3_lut (.I0(\data_out_frame2[6] [2]), .I1(rand_data[18]), 
            .I2(n10725), .I3(GND_net), .O(n11159));   // coms.v(416[12] 543[6])
    defparam i8473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8474_3_lut (.I0(\data_out_frame2[6] [3]), .I1(rand_data[19]), 
            .I2(n10725), .I3(GND_net), .O(n11160));   // coms.v(416[12] 543[6])
    defparam i8474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8282_2_lut (.I0(n5142), .I1(n10966), .I2(GND_net), .I3(GND_net), 
            .O(n10968));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8282_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8475_3_lut (.I0(\data_out_frame2[6] [4]), .I1(rand_data[20]), 
            .I2(n10725), .I3(GND_net), .O(n11161));   // coms.v(416[12] 543[6])
    defparam i8475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8279_2_lut (.I0(n5142), .I1(n10963), .I2(GND_net), .I3(GND_net), 
            .O(n10965));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8279_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8476_3_lut (.I0(\data_out_frame2[6] [5]), .I1(rand_data[21]), 
            .I2(n10725), .I3(GND_net), .O(n11162));   // coms.v(416[12] 543[6])
    defparam i8476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8477_3_lut (.I0(\data_out_frame2[6] [6]), .I1(rand_data[22]), 
            .I2(n10725), .I3(GND_net), .O(n11163));   // coms.v(416[12] 543[6])
    defparam i8477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8276_2_lut (.I0(n5142), .I1(n10960), .I2(GND_net), .I3(GND_net), 
            .O(n10962));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8276_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8273_2_lut (.I0(n5142), .I1(n10957), .I2(GND_net), .I3(GND_net), 
            .O(n10959));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8273_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8478_3_lut (.I0(\data_out_frame2[6] [7]), .I1(rand_data[23]), 
            .I2(n10725), .I3(GND_net), .O(n11164));   // coms.v(416[12] 543[6])
    defparam i8478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8270_2_lut (.I0(n5142), .I1(n10954), .I2(GND_net), .I3(GND_net), 
            .O(n10956));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8270_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8479_3_lut (.I0(\data_out_frame2[7] [0]), .I1(rand_data[8]), 
            .I2(n10725), .I3(GND_net), .O(n11165));   // coms.v(416[12] 543[6])
    defparam i8479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8480_3_lut (.I0(\data_out_frame2[7] [1]), .I1(rand_data[9]), 
            .I2(n10725), .I3(GND_net), .O(n11166));   // coms.v(416[12] 543[6])
    defparam i8480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8481_3_lut (.I0(\data_out_frame2[7] [2]), .I1(rand_data[10]), 
            .I2(n10725), .I3(GND_net), .O(n11167));   // coms.v(416[12] 543[6])
    defparam i8481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8482_3_lut (.I0(\data_out_frame2[7] [3]), .I1(rand_data[11]), 
            .I2(n10725), .I3(GND_net), .O(n11168));   // coms.v(416[12] 543[6])
    defparam i8482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8483_3_lut (.I0(\data_out_frame2[7] [4]), .I1(rand_data[12]), 
            .I2(n10725), .I3(GND_net), .O(n11169));   // coms.v(416[12] 543[6])
    defparam i8483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8267_2_lut (.I0(n5142), .I1(n10951), .I2(GND_net), .I3(GND_net), 
            .O(n10953));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8267_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8484_3_lut (.I0(\data_out_frame2[7] [5]), .I1(rand_data[13]), 
            .I2(n10725), .I3(GND_net), .O(n11170));   // coms.v(416[12] 543[6])
    defparam i8484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8485_3_lut (.I0(\data_out_frame2[7] [6]), .I1(rand_data[14]), 
            .I2(n10725), .I3(GND_net), .O(n11171));   // coms.v(416[12] 543[6])
    defparam i8485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8486_3_lut (.I0(\data_out_frame2[7] [7]), .I1(rand_data[15]), 
            .I2(n10725), .I3(GND_net), .O(n11172));   // coms.v(416[12] 543[6])
    defparam i8486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8487_3_lut (.I0(\data_out_frame2[8] [0]), .I1(rand_data[0]), 
            .I2(n10725), .I3(GND_net), .O(n11173));   // coms.v(416[12] 543[6])
    defparam i8487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8488_3_lut (.I0(\data_out_frame2[8] [1]), .I1(rand_data[1]), 
            .I2(n10725), .I3(GND_net), .O(n11174));   // coms.v(416[12] 543[6])
    defparam i8488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8489_3_lut (.I0(\data_out_frame2[8] [2]), .I1(rand_data[2]), 
            .I2(n10725), .I3(GND_net), .O(n11175));   // coms.v(416[12] 543[6])
    defparam i8489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2360_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[25]), .I3(n16065), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2360_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[24]), .I3(n16064), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_26 (.CI(n16064), .I0(GND_net), .I1(blink_counter[24]), 
            .CO(n16065));
    SB_LUT4 rand_setpoint_2359_add_4_32_lut (.I0(GND_net), .I1(rand_data[30]), 
            .I2(rand_setpoint[30]), .I3(n16039), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_5 (.CI(n16012), .I0(rand_data[3]), 
            .I1(rand_setpoint[3]), .CO(n16013));
    SB_CARRY rand_setpoint_2359_add_4_32 (.CI(n16039), .I0(rand_data[30]), 
            .I1(rand_setpoint[30]), .CO(n16040));
    SB_LUT4 blink_counter_2360_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[23]), .I3(n16063), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_31_lut (.I0(GND_net), .I1(rand_data[29]), 
            .I2(rand_setpoint[29]), .I3(n16038), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_4_lut (.I0(GND_net), .I1(rand_data[2]), 
            .I2(rand_setpoint[2]), .I3(n16011), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_25 (.CI(n16063), .I0(GND_net), .I1(blink_counter[23]), 
            .CO(n16064));
    SB_CARRY rand_setpoint_2359_add_4_31 (.CI(n16038), .I0(rand_data[29]), 
            .I1(rand_setpoint[29]), .CO(n16039));
    SB_CARRY rand_setpoint_2359_add_4_4 (.CI(n16011), .I0(rand_data[2]), 
            .I1(rand_setpoint[2]), .CO(n16012));
    SB_LUT4 rand_setpoint_2359_add_4_30_lut (.I0(GND_net), .I1(rand_data[28]), 
            .I2(rand_setpoint[28]), .I3(n16037), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2360_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[22]), .I3(n16062), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_30 (.CI(n16037), .I0(rand_data[28]), 
            .I1(rand_setpoint[28]), .CO(n16038));
    SB_LUT4 rand_setpoint_2359_add_4_3_lut (.I0(GND_net), .I1(rand_data[1]), 
            .I2(rand_setpoint[1]), .I3(n16010), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_24 (.CI(n16062), .I0(GND_net), .I1(blink_counter[22]), 
            .CO(n16063));
    SB_LUT4 rand_setpoint_2359_add_4_29_lut (.I0(GND_net), .I1(rand_data[27]), 
            .I2(rand_setpoint[27]), .I3(n16036), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_3 (.CI(n16010), .I0(rand_data[1]), 
            .I1(rand_setpoint[1]), .CO(n16011));
    SB_CARRY rand_setpoint_2359_add_4_29 (.CI(n16036), .I0(rand_data[27]), 
            .I1(rand_setpoint[27]), .CO(n16037));
    SB_LUT4 blink_counter_2360_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[21]), .I3(n16061), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_28_lut (.I0(GND_net), .I1(rand_data[26]), 
            .I2(rand_setpoint[26]), .I3(n16035), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8490_3_lut (.I0(\data_out_frame2[8] [3]), .I1(rand_data[3]), 
            .I2(n10725), .I3(GND_net), .O(n11176));   // coms.v(416[12] 543[6])
    defparam i8490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2359_add_4_2_lut (.I0(GND_net), .I1(rand_data[0]), 
            .I2(rand_setpoint[0]), .I3(GND_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_23 (.CI(n16061), .I0(GND_net), .I1(blink_counter[21]), 
            .CO(n16062));
    SB_LUT4 i8491_3_lut (.I0(\data_out_frame2[8] [4]), .I1(rand_data[4]), 
            .I2(n10725), .I3(GND_net), .O(n11177));   // coms.v(416[12] 543[6])
    defparam i8491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2360_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_2429), .I3(n16060), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_28 (.CI(n16035), .I0(rand_data[26]), 
            .I1(rand_setpoint[26]), .CO(n16036));
    SB_CARRY rand_setpoint_2359_add_4_2 (.CI(GND_net), .I0(rand_data[0]), 
            .I1(rand_setpoint[0]), .CO(n16010));
    SB_LUT4 rand_setpoint_2359_add_4_27_lut (.I0(GND_net), .I1(rand_data[25]), 
            .I2(rand_setpoint[25]), .I3(n16034), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_22 (.CI(n16060), .I0(GND_net), .I1(n6_adj_2429), 
            .CO(n16061));
    SB_CARRY rand_setpoint_2359_add_4_27 (.CI(n16034), .I0(rand_data[25]), 
            .I1(rand_setpoint[25]), .CO(n16035));
    SB_LUT4 rand_data_2358_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[31]), 
            .I3(n16009), .O(n134_adj_2451)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2360_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7), .I3(n16059), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_26_lut (.I0(GND_net), .I1(rand_data[24]), 
            .I2(rand_setpoint[24]), .I3(n16033), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[30]), 
            .I3(n16008), .O(n135_adj_2452)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[9]), 
            .I3(n15987), .O(n156_adj_2473)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_32 (.CI(n16008), .I0(GND_net), .I1(rand_data[30]), 
            .CO(n16009));
    SB_CARRY blink_counter_2360_add_4_21 (.CI(n16059), .I0(GND_net), .I1(n7), 
            .CO(n16060));
    SB_CARRY rand_setpoint_2359_add_4_26 (.CI(n16033), .I0(rand_data[24]), 
            .I1(rand_setpoint[24]), .CO(n16034));
    SB_LUT4 rand_data_2358_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[29]), 
            .I3(n16007), .O(n136_adj_2453)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_11 (.CI(n15987), .I0(GND_net), .I1(rand_data[9]), 
            .CO(n15988));
    SB_LUT4 blink_counter_2360_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_2412), .I3(n16058), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_25_lut (.I0(GND_net), .I1(rand_data[23]), 
            .I2(rand_setpoint[23]), .I3(n16032), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_31 (.CI(n16007), .I0(GND_net), .I1(rand_data[29]), 
            .CO(n16008));
    SB_LUT4 i53_4_lut_adj_776 (.I0(\data_out[5] [1]), .I1(n5_adj_2448), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n31));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i53_4_lut_adj_776.LUT_INIT = 16'hcac0;
    SB_LUT4 rand_data_2358_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[8]), 
            .I3(n15986), .O(n157_adj_2474)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[28]), 
            .I3(n16006), .O(n137_adj_2454)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut_15385 (.I0(r_Bit_Index[2]), .I1(r_Tx_Data[3]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n18070));
    defparam r_Bit_Index_2__bdd_4_lut_15385.LUT_INIT = 16'he4aa;
    SB_CARRY blink_counter_2360_add_4_20 (.CI(n16058), .I0(GND_net), .I1(n8_adj_2412), 
            .CO(n16059));
    SB_CARRY rand_setpoint_2359_add_4_25 (.CI(n16032), .I0(rand_data[23]), 
            .I1(rand_setpoint[23]), .CO(n16033));
    SB_CARRY rand_data_2358_add_4_30 (.CI(n16006), .I0(GND_net), .I1(rand_data[28]), 
            .CO(n16007));
    SB_CARRY rand_data_2358_add_4_10 (.CI(n15986), .I0(GND_net), .I1(rand_data[8]), 
            .CO(n15987));
    SB_LUT4 blink_counter_2360_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_2421), .I3(n16057), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_24_lut (.I0(GND_net), .I1(rand_data[22]), 
            .I2(rand_setpoint[22]), .I3(n16031), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_24 (.CI(n16031), .I0(rand_data[22]), 
            .I1(rand_setpoint[22]), .CO(n16032));
    SB_LUT4 rand_data_2358_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[27]), 
            .I3(n16005), .O(n138_adj_2455)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[7]), 
            .I3(n15985), .O(n158_adj_2475)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52_4_lut (.I0(n8_adj_2447), .I1(\data_out[10] [1]), .I2(byte_transmit_counter[1]), 
            .I3(byte_transmit_counter[0]), .O(n25));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i52_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY rand_data_2358_add_4_9 (.CI(n15985), .I0(GND_net), .I1(rand_data[7]), 
            .CO(n15986));
    SB_LUT4 i49_4_lut_adj_777 (.I0(n1_adj_2449), .I1(n31), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n22));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i49_4_lut_adj_777.LUT_INIT = 16'hc0ca;
    SB_LUT4 i51_4_lut_adj_778 (.I0(n22), .I1(n25), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n28));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i51_4_lut_adj_778.LUT_INIT = 16'h0aca;
    SB_CARRY blink_counter_2360_add_4_19 (.CI(n16057), .I0(GND_net), .I1(n9_adj_2421), 
            .CO(n16058));
    SB_LUT4 rand_setpoint_2359_add_4_23_lut (.I0(GND_net), .I1(rand_data[21]), 
            .I2(rand_setpoint[21]), .I3(n16030), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50_4_lut_adj_779 (.I0(r_Tx_Data[1]), .I1(n28), .I2(n9257), 
            .I3(byte_transmit_counter[4]), .O(n16926));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i50_4_lut_adj_779.LUT_INIT = 16'h0aca;
    SB_LUT4 blink_counter_2360_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_2420), .I3(n16056), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_18 (.CI(n16056), .I0(GND_net), .I1(n10_adj_2420), 
            .CO(n16057));
    SB_CARRY rand_setpoint_2359_add_4_23 (.CI(n16030), .I0(rand_data[21]), 
            .I1(rand_setpoint[21]), .CO(n16031));
    SB_CARRY rand_data_2358_add_4_29 (.CI(n16005), .I0(GND_net), .I1(rand_data[27]), 
            .CO(n16006));
    SB_LUT4 rand_data_2358_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[6]), 
            .I3(n15984), .O(n159_adj_2476)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[26]), 
            .I3(n16004), .O(n139_adj_2456)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2360_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11), .I3(n16055), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24_4_lut_adj_780 (.I0(n18169), .I1(n10_adj_2450), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10_adj_2411));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_4_lut_adj_780.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut_adj_781 (.I0(r_Tx_Data[2]), .I1(n10_adj_2411), .I2(n9257), 
            .I3(byte_transmit_counter[4]), .O(n16928));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i23_4_lut_adj_781.LUT_INIT = 16'h0aca;
    SB_LUT4 rand_setpoint_2359_add_4_22_lut (.I0(GND_net), .I1(rand_data[20]), 
            .I2(rand_setpoint[20]), .I3(n16029), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_28 (.CI(n16004), .I0(GND_net), .I1(rand_data[26]), 
            .CO(n16005));
    SB_CARRY rand_data_2358_add_4_8 (.CI(n15984), .I0(GND_net), .I1(rand_data[6]), 
            .CO(n15985));
    SB_CARRY blink_counter_2360_add_4_17 (.CI(n16055), .I0(GND_net), .I1(n11), 
            .CO(n16056));
    SB_CARRY rand_setpoint_2359_add_4_22 (.CI(n16029), .I0(rand_data[20]), 
            .I1(rand_setpoint[20]), .CO(n16030));
    SB_LUT4 i24_4_lut_adj_782 (.I0(n18175), .I1(n10_adj_2431), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10_adj_2409));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_4_lut_adj_782.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut_adj_783 (.I0(r_Tx_Data[3]), .I1(n10_adj_2409), .I2(n9257), 
            .I3(byte_transmit_counter[4]), .O(n16930));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i23_4_lut_adj_783.LUT_INIT = 16'h0aca;
    SB_LUT4 rand_data_2358_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[25]), 
            .I3(n16003), .O(n140_adj_2457)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2360_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12), .I3(n16054), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_21_lut (.I0(GND_net), .I1(rand_data[19]), 
            .I2(rand_setpoint[19]), .I3(n16028), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[5]), 
            .I3(n15983), .O(n160_adj_2477)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[3]), 
            .I3(n15981), .O(n162_adj_2479)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_27 (.CI(n16003), .I0(GND_net), .I1(rand_data[25]), 
            .CO(n16004));
    SB_CARRY blink_counter_2360_add_4_16 (.CI(n16054), .I0(GND_net), .I1(n12), 
            .CO(n16055));
    SB_CARRY rand_setpoint_2359_add_4_21 (.CI(n16028), .I0(rand_data[19]), 
            .I1(rand_setpoint[19]), .CO(n16029));
    SB_LUT4 rand_data_2358_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[24]), 
            .I3(n16002), .O(n141_adj_2458)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_7 (.CI(n15983), .I0(GND_net), .I1(rand_data[5]), 
            .CO(n15984));
    SB_LUT4 blink_counter_2360_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n16053), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_20_lut (.I0(GND_net), .I1(rand_data[18]), 
            .I2(rand_setpoint[18]), .I3(n16027), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24_4_lut_adj_784 (.I0(n18271), .I1(n10_adj_2430), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10_adj_2408));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_4_lut_adj_784.LUT_INIT = 16'h0aca;
    SB_CARRY rand_data_2358_add_4_26 (.CI(n16002), .I0(GND_net), .I1(rand_data[24]), 
            .CO(n16003));
    SB_LUT4 i23_4_lut_adj_785 (.I0(r_Tx_Data[4]), .I1(n10_adj_2408), .I2(n9257), 
            .I3(byte_transmit_counter[4]), .O(n16932));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i23_4_lut_adj_785.LUT_INIT = 16'h0aca;
    SB_LUT4 rand_data_2358_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[23]), 
            .I3(n16001), .O(n142_adj_2459)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_20 (.CI(n16027), .I0(rand_data[18]), 
            .I1(rand_setpoint[18]), .CO(n16028));
    SB_LUT4 rand_data_2358_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[4]), 
            .I3(n15982), .O(n161_adj_2478)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_15 (.CI(n16053), .I0(GND_net), .I1(n13), 
            .CO(n16054));
    SB_LUT4 rand_setpoint_2359_add_4_19_lut (.I0(GND_net), .I1(rand_data[17]), 
            .I2(rand_setpoint[17]), .I3(n16026), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2360_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n16052), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_19 (.CI(n16026), .I0(rand_data[17]), 
            .I1(rand_setpoint[17]), .CO(n16027));
    SB_CARRY rand_data_2358_add_4_25 (.CI(n16001), .I0(GND_net), .I1(rand_data[23]), 
            .CO(n16002));
    SB_LUT4 rand_setpoint_2359_add_4_18_lut (.I0(GND_net), .I1(rand_data[16]), 
            .I2(rand_setpoint[16]), .I3(n16025), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23_4_lut_adj_786 (.I0(byte_transmit_counter[5]), .I1(tx_transmit_N_1947[5]), 
            .I2(n10705), .I3(n10_adj_2444), .O(n16630));   // coms.v(280[12] 370[6])
    defparam i23_4_lut_adj_786.LUT_INIT = 16'hca0a;
    SB_CARRY blink_counter_2360_add_4_14 (.CI(n16052), .I0(GND_net), .I1(n14), 
            .CO(n16053));
    SB_CARRY rand_setpoint_2359_add_4_18 (.CI(n16025), .I0(rand_data[16]), 
            .I1(rand_setpoint[16]), .CO(n16026));
    SB_LUT4 rand_data_2358_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[22]), 
            .I3(n16000), .O(n143_adj_2460)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_DFF blink_counter_2360__i25 (.Q(blink_counter[25]), .C(CLK_c), .D(n110));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i24 (.Q(blink_counter[24]), .C(CLK_c), .D(n111));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i23 (.Q(blink_counter[23]), .C(CLK_c), .D(n112));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i22 (.Q(blink_counter[22]), .C(CLK_c), .D(n113));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i21 (.Q(blink_counter[21]), .C(CLK_c), .D(n114));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 blink_counter_2360_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15), .I3(n16051), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rand_setpoint_2359_add_4_17_lut (.I0(GND_net), .I1(rand_data[15]), 
            .I2(rand_setpoint[15]), .I3(n16024), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF blink_counter_2360__i20 (.Q(n6_adj_2429), .C(CLK_c), .D(n115));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i23_4_lut_adj_787 (.I0(byte_transmit_counter[6]), .I1(tx_transmit_N_1947[6]), 
            .I2(n10705), .I3(n10_adj_2444), .O(n16632));   // coms.v(280[12] 370[6])
    defparam i23_4_lut_adj_787.LUT_INIT = 16'hca0a;
    SB_DFF blink_counter_2360__i19 (.Q(n7), .C(CLK_c), .D(n116));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i18 (.Q(n8_adj_2412), .C(CLK_c), .D(n117));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_CARRY rand_data_2358_add_4_24 (.CI(n16000), .I0(GND_net), .I1(rand_data[22]), 
            .CO(n16001));
    SB_CARRY rand_setpoint_2359_add_4_17 (.CI(n16024), .I0(rand_data[15]), 
            .I1(rand_setpoint[15]), .CO(n16025));
    SB_LUT4 i2_2_lut (.I0(\UART_TRANSMITTER.state [1]), .I1(n4_adj_2419), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_2407));   // coms.v(280[12] 370[6])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_DFF blink_counter_2360__i17 (.Q(n9_adj_2421), .C(CLK_c), .D(n118));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i16 (.Q(n10_adj_2420), .C(CLK_c), .D(n119));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i15 (.Q(n11), .C(CLK_c), .D(n120));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i14 (.Q(n12), .C(CLK_c), .D(n121));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_CARRY blink_counter_2360_add_4_13 (.CI(n16051), .I0(GND_net), .I1(n15), 
            .CO(n16052));
    SB_LUT4 rand_setpoint_2359_add_4_16_lut (.I0(GND_net), .I1(rand_data[14]), 
            .I2(rand_setpoint[14]), .I3(n16023), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n18070_bdd_4_lut (.I0(n18070), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[1]), 
            .I3(r_Bit_Index[1]), .O(n18073));
    defparam n18070_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rand_data_2358_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[21]), 
            .I3(n15999), .O(n144_adj_2461)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF blink_counter_2360__i13 (.Q(n13), .C(CLK_c), .D(n122));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i12 (.Q(n14), .C(CLK_c), .D(n123));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i11 (.Q(n15), .C(CLK_c), .D(n124));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i10 (.Q(n16), .C(CLK_c), .D(n125));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i9 (.Q(n17), .C(CLK_c), .D(n126));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i8 (.Q(n18), .C(CLK_c), .D(n127));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i7 (.Q(n19), .C(CLK_c), .D(n128));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i6 (.Q(n20), .C(CLK_c), .D(n129));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i5 (.Q(n21), .C(CLK_c), .D(n130));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i4 (.Q(n22_adj_2426), .C(CLK_c), .D(n131));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i3 (.Q(n23_adj_2425), .C(CLK_c), .D(n132));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2360__i2 (.Q(n24), .C(CLK_c), .D(n133));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i15020_4_lut (.I0(n9524), .I1(n444), .I2(n17327), .I3(tx_transmit_N_1947[3]), 
            .O(n17664));   // coms.v(280[12] 370[6])
    defparam i15020_4_lut.LUT_INIT = 16'hcddd;
    SB_LUT4 blink_counter_2360_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n16050), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF blink_counter_2360__i1 (.Q(n25_adj_2424), .C(CLK_c), .D(n134_adj_2434));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i24_4_lut_adj_788 (.I0(n5_adj_2407), .I1(n17664), .I2(\UART_TRANSMITTER.state [2]), 
            .I3(\UART_TRANSMITTER.state [0]), .O(n10_adj_2444));   // coms.v(280[12] 370[6])
    defparam i24_4_lut_adj_788.LUT_INIT = 16'h0aca;
    SB_CARRY rand_setpoint_2359_add_4_16 (.CI(n16023), .I0(rand_data[14]), 
            .I1(rand_setpoint[14]), .CO(n16024));
    SB_CARRY rand_data_2358_add_4_23 (.CI(n15999), .I0(GND_net), .I1(rand_data[21]), 
            .CO(n16000));
    SB_LUT4 rand_setpoint_2359_add_4_15_lut (.I0(GND_net), .I1(rand_data[13]), 
            .I2(rand_setpoint[13]), .I3(n16022), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_12 (.CI(n16050), .I0(GND_net), .I1(n16), 
            .CO(n16051));
    SB_CARRY rand_setpoint_2359_add_4_15 (.CI(n16022), .I0(rand_data[13]), 
            .I1(rand_setpoint[13]), .CO(n16023));
    SB_LUT4 i23_4_lut_adj_789 (.I0(byte_transmit_counter[7]), .I1(tx_transmit_N_1947[7]), 
            .I2(n10705), .I3(n10_adj_2444), .O(n16634));   // coms.v(280[12] 370[6])
    defparam i23_4_lut_adj_789.LUT_INIT = 16'hca0a;
    SB_LUT4 i8237_4_lut (.I0(n10976), .I1(r_Bit_Index_adj_2505[1]), .I2(r_Bit_Index_adj_2505[0]), 
            .I3(n17412), .O(n10923));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8237_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 rand_data_2358_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[20]), 
            .I3(n15998), .O(n145_adj_2462)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_22 (.CI(n15998), .I0(GND_net), .I1(rand_data[20]), 
            .CO(n15999));
    SB_LUT4 blink_counter_2360_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17), .I3(n16049), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_14_lut (.I0(GND_net), .I1(rand_data[12]), 
            .I2(rand_setpoint[12]), .I3(n16021), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[19]), 
            .I3(n15997), .O(n146_adj_2463)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_14 (.CI(n16021), .I0(rand_data[12]), 
            .I1(rand_setpoint[12]), .CO(n16022));
    SB_CARRY blink_counter_2360_add_4_11 (.CI(n16049), .I0(GND_net), .I1(n17), 
            .CO(n16050));
    SB_LUT4 rand_setpoint_2359_add_4_13_lut (.I0(GND_net), .I1(rand_data[11]), 
            .I2(rand_setpoint[11]), .I3(n16020), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_21 (.CI(n15997), .I0(GND_net), .I1(rand_data[19]), 
            .CO(n15998));
    SB_LUT4 rand_data_2358_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[18]), 
            .I3(n15996), .O(n147_adj_2464)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8492_3_lut (.I0(\data_out_frame2[8] [5]), .I1(rand_data[5]), 
            .I2(n10725), .I3(GND_net), .O(n11178));   // coms.v(416[12] 543[6])
    defparam i8492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2360_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18), .I3(n16048), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_13 (.CI(n16020), .I0(rand_data[11]), 
            .I1(rand_setpoint[11]), .CO(n16021));
    SB_CARRY rand_data_2358_add_4_20 (.CI(n15996), .I0(GND_net), .I1(rand_data[18]), 
            .CO(n15997));
    SB_LUT4 i8493_3_lut (.I0(\data_out_frame2[8] [6]), .I1(rand_data[6]), 
            .I2(n10725), .I3(GND_net), .O(n11179));   // coms.v(416[12] 543[6])
    defparam i8493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2358_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[17]), 
            .I3(n15995), .O(n148_adj_2465)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_10 (.CI(n16048), .I0(GND_net), .I1(n18), 
            .CO(n16049));
    SB_LUT4 rand_setpoint_2359_add_4_12_lut (.I0(GND_net), .I1(rand_data[10]), 
            .I2(rand_setpoint[10]), .I3(n16019), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_19 (.CI(n15995), .I0(GND_net), .I1(rand_data[17]), 
            .CO(n15996));
    SB_LUT4 blink_counter_2360_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19), .I3(n16047), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_12 (.CI(n16019), .I0(rand_data[10]), 
            .I1(rand_setpoint[10]), .CO(n16020));
    SB_LUT4 rand_data_2358_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[16]), 
            .I3(n15994), .O(n149_adj_2466)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_5 (.CI(n15981), .I0(GND_net), .I1(rand_data[3]), 
            .CO(n15982));
    SB_CARRY rand_data_2358_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(rand_data[0]), 
            .CO(n15979));
    SB_CARRY rand_data_2358_add_4_18 (.CI(n15994), .I0(GND_net), .I1(rand_data[16]), 
            .CO(n15995));
    SB_CARRY blink_counter_2360_add_4_9 (.CI(n16047), .I0(GND_net), .I1(n19), 
            .CO(n16048));
    SB_LUT4 rand_setpoint_2359_add_4_11_lut (.I0(GND_net), .I1(rand_data[9]), 
            .I2(rand_setpoint[9]), .I3(n16018), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[15]), 
            .I3(n15993), .O(n150_adj_2467)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[2]), 
            .I3(n15980), .O(n163_adj_2480)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2360_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20), .I3(n16046), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2359_add_4_11 (.CI(n16018), .I0(rand_data[9]), 
            .I1(rand_setpoint[9]), .CO(n16019));
    SB_CARRY rand_data_2358_add_4_17 (.CI(n15993), .I0(GND_net), .I1(rand_data[15]), 
            .CO(n15994));
    SB_CARRY rand_data_2358_add_4_4 (.CI(n15980), .I0(GND_net), .I1(rand_data[2]), 
            .CO(n15981));
    SB_CARRY blink_counter_2360_add_4_8 (.CI(n16046), .I0(GND_net), .I1(n20), 
            .CO(n16047));
    SB_LUT4 rand_data_2358_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[14]), 
            .I3(n15992), .O(n151_adj_2468)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_setpoint_2359__i31 (.Q(rand_setpoint[31]), .C(CLK_c), .D(n134));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 blink_counter_2360_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21), .I3(n16045), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8494_3_lut (.I0(\data_out_frame2[8] [7]), .I1(rand_data[7]), 
            .I2(n10725), .I3(GND_net), .O(n11180));   // coms.v(416[12] 543[6])
    defparam i8494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2359_add_4_10_lut (.I0(GND_net), .I1(rand_data[8]), 
            .I2(rand_setpoint[8]), .I3(n16017), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_16 (.CI(n15992), .I0(GND_net), .I1(rand_data[14]), 
            .CO(n15993));
    SB_LUT4 rand_data_2358_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[13]), 
            .I3(n15991), .O(n152_adj_2469)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_7 (.CI(n16045), .I0(GND_net), .I1(n21), 
            .CO(n16046));
    SB_CARRY rand_setpoint_2359_add_4_10 (.CI(n16017), .I0(rand_data[8]), 
            .I1(rand_setpoint[8]), .CO(n16018));
    SB_LUT4 i8495_3_lut (.I0(\data_out_frame2[9] [0]), .I1(rand_data[24]), 
            .I2(n10725), .I3(GND_net), .O(n11181));   // coms.v(416[12] 543[6])
    defparam i8495_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2358_add_4_15 (.CI(n15991), .I0(GND_net), .I1(rand_data[13]), 
            .CO(n15992));
    SB_LUT4 i8496_3_lut (.I0(\data_out_frame2[9] [1]), .I1(rand_data[25]), 
            .I2(n10725), .I3(GND_net), .O(n11182));   // coms.v(416[12] 543[6])
    defparam i8496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2360_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_2426), .I3(n16044), .O(n131)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2359_add_4_9_lut (.I0(GND_net), .I1(rand_data[7]), 
            .I2(rand_setpoint[7]), .I3(n16016), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[12]), 
            .I3(n15990), .O(n153_adj_2470)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2358_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[1]), 
            .I3(n15979), .O(n164_adj_2481)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_14 (.CI(n15990), .I0(GND_net), .I1(rand_data[12]), 
            .CO(n15991));
    SB_CARRY blink_counter_2360_add_4_6 (.CI(n16044), .I0(GND_net), .I1(n22_adj_2426), 
            .CO(n16045));
    SB_CARRY rand_setpoint_2359_add_4_9 (.CI(n16016), .I0(rand_data[7]), 
            .I1(rand_setpoint[7]), .CO(n16017));
    SB_LUT4 rand_data_2358_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[11]), 
            .I3(n15989), .O(n154_adj_2471)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2358_add_4_3 (.CI(n15979), .I0(GND_net), .I1(rand_data[1]), 
            .CO(n15980));
    SB_LUT4 rand_data_2358_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[0]), 
            .I3(VCC_net), .O(n165_adj_2482)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8234_4_lut (.I0(n10976), .I1(r_Bit_Index_adj_2505[2]), .I2(n5266), 
            .I3(n17412), .O(n10920));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8234_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 i8497_3_lut (.I0(\data_out_frame2[9] [2]), .I1(rand_data[26]), 
            .I2(n10725), .I3(GND_net), .O(n11183));   // coms.v(416[12] 543[6])
    defparam i8497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8498_3_lut (.I0(\data_out_frame2[9] [3]), .I1(rand_data[27]), 
            .I2(n10725), .I3(GND_net), .O(n11184));   // coms.v(416[12] 543[6])
    defparam i8498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8499_3_lut (.I0(\data_out_frame2[9] [4]), .I1(rand_data[28]), 
            .I2(n10725), .I3(GND_net), .O(n11185));   // coms.v(416[12] 543[6])
    defparam i8499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2360_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_2425), .I3(n16043), .O(n132)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_5 (.CI(n16043), .I0(GND_net), .I1(n23_adj_2425), 
            .CO(n16044));
    SB_LUT4 i8500_3_lut (.I0(\data_out_frame2[9] [5]), .I1(rand_data[29]), 
            .I2(n10725), .I3(GND_net), .O(n11186));   // coms.v(416[12] 543[6])
    defparam i8500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2360_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24), .I3(n16042), .O(n133)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8501_3_lut (.I0(\data_out_frame2[9] [6]), .I1(rand_data[30]), 
            .I2(n10725), .I3(GND_net), .O(n11187));   // coms.v(416[12] 543[6])
    defparam i8501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8502_3_lut (.I0(\data_out_frame2[9] [7]), .I1(rand_data[31]), 
            .I2(n10725), .I3(GND_net), .O(n11188));   // coms.v(416[12] 543[6])
    defparam i8502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8503_3_lut (.I0(\data_out_frame2[10] [0]), .I1(rand_data[16]), 
            .I2(n10725), .I3(GND_net), .O(n11189));   // coms.v(416[12] 543[6])
    defparam i8503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8504_3_lut (.I0(\data_out_frame2[10] [1]), .I1(rand_data[17]), 
            .I2(n10725), .I3(GND_net), .O(n11190));   // coms.v(416[12] 543[6])
    defparam i8504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8505_3_lut (.I0(\data_out_frame2[10] [2]), .I1(rand_data[18]), 
            .I2(n10725), .I3(GND_net), .O(n11191));   // coms.v(416[12] 543[6])
    defparam i8505_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2360_add_4_4 (.CI(n16042), .I0(GND_net), .I1(n24), 
            .CO(n16043));
    SB_LUT4 rand_setpoint_2359_add_4_8_lut (.I0(GND_net), .I1(rand_data[6]), 
            .I2(rand_setpoint[6]), .I3(n16015), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8506_3_lut (.I0(\data_out_frame2[10] [3]), .I1(rand_data[19]), 
            .I2(n10725), .I3(GND_net), .O(n11192));   // coms.v(416[12] 543[6])
    defparam i8506_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2359_add_4_8 (.CI(n16015), .I0(rand_data[6]), 
            .I1(rand_setpoint[6]), .CO(n16016));
    SB_CARRY rand_data_2358_add_4_13 (.CI(n15989), .I0(GND_net), .I1(rand_data[11]), 
            .CO(n15990));
    SB_LUT4 i8507_3_lut (.I0(\data_out_frame2[10] [4]), .I1(rand_data[20]), 
            .I2(n10725), .I3(GND_net), .O(n11193));   // coms.v(416[12] 543[6])
    defparam i8507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8508_3_lut (.I0(\data_out_frame2[10] [5]), .I1(rand_data[21]), 
            .I2(n10725), .I3(GND_net), .O(n11194));   // coms.v(416[12] 543[6])
    defparam i8508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2359_add_4_7_lut (.I0(GND_net), .I1(rand_data[5]), 
            .I2(rand_setpoint[5]), .I3(n16014), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_setpoint_2359__i30 (.Q(rand_setpoint[30]), .C(CLK_c), .D(n135));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i29 (.Q(rand_setpoint[29]), .C(CLK_c), .D(n136));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i28 (.Q(rand_setpoint[28]), .C(CLK_c), .D(n137));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i27 (.Q(rand_setpoint[27]), .C(CLK_c), .D(n138));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i26 (.Q(rand_setpoint[26]), .C(CLK_c), .D(n139));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i25 (.Q(rand_setpoint[25]), .C(CLK_c), .D(n140));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i24 (.Q(rand_setpoint[24]), .C(CLK_c), .D(n141));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i23 (.Q(rand_setpoint[23]), .C(CLK_c), .D(n142));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i22 (.Q(rand_setpoint[22]), .C(CLK_c), .D(n143));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i21 (.Q(rand_setpoint[21]), .C(CLK_c), .D(n144));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i20 (.Q(rand_setpoint[20]), .C(CLK_c), .D(n145));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i19 (.Q(rand_setpoint[19]), .C(CLK_c), .D(n146));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i18 (.Q(rand_setpoint[18]), .C(CLK_c), .D(n147));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i17 (.Q(rand_setpoint[17]), .C(CLK_c), .D(n148));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i16 (.Q(rand_setpoint[16]), .C(CLK_c), .D(n149));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i15 (.Q(rand_setpoint[15]), .C(CLK_c), .D(n150));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i14 (.Q(rand_setpoint[14]), .C(CLK_c), .D(n151));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i13 (.Q(rand_setpoint[13]), .C(CLK_c), .D(n152));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i12 (.Q(rand_setpoint[12]), .C(CLK_c), .D(n153));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i11 (.Q(rand_setpoint[11]), .C(CLK_c), .D(n154));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i10 (.Q(rand_setpoint[10]), .C(CLK_c), .D(n155));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i9 (.Q(rand_setpoint[9]), .C(CLK_c), .D(n156));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i8 (.Q(rand_setpoint[8]), .C(CLK_c), .D(n157));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i7 (.Q(rand_setpoint[7]), .C(CLK_c), .D(n158));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i6 (.Q(rand_setpoint[6]), .C(CLK_c), .D(n159));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i5 (.Q(rand_setpoint[5]), .C(CLK_c), .D(n160));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i4 (.Q(rand_setpoint[4]), .C(CLK_c), .D(n161));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2359__i3 (.Q(rand_setpoint[3]), .C(CLK_c), .D(n162));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 i8509_3_lut (.I0(\data_out_frame2[10] [6]), .I1(rand_data[22]), 
            .I2(n10725), .I3(GND_net), .O(n11195));   // coms.v(416[12] 543[6])
    defparam i8509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8510_3_lut (.I0(\data_out_frame2[10] [7]), .I1(rand_data[23]), 
            .I2(n10725), .I3(GND_net), .O(n11196));   // coms.v(416[12] 543[6])
    defparam i8510_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_setpoint_2359__i2 (.Q(rand_setpoint[2]), .C(CLK_c), .D(n163));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 rand_data_2358_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[10]), 
            .I3(n15988), .O(n155_adj_2472)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2358_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_setpoint_2359__i1 (.Q(rand_setpoint[1]), .C(CLK_c), .D(n164));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 blink_counter_2360_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_2424), .I3(n16041), .O(n134_adj_2434)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_data_2358__i31 (.Q(rand_data[31]), .C(CLK_c), .D(n134_adj_2451));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i30 (.Q(rand_data[30]), .C(CLK_c), .D(n135_adj_2452));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_CARRY rand_data_2358_add_4_12 (.CI(n15988), .I0(GND_net), .I1(rand_data[10]), 
            .CO(n15989));
    SB_LUT4 i8511_3_lut (.I0(\data_out_frame2[11] [0]), .I1(rand_data[8]), 
            .I2(n10725), .I3(GND_net), .O(n11197));   // coms.v(416[12] 543[6])
    defparam i8511_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_data_2358__i29 (.Q(rand_data[29]), .C(CLK_c), .D(n136_adj_2453));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i28 (.Q(rand_data[28]), .C(CLK_c), .D(n137_adj_2454));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_CARRY blink_counter_2360_add_4_3 (.CI(n16041), .I0(GND_net), .I1(n25_adj_2424), 
            .CO(n16042));
    SB_LUT4 i8512_3_lut (.I0(\data_out_frame2[11] [1]), .I1(rand_data[9]), 
            .I2(n10725), .I3(GND_net), .O(n11198));   // coms.v(416[12] 543[6])
    defparam i8512_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_data_2358__i27 (.Q(rand_data[27]), .C(CLK_c), .D(n138_adj_2455));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i26 (.Q(rand_data[26]), .C(CLK_c), .D(n139_adj_2456));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i25 (.Q(rand_data[25]), .C(CLK_c), .D(n140_adj_2457));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i24 (.Q(rand_data[24]), .C(CLK_c), .D(n141_adj_2458));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i8513_3_lut (.I0(\data_out_frame2[11] [2]), .I1(rand_data[10]), 
            .I2(n10725), .I3(GND_net), .O(n11199));   // coms.v(416[12] 543[6])
    defparam i8513_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_data_2358__i23 (.Q(rand_data[23]), .C(CLK_c), .D(n142_adj_2459));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i22 (.Q(rand_data[22]), .C(CLK_c), .D(n143_adj_2460));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i21 (.Q(rand_data[21]), .C(CLK_c), .D(n144_adj_2461));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i20 (.Q(rand_data[20]), .C(CLK_c), .D(n145_adj_2462));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_CARRY rand_setpoint_2359_add_4_7 (.CI(n16014), .I0(rand_data[5]), 
            .I1(rand_setpoint[5]), .CO(n16015));
    SB_DFF rand_data_2358__i19 (.Q(rand_data[19]), .C(CLK_c), .D(n146_adj_2463));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i18 (.Q(rand_data[18]), .C(CLK_c), .D(n147_adj_2464));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i17 (.Q(rand_data[17]), .C(CLK_c), .D(n148_adj_2465));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i16 (.Q(rand_data[16]), .C(CLK_c), .D(n149_adj_2466));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 rand_setpoint_2359_add_4_6_lut (.I0(GND_net), .I1(rand_data[4]), 
            .I2(rand_setpoint[4]), .I3(n16013), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_data_2358__i15 (.Q(rand_data[15]), .C(CLK_c), .D(n150_adj_2467));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i14 (.Q(rand_data[14]), .C(CLK_c), .D(n151_adj_2468));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i13 (.Q(rand_data[13]), .C(CLK_c), .D(n152_adj_2469));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i12 (.Q(rand_data[12]), .C(CLK_c), .D(n153_adj_2470));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i8514_3_lut (.I0(\data_out_frame2[11] [3]), .I1(rand_data[11]), 
            .I2(n10725), .I3(GND_net), .O(n11200));   // coms.v(416[12] 543[6])
    defparam i8514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8515_3_lut (.I0(\data_out_frame2[11] [4]), .I1(rand_data[12]), 
            .I2(n10725), .I3(GND_net), .O(n11201));   // coms.v(416[12] 543[6])
    defparam i8515_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2359_add_4_6 (.CI(n16013), .I0(rand_data[4]), 
            .I1(rand_setpoint[4]), .CO(n16014));
    SB_LUT4 i8516_3_lut (.I0(\data_out_frame2[11] [5]), .I1(rand_data[13]), 
            .I2(n10725), .I3(GND_net), .O(n11202));   // coms.v(416[12] 543[6])
    defparam i8516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8517_3_lut (.I0(\data_out_frame2[11] [6]), .I1(rand_data[14]), 
            .I2(n10725), .I3(GND_net), .O(n11203));   // coms.v(416[12] 543[6])
    defparam i8517_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2358_add_4_6 (.CI(n15982), .I0(GND_net), .I1(rand_data[4]), 
            .CO(n15983));
    SB_LUT4 i8518_3_lut (.I0(\data_out_frame2[11] [7]), .I1(rand_data[15]), 
            .I2(n10725), .I3(GND_net), .O(n11204));   // coms.v(416[12] 543[6])
    defparam i8518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8519_3_lut (.I0(\data_out_frame2[12] [0]), .I1(rand_data[0]), 
            .I2(n10725), .I3(GND_net), .O(n11205));   // coms.v(416[12] 543[6])
    defparam i8519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8225_3_lut (.I0(\data_out[0] [5]), .I1(n2699), .I2(n10596), 
            .I3(GND_net), .O(n10911));   // coms.v(280[12] 370[6])
    defparam i8225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8520_3_lut (.I0(\data_out_frame2[12] [1]), .I1(rand_data[1]), 
            .I2(n10725), .I3(GND_net), .O(n11206));   // coms.v(416[12] 543[6])
    defparam i8520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8521_3_lut (.I0(\data_out_frame2[12] [2]), .I1(rand_data[2]), 
            .I2(n10725), .I3(GND_net), .O(n11207));   // coms.v(416[12] 543[6])
    defparam i8521_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_data_2358__i11 (.Q(rand_data[11]), .C(CLK_c), .D(n154_adj_2471));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i10 (.Q(rand_data[10]), .C(CLK_c), .D(n155_adj_2472));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i9 (.Q(rand_data[9]), .C(CLK_c), .D(n156_adj_2473));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i8 (.Q(rand_data[8]), .C(CLK_c), .D(n157_adj_2474));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i7 (.Q(rand_data[7]), .C(CLK_c), .D(n158_adj_2475));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i6 (.Q(rand_data[6]), .C(CLK_c), .D(n159_adj_2476));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i5 (.Q(rand_data[5]), .C(CLK_c), .D(n160_adj_2477));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i4 (.Q(rand_data[4]), .C(CLK_c), .D(n161_adj_2478));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i3 (.Q(rand_data[3]), .C(CLK_c), .D(n162_adj_2479));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i2 (.Q(rand_data[2]), .C(CLK_c), .D(n163_adj_2480));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2358__i1 (.Q(rand_data[1]), .C(CLK_c), .D(n164_adj_2481));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i8522_3_lut (.I0(\data_out_frame2[12] [3]), .I1(rand_data[3]), 
            .I2(n10725), .I3(GND_net), .O(n11208));   // coms.v(416[12] 543[6])
    defparam i8522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8301_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n9999), 
            .I3(n4_adj_2416), .O(n10987));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8301_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8330_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n17075), 
            .I3(GND_net), .O(n11016));   // coms.v(416[12] 543[6])
    defparam i8330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 blink_counter_2360_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26_adj_2423), .I3(VCC_net), .O(n135_adj_2433)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2360_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8337_3_lut (.I0(\data_in_frame[6] [6]), .I1(rx_data[6]), .I2(n17075), 
            .I3(GND_net), .O(n11023));   // coms.v(416[12] 543[6])
    defparam i8337_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8338_3_lut (.I0(\data_in_frame[6] [5]), .I1(rx_data[5]), .I2(n17075), 
            .I3(GND_net), .O(n11024));   // coms.v(416[12] 543[6])
    defparam i8338_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8339_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n17075), 
            .I3(GND_net), .O(n11025));   // coms.v(416[12] 543[6])
    defparam i8339_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8340_4_lut (.I0(r_SM_Main_adj_2500[2]), .I1(n1), .I2(n13692), 
            .I3(r_SM_Main_adj_2500[1]), .O(n11026));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8340_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i8341_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n17075), 
            .I3(GND_net), .O(n11027));   // coms.v(416[12] 543[6])
    defparam i8341_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8342_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n17075), 
            .I3(GND_net), .O(n11028));   // coms.v(416[12] 543[6])
    defparam i8342_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8346_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n17075), 
            .I3(GND_net), .O(n11032));   // coms.v(416[12] 543[6])
    defparam i8346_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8347_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n17075), 
            .I3(GND_net), .O(n11033));   // coms.v(416[12] 543[6])
    defparam i8347_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8348_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n10010), 
            .I3(n13116), .O(n11034));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8348_4_lut.LUT_INIT = 16'hcacc;
    SB_LUT4 i8351_3_lut (.I0(tx2_o), .I1(n3), .I2(n10674), .I3(GND_net), 
            .O(n11037));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8221_3_lut_4_lut (.I0(\data_out[1] [6]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n10596), .O(n10907));   // coms.v(280[12] 370[6])
    defparam i8221_3_lut_4_lut.LUT_INIT = 16'hc0aa;
    SB_LUT4 i8226_3_lut (.I0(\data_out[0] [3]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n10596), .I3(GND_net), .O(n10912));   // coms.v(280[12] 370[6])
    defparam i8226_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i15178_4_lut (.I0(n450), .I1(\UART_TRANSMITTER.state [0]), .I2(\UART_TRANSMITTER.state [1]), 
            .I3(n4_adj_2414), .O(n17759));   // coms.v(280[12] 370[6])
    defparam i15178_4_lut.LUT_INIT = 16'h0032;
    SB_LUT4 i30_4_lut (.I0(n2594), .I1(n17759), .I2(\UART_TRANSMITTER.state [2]), 
            .I3(n5_adj_2407), .O(n13_adj_2437));   // coms.v(280[12] 370[6])
    defparam i30_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i36_4_lut (.I0(\UART_TRANSMITTER.state [1]), .I1(n4_adj_2414), 
            .I2(\UART_TRANSMITTER.state [2]), .I3(\UART_TRANSMITTER.state [0]), 
            .O(n16618));   // coms.v(280[12] 370[6])
    defparam i36_4_lut.LUT_INIT = 16'hb58a;
    SB_LUT4 i24_4_lut_adj_790 (.I0(n18091), .I1(n10_adj_2432), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10_adj_2483));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_4_lut_adj_790.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut_adj_791 (.I0(r_Tx_Data[5]), .I1(n10_adj_2483), .I2(n9257), 
            .I3(byte_transmit_counter[4]), .O(n16912));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i23_4_lut_adj_791.LUT_INIT = 16'h0aca;
    SB_LUT4 i8227_3_lut (.I0(\data_out[0] [1]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n10596), .I3(GND_net), .O(n10913));   // coms.v(280[12] 370[6])
    defparam i8227_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8403_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n9999), 
            .I3(n13116), .O(n11089));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8403_4_lut.LUT_INIT = 16'hcacc;
    SB_LUT4 i8404_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n10010), 
            .I3(n4), .O(n11090));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8404_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8405_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11091));   // coms.v(416[12] 543[6])
    defparam i8405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8406_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11092));   // coms.v(416[12] 543[6])
    defparam i8406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8407_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11093));   // coms.v(416[12] 543[6])
    defparam i8407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8408_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11094));   // coms.v(416[12] 543[6])
    defparam i8408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8409_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11095));   // coms.v(416[12] 543[6])
    defparam i8409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8410_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11096));   // coms.v(416[12] 543[6])
    defparam i8410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8411_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11097));   // coms.v(416[12] 543[6])
    defparam i8411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8412_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11098));   // coms.v(416[12] 543[6])
    defparam i8412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8413_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11099));   // coms.v(416[12] 543[6])
    defparam i8413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8414_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11100));   // coms.v(416[12] 543[6])
    defparam i8414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8415_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11101));   // coms.v(416[12] 543[6])
    defparam i8415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8416_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11102));   // coms.v(416[12] 543[6])
    defparam i8416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8417_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11103));   // coms.v(416[12] 543[6])
    defparam i8417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14574_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n5), 
            .I2(n2061), .I3(GND_net), .O(n17349));
    defparam i14574_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i8418_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11104));   // coms.v(416[12] 543[6])
    defparam i8418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8419_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11105));   // coms.v(416[12] 543[6])
    defparam i8419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8420_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11106));   // coms.v(416[12] 543[6])
    defparam i8420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8421_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11107));   // coms.v(416[12] 543[6])
    defparam i8421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8422_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11108));   // coms.v(416[12] 543[6])
    defparam i8422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8423_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11109));   // coms.v(416[12] 543[6])
    defparam i8423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8424_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11110));   // coms.v(416[12] 543[6])
    defparam i8424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8425_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11111));   // coms.v(416[12] 543[6])
    defparam i8425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8426_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n9999), 
            .I3(n4), .O(n11112));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8426_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8427_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11113));   // coms.v(416[12] 543[6])
    defparam i8427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8428_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11114));   // coms.v(416[12] 543[6])
    defparam i8428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8429_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11115));   // coms.v(416[12] 543[6])
    defparam i8429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8228_3_lut_4_lut (.I0(\data_out[0] [0]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n10596), .O(n10914));   // coms.v(280[12] 370[6])
    defparam i8228_3_lut_4_lut.LUT_INIT = 16'hc0aa;
    SB_LUT4 i8430_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11116));   // coms.v(416[12] 543[6])
    defparam i8430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.i_31__N_1272 ), .I1(n488), .I2(GND_net), 
            .I3(GND_net), .O(n3_adj_2485));   // coms.v(416[12] 543[6])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(n10140), .I1(\FRAME_MATCHER.i_31__N_1275 ), .I2(n4408), 
            .I3(GND_net), .O(n17089));   // coms.v(416[12] 543[6])
    defparam i1_3_lut.LUT_INIT = 16'h5d5d;
    SB_LUT4 i8353_4_lut_4_lut (.I0(r_SM_Main_adj_2503[2]), .I1(n8191), .I2(r_SM_Main_2__N_2031_adj_2510[1]), 
            .I3(r_SM_Main_adj_2503[0]), .O(n11039));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8353_4_lut_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i8352_4_lut_4_lut (.I0(tx2_active), .I1(r_SM_Main_adj_2503[1]), 
            .I2(r_SM_Main_adj_2503[2]), .I3(n4_adj_2484), .O(n11038));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8352_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i8523_3_lut (.I0(\data_out_frame2[12] [4]), .I1(rand_data[4]), 
            .I2(n10725), .I3(GND_net), .O(n11209));   // coms.v(416[12] 543[6])
    defparam i8523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8524_3_lut (.I0(\data_out_frame2[12] [5]), .I1(rand_data[5]), 
            .I2(n10725), .I3(GND_net), .O(n11210));   // coms.v(416[12] 543[6])
    defparam i8524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8431_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11117));   // coms.v(416[12] 543[6])
    defparam i8431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8432_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11118));   // coms.v(416[12] 543[6])
    defparam i8432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8433_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11119));   // coms.v(416[12] 543[6])
    defparam i8433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8434_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11120));   // coms.v(416[12] 543[6])
    defparam i8434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8435_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11121));   // coms.v(416[12] 543[6])
    defparam i8435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8437_3_lut (.I0(\data_out[8] [1]), .I1(rand_setpoint[1]), .I2(data_out_10__7__N_110), 
            .I3(GND_net), .O(n11123));   // coms.v(280[12] 370[6])
    defparam i8437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8438_3_lut (.I0(\data_out[9] [2]), .I1(data_out_9__2__N_367), 
            .I2(data_out_10__7__N_110), .I3(GND_net), .O(n11124));   // coms.v(280[12] 370[6])
    defparam i8438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8439_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11125));   // coms.v(416[12] 543[6])
    defparam i8439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8440_3_lut (.I0(\data_out[8] [7]), .I1(rand_setpoint[7]), .I2(data_out_10__7__N_110), 
            .I3(GND_net), .O(n11126));   // coms.v(280[12] 370[6])
    defparam i8440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8441_3_lut (.I0(\data_out[8] [6]), .I1(rand_setpoint[6]), .I2(data_out_10__7__N_110), 
            .I3(GND_net), .O(n11127));   // coms.v(280[12] 370[6])
    defparam i8441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_792 (.I0(\FRAME_MATCHER.i_31__N_1273 ), .I1(n3779), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2488));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_792.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut (.I0(n17089), .I1(n17349), .I2(n6_adj_2488), .I3(n3_adj_2485), 
            .O(n17090));   // coms.v(416[12] 543[6])
    defparam i2_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_4_lut (.I0(n1_adj_2486), .I1(\FRAME_MATCHER.state [0]), .I2(n17090), 
            .I3(n9378), .O(n16662));   // coms.v(416[12] 543[6])
    defparam i1_4_lut.LUT_INIT = 16'heafa;
    SB_LUT4 i8442_3_lut (.I0(\data_out[8] [5]), .I1(rand_setpoint[5]), .I2(data_out_10__7__N_110), 
            .I3(GND_net), .O(n11128));   // coms.v(280[12] 370[6])
    defparam i8442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8443_3_lut (.I0(\data_out[8] [4]), .I1(rand_setpoint[4]), .I2(data_out_10__7__N_110), 
            .I3(GND_net), .O(n11129));   // coms.v(280[12] 370[6])
    defparam i8443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8444_3_lut (.I0(\data_out[8] [3]), .I1(rand_setpoint[3]), .I2(data_out_10__7__N_110), 
            .I3(GND_net), .O(n11130));   // coms.v(280[12] 370[6])
    defparam i8444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8445_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n11131));   // coms.v(416[12] 543[6])
    defparam i8445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8446_3_lut (.I0(\data_out[8] [2]), .I1(rand_setpoint[2]), .I2(data_out_10__7__N_110), 
            .I3(GND_net), .O(n11132));   // coms.v(280[12] 370[6])
    defparam i8446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_793 (.I0(\FRAME_MATCHER.state [2]), .I1(n63), .I2(n63_adj_2428), 
            .I3(n63_adj_2418), .O(\FRAME_MATCHER.state_31__N_1406 [2]));   // coms.v(416[12] 543[6])
    defparam i1_4_lut_adj_793.LUT_INIT = 16'h8c0c;
    SB_LUT4 i1_4_lut_adj_794 (.I0(n1_adj_2486), .I1(\FRAME_MATCHER.state_31__N_1406 [2]), 
            .I2(\FRAME_MATCHER.i_31__N_1275 ), .I3(n4408), .O(n6));   // coms.v(416[12] 543[6])
    defparam i1_4_lut_adj_794.LUT_INIT = 16'hfaea;
    SB_LUT4 i3_4_lut_adj_795 (.I0(n17349), .I1(n6), .I2(\FRAME_MATCHER.state_31__N_1406 [2]), 
            .I3(n3_adj_2485), .O(n8));   // coms.v(416[12] 543[6])
    defparam i3_4_lut_adj_795.LUT_INIT = 16'hfcdc;
    SB_LUT4 i4_4_lut (.I0(n4_adj_2417), .I1(n8), .I2(\FRAME_MATCHER.state_31__N_1406 [2]), 
            .I3(n10140), .O(n18287));   // coms.v(416[12] 543[6])
    defparam i4_4_lut.LUT_INIT = 16'heefe;
    SB_LUT4 rand_setpoint_2359_add_4_5_lut (.I0(GND_net), .I1(rand_data[3]), 
            .I2(rand_setpoint[3]), .I3(n16012), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2360_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n26_adj_2423), 
            .CO(n16041));
    SB_LUT4 i14639_4_lut (.I0(\UART_TRANSMITTER.state [1]), .I1(n450), .I2(\UART_TRANSMITTER.state [2]), 
            .I3(n4_adj_2414), .O(n17416));
    defparam i14639_4_lut.LUT_INIT = 16'hfaea;
    SB_LUT4 i1_4_lut_adj_796 (.I0(n10088), .I1(n17089), .I2(n3_adj_2485), 
            .I3(n17086), .O(n17063));   // coms.v(416[12] 543[6])
    defparam i1_4_lut_adj_796.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_4_lut_adj_797 (.I0(\FRAME_MATCHER.state [1]), .I1(n9), .I2(n17063), 
            .I3(n31_adj_2415), .O(n21_adj_2487));   // coms.v(416[12] 543[6])
    defparam i1_4_lut_adj_797.LUT_INIT = 16'ha0a2;
    SB_LUT4 i15147_4_lut (.I0(n4_adj_2414), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [2]), .I3(n4_adj_2419), .O(n17765));   // coms.v(280[12] 370[6])
    defparam i15147_4_lut.LUT_INIT = 16'hece0;
    SB_LUT4 i8525_3_lut (.I0(\data_out_frame2[12] [6]), .I1(rand_data[6]), 
            .I2(n10725), .I3(GND_net), .O(n11211));   // coms.v(416[12] 543[6])
    defparam i8525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8211_3_lut_4_lut (.I0(\data_out[3] [5]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n10596), .O(n10897));   // coms.v(280[12] 370[6])
    defparam i8211_3_lut_4_lut.LUT_INIT = 16'hc0aa;
    SB_LUT4 i8526_3_lut (.I0(\data_out_frame2[12] [7]), .I1(rand_data[7]), 
            .I2(n10725), .I3(GND_net), .O(n11212));   // coms.v(416[12] 543[6])
    defparam i8526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_798 (.I0(\FRAME_MATCHER.i_31__N_1273 ), .I1(n63_adj_2418), 
            .I2(n3779), .I3(n17063), .O(n6_adj_2410));   // coms.v(416[12] 543[6])
    defparam i2_4_lut_adj_798.LUT_INIT = 16'hb3a0;
    SB_LUT4 i8527_3_lut (.I0(\data_out_frame2[13] [0]), .I1(rand_data[24]), 
            .I2(n10725), .I3(GND_net), .O(n11213));   // coms.v(416[12] 543[6])
    defparam i8527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_799 (.I0(n44), .I1(n6_adj_2410), .I2(n21_adj_2487), 
            .I3(n2061), .O(n18286));   // coms.v(416[12] 543[6])
    defparam i3_4_lut_adj_799.LUT_INIT = 16'hfdfc;
    SB_LUT4 i8528_3_lut (.I0(\data_out_frame2[13] [1]), .I1(rand_data[25]), 
            .I2(n10725), .I3(GND_net), .O(n11214));   // coms.v(416[12] 543[6])
    defparam i8528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8529_3_lut (.I0(\data_out_frame2[13] [2]), .I1(rand_data[26]), 
            .I2(n10725), .I3(GND_net), .O(n11215));   // coms.v(416[12] 543[6])
    defparam i8529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43_4_lut (.I0(n17392), .I1(n17765), .I2(\UART_TRANSMITTER.state [0]), 
            .I3(n17416), .O(n16614));   // coms.v(280[12] 370[6])
    defparam i43_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i8530_3_lut (.I0(\data_out_frame2[13] [3]), .I1(rand_data[27]), 
            .I2(n10725), .I3(GND_net), .O(n11216));   // coms.v(416[12] 543[6])
    defparam i8530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8212_3_lut (.I0(\data_out[3] [4]), .I1(n2699), .I2(n10596), 
            .I3(GND_net), .O(n10898));   // coms.v(280[12] 370[6])
    defparam i8212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8531_3_lut (.I0(\data_out_frame2[13] [4]), .I1(rand_data[28]), 
            .I2(n10725), .I3(GND_net), .O(n11217));   // coms.v(416[12] 543[6])
    defparam i8531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8213_3_lut (.I0(\data_out[3] [2]), .I1(n2699), .I2(n10596), 
            .I3(GND_net), .O(n10899));   // coms.v(280[12] 370[6])
    defparam i8213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14651_4_lut (.I0(blink_counter[22]), .I1(blink_counter[23]), 
            .I2(blink_counter[24]), .I3(blink_counter[21]), .O(n17428));
    defparam i14651_4_lut.LUT_INIT = 16'hfec4;
    SB_LUT4 i14650_4_lut (.I0(blink_counter[23]), .I1(blink_counter[22]), 
            .I2(blink_counter[24]), .I3(blink_counter[21]), .O(n17427));
    defparam i14650_4_lut.LUT_INIT = 16'hcf08;
    SB_LUT4 i14652_3_lut (.I0(n17427), .I1(n17428), .I2(blink_counter[25]), 
            .I3(GND_net), .O(LED_c));
    defparam i14652_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i8209_3_lut_4_lut (.I0(\data_out[3] [7]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n10596), .O(n10895));   // coms.v(280[12] 370[6])
    defparam i8209_3_lut_4_lut.LUT_INIT = 16'hc0aa;
    SB_LUT4 i8532_3_lut (.I0(\data_out_frame2[13] [5]), .I1(rand_data[29]), 
            .I2(n10725), .I3(GND_net), .O(n11218));   // coms.v(416[12] 543[6])
    defparam i8532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8214_3_lut (.I0(\data_out[3] [0]), .I1(n2699), .I2(n10596), 
            .I3(GND_net), .O(n10900));   // coms.v(280[12] 370[6])
    defparam i8214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8533_3_lut (.I0(\data_out_frame2[13] [6]), .I1(rand_data[30]), 
            .I2(n10725), .I3(GND_net), .O(n11219));   // coms.v(416[12] 543[6])
    defparam i8533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8215_3_lut (.I0(\data_out[2] [7]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n10596), .I3(GND_net), .O(n10901));   // coms.v(280[12] 370[6])
    defparam i8215_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8534_3_lut (.I0(\data_out_frame2[13] [7]), .I1(rand_data[31]), 
            .I2(n10725), .I3(GND_net), .O(n11220));   // coms.v(416[12] 543[6])
    defparam i8534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8535_3_lut (.I0(\data_out_frame2[14] [0]), .I1(rand_data[16]), 
            .I2(n10725), .I3(GND_net), .O(n11221));   // coms.v(416[12] 543[6])
    defparam i8535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8536_3_lut (.I0(\data_out_frame2[14] [1]), .I1(rand_data[17]), 
            .I2(n10725), .I3(GND_net), .O(n11222));   // coms.v(416[12] 543[6])
    defparam i8536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8537_3_lut (.I0(\data_out_frame2[14] [2]), .I1(rand_data[18]), 
            .I2(n10725), .I3(GND_net), .O(n11223));   // coms.v(416[12] 543[6])
    defparam i8537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8538_3_lut (.I0(\data_out_frame2[14] [3]), .I1(rand_data[19]), 
            .I2(n10725), .I3(GND_net), .O(n11224));   // coms.v(416[12] 543[6])
    defparam i8538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8539_3_lut (.I0(\data_out_frame2[14] [4]), .I1(rand_data[20]), 
            .I2(n10725), .I3(GND_net), .O(n11225));   // coms.v(416[12] 543[6])
    defparam i8539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8540_3_lut (.I0(\data_out_frame2[14] [5]), .I1(rand_data[21]), 
            .I2(n10725), .I3(GND_net), .O(n11226));   // coms.v(416[12] 543[6])
    defparam i8540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8541_3_lut (.I0(\data_out_frame2[14] [6]), .I1(rand_data[22]), 
            .I2(n10725), .I3(GND_net), .O(n11227));   // coms.v(416[12] 543[6])
    defparam i8541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8542_3_lut (.I0(\data_out_frame2[14] [7]), .I1(rand_data[23]), 
            .I2(n10725), .I3(GND_net), .O(n11228));   // coms.v(416[12] 543[6])
    defparam i8542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2359_add_4_33_lut (.I0(GND_net), .I1(rand_data[31]), 
            .I2(rand_setpoint[31]), .I3(n16040), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2359_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8543_3_lut (.I0(\data_out_frame2[15] [0]), .I1(rand_data[8]), 
            .I2(n10725), .I3(GND_net), .O(n11229));   // coms.v(416[12] 543[6])
    defparam i8543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8544_3_lut (.I0(\data_out_frame2[15] [1]), .I1(rand_data[9]), 
            .I2(n10725), .I3(GND_net), .O(n11230));   // coms.v(416[12] 543[6])
    defparam i8544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8545_3_lut (.I0(\data_out_frame2[15] [2]), .I1(rand_data[10]), 
            .I2(n10725), .I3(GND_net), .O(n11231));   // coms.v(416[12] 543[6])
    defparam i8545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8546_3_lut (.I0(\data_out_frame2[15] [3]), .I1(rand_data[11]), 
            .I2(n10725), .I3(GND_net), .O(n11232));   // coms.v(416[12] 543[6])
    defparam i8546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8547_3_lut (.I0(\data_out_frame2[15] [4]), .I1(rand_data[12]), 
            .I2(n10725), .I3(GND_net), .O(n11233));   // coms.v(416[12] 543[6])
    defparam i8547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8548_3_lut (.I0(\data_out_frame2[15] [5]), .I1(rand_data[13]), 
            .I2(n10725), .I3(GND_net), .O(n11234));   // coms.v(416[12] 543[6])
    defparam i8548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8549_3_lut (.I0(\data_out_frame2[15] [6]), .I1(rand_data[14]), 
            .I2(n10725), .I3(GND_net), .O(n11235));   // coms.v(416[12] 543[6])
    defparam i8549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8550_3_lut (.I0(\data_out_frame2[15] [7]), .I1(rand_data[15]), 
            .I2(n10725), .I3(GND_net), .O(n11236));   // coms.v(416[12] 543[6])
    defparam i8550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8551_3_lut (.I0(\data_out_frame2[16] [0]), .I1(rand_data[0]), 
            .I2(n10725), .I3(GND_net), .O(n11237));   // coms.v(416[12] 543[6])
    defparam i8551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8552_3_lut (.I0(\data_out_frame2[16] [1]), .I1(rand_data[1]), 
            .I2(n10725), .I3(GND_net), .O(n11238));   // coms.v(416[12] 543[6])
    defparam i8552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8553_3_lut (.I0(\data_out_frame2[16] [2]), .I1(rand_data[2]), 
            .I2(n10725), .I3(GND_net), .O(n11239));   // coms.v(416[12] 543[6])
    defparam i8553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8554_3_lut (.I0(\data_out_frame2[16] [3]), .I1(rand_data[3]), 
            .I2(n10725), .I3(GND_net), .O(n11240));   // coms.v(416[12] 543[6])
    defparam i8554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8555_3_lut (.I0(\data_out_frame2[16] [4]), .I1(rand_data[4]), 
            .I2(n10725), .I3(GND_net), .O(n11241));   // coms.v(416[12] 543[6])
    defparam i8555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8556_3_lut (.I0(\data_out_frame2[16] [5]), .I1(rand_data[5]), 
            .I2(n10725), .I3(GND_net), .O(n11242));   // coms.v(416[12] 543[6])
    defparam i8556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8557_3_lut (.I0(\data_out_frame2[16] [6]), .I1(rand_data[6]), 
            .I2(n10725), .I3(GND_net), .O(n11243));   // coms.v(416[12] 543[6])
    defparam i8557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8216_3_lut (.I0(\data_out[2] [5]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n10596), .I3(GND_net), .O(n10902));   // coms.v(280[12] 370[6])
    defparam i8216_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8558_3_lut (.I0(\data_out_frame2[16] [7]), .I1(rand_data[7]), 
            .I2(n10725), .I3(GND_net), .O(n11244));   // coms.v(416[12] 543[6])
    defparam i8558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8559_3_lut (.I0(\data_out_frame2[17] [0]), .I1(rand_data[8]), 
            .I2(n10725), .I3(GND_net), .O(n11245));   // coms.v(416[12] 543[6])
    defparam i8559_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 i8218_3_lut (.I0(\data_out[2] [2]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n10596), .I3(GND_net), .O(n10904));   // coms.v(280[12] 370[6])
    defparam i8218_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8219_3_lut (.I0(\data_out[2] [0]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n10596), .I3(GND_net), .O(n10905));   // coms.v(280[12] 370[6])
    defparam i8219_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8220_3_lut (.I0(\data_out[1] [7]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n10596), .I3(GND_net), .O(n10906));   // coms.v(280[12] 370[6])
    defparam i8220_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8560_3_lut (.I0(\data_out_frame2[17] [1]), .I1(rand_data[9]), 
            .I2(n10725), .I3(GND_net), .O(n11246));   // coms.v(416[12] 543[6])
    defparam i8560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8449_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n10010), 
            .I3(n4_adj_2427), .O(n11135));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8449_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8450_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n9999), 
            .I3(n4_adj_2427), .O(n11136));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8450_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8561_3_lut (.I0(\data_out_frame2[17] [2]), .I1(rand_data[10]), 
            .I2(n10725), .I3(GND_net), .O(n11247));   // coms.v(416[12] 543[6])
    defparam i8561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15221_4_lut (.I0(r_SM_Main_adj_2500[2]), .I1(n17707), .I2(n17708), 
            .I3(r_SM_Main_adj_2500[1]), .O(n13744));
    defparam i15221_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i8562_3_lut (.I0(\data_out_frame2[17] [3]), .I1(rand_data[11]), 
            .I2(n10725), .I3(GND_net), .O(n11248));   // coms.v(416[12] 543[6])
    defparam i8562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8453_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n10010), 
            .I3(n4_adj_2416), .O(n11139));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8453_4_lut.LUT_INIT = 16'hccca;
    coms c0 (.tx_transmit_N_1947({tx_transmit_N_1947}), .\UART_TRANSMITTER.state[1] (\UART_TRANSMITTER.state [1]), 
         .\UART_TRANSMITTER.state[2] (\UART_TRANSMITTER.state [2]), .byte_transmit_counter({byte_transmit_counter}), 
         .\FRAME_MATCHER.i_31__N_1273 (\FRAME_MATCHER.i_31__N_1273 ), .n3779(n3779), 
         .GND_net(GND_net), .n444(n444), .\UART_TRANSMITTER.state[0] (\UART_TRANSMITTER.state [0]), 
         .n2061(n2061), .n18175(n18175), .n4408(n4408), .\FRAME_MATCHER.i_31__N_1275 (\FRAME_MATCHER.i_31__N_1275 ), 
         .\data_out_frame2[9] ({\data_out_frame2[9] }), .\data_out_frame2[8] ({\data_out_frame2[8] }), 
         .\data_out_frame2[18] ({\data_out_frame2[18] }), .\data_out_frame2[17] ({\data_out_frame2[17] }), 
         .\data_out_frame2[16] ({\data_out_frame2[16] }), .n2593({n2594}), 
         .\rand_setpoint[15] (rand_setpoint[15]), .n18271(n18271), .\data_out_frame2[6] ({\data_out_frame2[6] }), 
         .\data_out_frame2[7] ({\data_out_frame2[7] }), .\data_out_frame2[5] ({\data_out_frame2[5] }), 
         .\data_out_frame2[14] ({\data_out_frame2[14] }), .\data_out_frame2[15] ({\data_out_frame2[15] }), 
         .\data_out[8] ({\data_out[8] [7], Open_0, Open_1, Open_2, Open_3, 
         Open_4, Open_5, Open_6}), .n10(n10_adj_2413), .\data_out[1][7] (\data_out[1] [7]), 
         .\rand_setpoint[16] (rand_setpoint[16]), .n10596(n10596), .\rand_setpoint[31] (rand_setpoint[31]), 
         .\data_out_frame2[13] ({\data_out_frame2[13] }), .\data_out_frame2[12] ({\data_out_frame2[12] }), 
         .n8(n8_adj_2445), .n18169(n18169), .CLK_c(CLK_c), .\data_out[2][0] (\data_out[2] [0]), 
         .\data_out[3][0] (\data_out[3] [0]), .n2(n2), .n6(n6_adj_2446), 
         .n18223(n18223), .\data_out[2][7] (\data_out[2] [7]), .\data_out[3][7] (\data_out[3] [7]), 
         .\data_out[8][6] (\data_out[8] [6]), .\rand_setpoint[12] (rand_setpoint[12]), 
         .\rand_setpoint[30] (rand_setpoint[30]), .n10_adj_3(n10_adj_2422), 
         .\FRAME_MATCHER.i_31__N_1272 (\FRAME_MATCHER.i_31__N_1272 ), .\data_out_frame2[10] ({\data_out_frame2[10] }), 
         .\data_out_frame2[11] ({\data_out_frame2[11] }), .\data_out[5][1] (\data_out[5] [1]), 
         .n16614(n16614), .n16662(n16662), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n10914(n10914), .\data_out[0][0] (\data_out[0] [0]), .n10913(n10913), 
         .\data_out[0][1] (\data_out[0] [1]), .\rand_setpoint[29] (rand_setpoint[29]), 
         .n18187(n18187), .\rand_setpoint[28] (rand_setpoint[28]), .n10912(n10912), 
         .\data_out[0][3] (\data_out[0] [3]), .\rand_setpoint[27] (rand_setpoint[27]), 
         .\rand_setpoint[26] (rand_setpoint[26]), .\rand_setpoint[24] (rand_setpoint[24]), 
         .\FRAME_MATCHER.state[2] (\FRAME_MATCHER.state [2]), .\FRAME_MATCHER.state[1] (\FRAME_MATCHER.state [1]), 
         .\rand_setpoint[13] (rand_setpoint[13]), .\rand_setpoint[14] (rand_setpoint[14]), 
         .n10911(n10911), .\data_out[0][5] (\data_out[0] [5]), .n5(n5_adj_2448), 
         .\data_out[8][5] (\data_out[8] [5]), .n18091(n18091), .n16634(n16634), 
         .n16632(n16632), .n16630(n16630), .\data_out[8][3] (\data_out[8] [3]), 
         .\data_out[8][4] (\data_out[8] [4]), .n16628(n16628), .\data_out[8][1] (\data_out[8] [1]), 
         .n8_adj_4(n8_adj_2447), .n1(n1_adj_2449), .n16626(n16626), .n16624(n16624), 
         .n16622(n16622), .n16620(n16620), .n11260(n11260), .\data_out[9][2] (\data_out[9] [2]), 
         .n11259(n11259), .n11258(n11258), .n11257(n11257), .n11256(n11256), 
         .\data_out[8][2] (\data_out[8] [2]), .n10_adj_5(n10_adj_2450), 
         .n11255(n11255), .n11254(n11254), .n11253(n11253), .n11252(n11252), 
         .n11251(n11251), .n11250(n11250), .n11249(n11249), .n11248(n11248), 
         .n11247(n11247), .n10907(n10907), .\data_out[1][6] (\data_out[1] [6]), 
         .data_out_9__2__N_367(data_out_9__2__N_367), .\data_out[10][1] (\data_out[10] [1]), 
         .n11246(n11246), .n10906(n10906), .n10905(n10905), .n10_adj_6(n10_adj_2431), 
         .n10904(n10904), .\data_out[2][2] (\data_out[2] [2]), .n11245(n11245), 
         .n11244(n11244), .n10902(n10902), .\data_out[2][5] (\data_out[2] [5]), 
         .n11243(n11243), .n11242(n11242), .n11241(n11241), .n11240(n11240), 
         .n10_adj_7(n10_adj_2430), .n11239(n11239), .n11238(n11238), .n11237(n11237), 
         .n11236(n11236), .n11235(n11235), .n11234(n11234), .n11233(n11233), 
         .n11232(n11232), .n11231(n11231), .n11230(n11230), .n11229(n11229), 
         .n11228(n11228), .\data_out[3][2] (\data_out[3] [2]), .VCC_net(VCC_net), 
         .rx_data({rx_data}), .n11227(n11227), .n11226(n11226), .n11225(n11225), 
         .n11224(n11224), .n11223(n11223), .n11222(n11222), .n11221(n11221), 
         .n11220(n11220), .n10901(n10901), .n11219(n11219), .n10900(n10900), 
         .n11218(n11218), .n10899(n10899), .n11217(n11217), .n10705(n10705), 
         .n10898(n10898), .\data_out[3][4] (\data_out[3] [4]), .n11216(n11216), 
         .n11215(n11215), .n11214(n11214), .n11213(n11213), .n11212(n11212), 
         .n31(n31_adj_2415), .n11211(n11211), .n11210(n11210), .n11209(n11209), 
         .n11208(n11208), .n11207(n11207), .n11206(n11206), .n11205(n11205), 
         .n11204(n11204), .\data_out[3][5] (\data_out[3] [5]), .n11203(n11203), 
         .n11202(n11202), .n11201(n11201), .n11200(n11200), .n11199(n11199), 
         .n11198(n11198), .n11197(n11197), .n11196(n11196), .n11195(n11195), 
         .n11194(n11194), .n11193(n11193), .n11192(n11192), .n11191(n11191), 
         .n11190(n11190), .n11189(n11189), .tx2_active(tx2_active), .n11188(n11188), 
         .n11187(n11187), .n11186(n11186), .n10897(n10897), .n10895(n10895), 
         .n11185(n11185), .n488(n488), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .n11184(n11184), .n11183(n11183), .n11182(n11182), .n11181(n11181), 
         .n11180(n11180), .n11179(n11179), .n11178(n11178), .data_out_10__7__N_110(data_out_10__7__N_110), 
         .\data_out[10][0] (\data_out[10] [0]), .n2698({n2699}), .n11177(n11177), 
         .n11176(n11176), .n11175(n11175), .n11174(n11174), .n11173(n11173), 
         .n11172(n11172), .n11171(n11171), .n11170(n11170), .n11169(n11169), 
         .n11168(n11168), .n11167(n11167), .n11166(n11166), .n11165(n11165), 
         .n11164(n11164), .n11163(n11163), .n11162(n11162), .n11161(n11161), 
         .n11160(n11160), .n11159(n11159), .n11158(n11158), .n11157(n11157), 
         .n11156(n11156), .n11155(n11155), .n11154(n11154), .n11153(n11153), 
         .n11152(n11152), .n11151(n11151), .n11150(n11150), .n11149(n11149), 
         .n18286(n18286), .n18287(n18287), .n17392(n17392), .n4(n4_adj_2419), 
         .n11132(n11132), .n11131(n11131), .\data_in[3] ({\data_in[3] }), 
         .n11130(n11130), .n11129(n11129), .n11128(n11128), .n11127(n11127), 
         .n11126(n11126), .n11125(n11125), .n11124(n11124), .n11123(n11123), 
         .n11121(n11121), .n11120(n11120), .n17075(n17075), .n9378(n9378), 
         .n11119(n11119), .n11118(n11118), .n5_adj_8(n5), .n17086(n17086), 
         .n9(n9), .n63(n63_adj_2418), .n63_adj_9(n63_adj_2428), .n63_adj_10(n63), 
         .n11117(n11117), .n11116(n11116), .n11115(n11115), .\data_in[2] ({\data_in[2] }), 
         .n10_adj_11(n10_adj_2432), .n11114(n11114), .n11113(n11113), 
         .n11111(n11111), .n11110(n11110), .n11109(n11109), .n10088(n10088), 
         .n11108(n11108), .n11107(n11107), .\data_in[0] ({\data_in[0] }), 
         .\data_in[1] ({\data_in[1] }), .n11106(n11106), .n44(n44), .n11105(n11105), 
         .n10140(n10140), .n11104(n11104), .n11103(n11103), .n11102(n11102), 
         .n11101(n11101), .n11100(n11100), .n11099(n11099), .n11098(n11098), 
         .n11097(n11097), .n11096(n11096), .n11095(n11095), .n11094(n11094), 
         .n11093(n11093), .n11092(n11092), .n11091(n11091), .n1_adj_12(n1_adj_2486), 
         .n10725(n10725), .n16618(n16618), .n13(n13_adj_2437), .\rand_setpoint[0] (rand_setpoint[0]), 
         .n9524(n9524), .n450(n450), .\FRAME_MATCHER.state_31__N_1406[2] (\FRAME_MATCHER.state_31__N_1406 [2]), 
         .n4_adj_13(n4_adj_2417), .n4_adj_14(n4_adj_2414), .n11033(n11033), 
         .n11032(n11032), .n11028(n11028), .\rand_setpoint[25] (rand_setpoint[25]), 
         .\rand_setpoint[17] (rand_setpoint[17]), .n11027(n11027), .n11025(n11025), 
         .\rand_setpoint[18] (rand_setpoint[18]), .n11024(n11024), .n11023(n11023), 
         .\rand_setpoint[19] (rand_setpoint[19]), .n11016(n11016), .\rand_setpoint[20] (rand_setpoint[20]), 
         .\rand_setpoint[21] (rand_setpoint[21]), .\rand_setpoint[22] (rand_setpoint[22]), 
         .\rand_setpoint[23] (rand_setpoint[23]), .\rand_setpoint[8] (rand_setpoint[8]), 
         .n17327(n17327), .rx_data_ready(rx_data_ready), .\rand_setpoint[9] (rand_setpoint[9]), 
         .\rand_setpoint[10] (rand_setpoint[10]), .\rand_setpoint[11] (rand_setpoint[11]), 
         .n10969(n10969), .n10966(n10966), .n10963(n10963), .n10960(n10960), 
         .n10957(n10957), .n10954(n10954), .n10951(n10951), .n10994(n10994), 
         .\r_Bit_Index[2] (r_Bit_Index[2]), .n16932(n16932), .r_Tx_Data({r_Tx_Data}), 
         .n16930(n16930), .n16928(n16928), .n16926(n16926), .\r_Bit_Index[1] (r_Bit_Index[1]), 
         .n10953(n10953), .n10956(n10956), .n10959(n10959), .n10962(n10962), 
         .n10965(n10965), .n10968(n10968), .n10971(n10971), .n10974(n10974), 
         .n16924(n16924), .n10996(n10996), .n16914(n16914), .n16902(n16902), 
         .n18199(n18199), .n18073(n18073), .tx_o(tx_o), .n9257(n9257), 
         .n16912(n16912), .n5142(n5142), .n10972(n10972), .tx_enable(tx_enable), 
         .\r_SM_Main_2__N_2031[1] (r_SM_Main_2__N_2031_adj_2510[1]), .r_SM_Main({r_SM_Main_adj_2503}), 
         .n4_adj_15(n4_adj_2484), .r_Bit_Index({r_Bit_Index_adj_2505}), 
         .n18280(n18280), .n10674(n10674), .n10920(n10920), .n10923(n10923), 
         .n10977(n10977), .n5266(n5266), .n17412(n17412), .n10976(n10976), 
         .n3(n3), .n8191(n8191), .n11039(n11039), .n11038(n11038), .n11037(n11037), 
         .tx2_o(tx2_o), .tx2_enable(tx2_enable), .r_Bit_Index_adj_27({r_Bit_Index_adj_2499}), 
         .n5244(n5244), .\r_SM_Main[1]_adj_21 (r_SM_Main_adj_2500[1]), .\r_SM_Main[2]_adj_22 (r_SM_Main_adj_2500[2]), 
         .n17361(n17361), .n10983(n10983), .n11019(n11019), .n11031(n11031), 
         .r_Rx_Data(r_Rx_Data), .rx_i(rx_i), .n11139(n11139), .n13744(n13744), 
         .n11136(n11136), .n11135(n11135), .n1_adj_23(n1), .n13116(n13116), 
         .n11112(n11112), .n4_adj_24(n4), .n11090(n11090), .n11089(n11089), 
         .n11034(n11034), .n11026(n11026), .n10987(n10987), .n13692(n13692), 
         .n11018(n11018), .n4_adj_25(n4_adj_2427), .n9999(n9999), .n17708(n17708), 
         .n17707(n17707), .n4_adj_26(n4_adj_2416), .n10010(n10010)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(84[8] 97[4])
    SB_LUT4 i8563_3_lut (.I0(\data_out_frame2[17] [4]), .I1(rand_data[12]), 
            .I2(n10725), .I3(GND_net), .O(n11249));   // coms.v(416[12] 543[6])
    defparam i8563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8564_3_lut (.I0(\data_out_frame2[17] [5]), .I1(rand_data[13]), 
            .I2(n10725), .I3(GND_net), .O(n11250));   // coms.v(416[12] 543[6])
    defparam i8564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8565_3_lut (.I0(\data_out_frame2[17] [6]), .I1(rand_data[14]), 
            .I2(n10725), .I3(GND_net), .O(n11251));   // coms.v(416[12] 543[6])
    defparam i8565_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module coms
//

module coms (tx_transmit_N_1947, \UART_TRANSMITTER.state[1] , \UART_TRANSMITTER.state[2] , 
            byte_transmit_counter, \FRAME_MATCHER.i_31__N_1273 , n3779, 
            GND_net, n444, \UART_TRANSMITTER.state[0] , n2061, n18175, 
            n4408, \FRAME_MATCHER.i_31__N_1275 , \data_out_frame2[9] , 
            \data_out_frame2[8] , \data_out_frame2[18] , \data_out_frame2[17] , 
            \data_out_frame2[16] , n2593, \rand_setpoint[15] , n18271, 
            \data_out_frame2[6] , \data_out_frame2[7] , \data_out_frame2[5] , 
            \data_out_frame2[14] , \data_out_frame2[15] , \data_out[8] , 
            n10, \data_out[1][7] , \rand_setpoint[16] , n10596, \rand_setpoint[31] , 
            \data_out_frame2[13] , \data_out_frame2[12] , n8, n18169, 
            CLK_c, \data_out[2][0] , \data_out[3][0] , n2, n6, n18223, 
            \data_out[2][7] , \data_out[3][7] , \data_out[8][6] , \rand_setpoint[12] , 
            \rand_setpoint[30] , n10_adj_3, \FRAME_MATCHER.i_31__N_1272 , 
            \data_out_frame2[10] , \data_out_frame2[11] , \data_out[5][1] , 
            n16614, n16662, \FRAME_MATCHER.state[0] , n10914, \data_out[0][0] , 
            n10913, \data_out[0][1] , \rand_setpoint[29] , n18187, \rand_setpoint[28] , 
            n10912, \data_out[0][3] , \rand_setpoint[27] , \rand_setpoint[26] , 
            \rand_setpoint[24] , \FRAME_MATCHER.state[2] , \FRAME_MATCHER.state[1] , 
            \rand_setpoint[13] , \rand_setpoint[14] , n10911, \data_out[0][5] , 
            n5, \data_out[8][5] , n18091, n16634, n16632, n16630, 
            \data_out[8][3] , \data_out[8][4] , n16628, \data_out[8][1] , 
            n8_adj_4, n1, n16626, n16624, n16622, n16620, n11260, 
            \data_out[9][2] , n11259, n11258, n11257, n11256, \data_out[8][2] , 
            n10_adj_5, n11255, n11254, n11253, n11252, n11251, n11250, 
            n11249, n11248, n11247, n10907, \data_out[1][6] , data_out_9__2__N_367, 
            \data_out[10][1] , n11246, n10906, n10905, n10_adj_6, 
            n10904, \data_out[2][2] , n11245, n11244, n10902, \data_out[2][5] , 
            n11243, n11242, n11241, n11240, n10_adj_7, n11239, n11238, 
            n11237, n11236, n11235, n11234, n11233, n11232, n11231, 
            n11230, n11229, n11228, \data_out[3][2] , VCC_net, rx_data, 
            n11227, n11226, n11225, n11224, n11223, n11222, n11221, 
            n11220, n10901, n11219, n10900, n11218, n10899, n11217, 
            n10705, n10898, \data_out[3][4] , n11216, n11215, n11214, 
            n11213, n11212, n31, n11211, n11210, n11209, n11208, 
            n11207, n11206, n11205, n11204, \data_out[3][5] , n11203, 
            n11202, n11201, n11200, n11199, n11198, n11197, n11196, 
            n11195, n11194, n11193, n11192, n11191, n11190, n11189, 
            tx2_active, n11188, n11187, n11186, n10897, n10895, 
            n11185, n488, \data_in_frame[6] , n11184, n11183, n11182, 
            n11181, n11180, n11179, n11178, data_out_10__7__N_110, 
            \data_out[10][0] , n2698, n11177, n11176, n11175, n11174, 
            n11173, n11172, n11171, n11170, n11169, n11168, n11167, 
            n11166, n11165, n11164, n11163, n11162, n11161, n11160, 
            n11159, n11158, n11157, n11156, n11155, n11154, n11153, 
            n11152, n11151, n11150, n11149, n18286, n18287, n17392, 
            n4, n11132, n11131, \data_in[3] , n11130, n11129, n11128, 
            n11127, n11126, n11125, n11124, n11123, n11121, n11120, 
            n17075, n9378, n11119, n11118, n5_adj_8, n17086, n9, 
            n63, n63_adj_9, n63_adj_10, n11117, n11116, n11115, 
            \data_in[2] , n10_adj_11, n11114, n11113, n11111, n11110, 
            n11109, n10088, n11108, n11107, \data_in[0] , \data_in[1] , 
            n11106, n44, n11105, n10140, n11104, n11103, n11102, 
            n11101, n11100, n11099, n11098, n11097, n11096, n11095, 
            n11094, n11093, n11092, n11091, n1_adj_12, n10725, n16618, 
            n13, \rand_setpoint[0] , n9524, n450, \FRAME_MATCHER.state_31__N_1406[2] , 
            n4_adj_13, n4_adj_14, n11033, n11032, n11028, \rand_setpoint[25] , 
            \rand_setpoint[17] , n11027, n11025, \rand_setpoint[18] , 
            n11024, n11023, \rand_setpoint[19] , n11016, \rand_setpoint[20] , 
            \rand_setpoint[21] , \rand_setpoint[22] , \rand_setpoint[23] , 
            \rand_setpoint[8] , n17327, rx_data_ready, \rand_setpoint[9] , 
            \rand_setpoint[10] , \rand_setpoint[11] , n10969, n10966, 
            n10963, n10960, n10957, n10954, n10951, n10994, \r_Bit_Index[2] , 
            n16932, r_Tx_Data, n16930, n16928, n16926, \r_Bit_Index[1] , 
            n10953, n10956, n10959, n10962, n10965, n10968, n10971, 
            n10974, n16924, n10996, n16914, n16902, n18199, n18073, 
            tx_o, n9257, n16912, n5142, n10972, tx_enable, \r_SM_Main_2__N_2031[1] , 
            r_SM_Main, n4_adj_15, r_Bit_Index, n18280, n10674, n10920, 
            n10923, n10977, n5266, n17412, n10976, n3, n8191, 
            n11039, n11038, n11037, tx2_o, tx2_enable, r_Bit_Index_adj_27, 
            n5244, \r_SM_Main[1]_adj_21 , \r_SM_Main[2]_adj_22 , n17361, 
            n10983, n11019, n11031, r_Rx_Data, rx_i, n11139, n13744, 
            n11136, n11135, n1_adj_23, n13116, n11112, n4_adj_24, 
            n11090, n11089, n11034, n11026, n10987, n13692, n11018, 
            n4_adj_25, n9999, n17708, n17707, n4_adj_26, n10010) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [7:0]tx_transmit_N_1947;
    output \UART_TRANSMITTER.state[1] ;
    output \UART_TRANSMITTER.state[2] ;
    output [7:0]byte_transmit_counter;
    output \FRAME_MATCHER.i_31__N_1273 ;
    output n3779;
    input GND_net;
    output n444;
    output \UART_TRANSMITTER.state[0] ;
    output n2061;
    output n18175;
    output n4408;
    output \FRAME_MATCHER.i_31__N_1275 ;
    output [7:0]\data_out_frame2[9] ;
    output [7:0]\data_out_frame2[8] ;
    output [7:0]\data_out_frame2[18] ;
    output [7:0]\data_out_frame2[17] ;
    output [7:0]\data_out_frame2[16] ;
    output [0:0]n2593;
    input \rand_setpoint[15] ;
    output n18271;
    output [7:0]\data_out_frame2[6] ;
    output [7:0]\data_out_frame2[7] ;
    output [7:0]\data_out_frame2[5] ;
    output [7:0]\data_out_frame2[14] ;
    output [7:0]\data_out_frame2[15] ;
    output [7:0]\data_out[8] ;
    output n10;
    output \data_out[1][7] ;
    input \rand_setpoint[16] ;
    output n10596;
    input \rand_setpoint[31] ;
    output [7:0]\data_out_frame2[13] ;
    output [7:0]\data_out_frame2[12] ;
    output n8;
    output n18169;
    input CLK_c;
    output \data_out[2][0] ;
    output \data_out[3][0] ;
    output n2;
    output n6;
    output n18223;
    output \data_out[2][7] ;
    output \data_out[3][7] ;
    output \data_out[8][6] ;
    input \rand_setpoint[12] ;
    input \rand_setpoint[30] ;
    output n10_adj_3;
    output \FRAME_MATCHER.i_31__N_1272 ;
    output [7:0]\data_out_frame2[10] ;
    output [7:0]\data_out_frame2[11] ;
    output \data_out[5][1] ;
    input n16614;
    input n16662;
    output \FRAME_MATCHER.state[0] ;
    input n10914;
    output \data_out[0][0] ;
    input n10913;
    output \data_out[0][1] ;
    input \rand_setpoint[29] ;
    output n18187;
    input \rand_setpoint[28] ;
    input n10912;
    output \data_out[0][3] ;
    input \rand_setpoint[27] ;
    input \rand_setpoint[26] ;
    input \rand_setpoint[24] ;
    output \FRAME_MATCHER.state[2] ;
    output \FRAME_MATCHER.state[1] ;
    input \rand_setpoint[13] ;
    input \rand_setpoint[14] ;
    input n10911;
    output \data_out[0][5] ;
    output n5;
    output \data_out[8][5] ;
    output n18091;
    input n16634;
    input n16632;
    input n16630;
    output \data_out[8][3] ;
    output \data_out[8][4] ;
    input n16628;
    output \data_out[8][1] ;
    output n8_adj_4;
    output n1;
    input n16626;
    input n16624;
    input n16622;
    input n16620;
    input n11260;
    output \data_out[9][2] ;
    input n11259;
    input n11258;
    input n11257;
    input n11256;
    output \data_out[8][2] ;
    output n10_adj_5;
    input n11255;
    input n11254;
    input n11253;
    input n11252;
    input n11251;
    input n11250;
    input n11249;
    input n11248;
    input n11247;
    input n10907;
    output \data_out[1][6] ;
    output data_out_9__2__N_367;
    output \data_out[10][1] ;
    input n11246;
    input n10906;
    input n10905;
    output n10_adj_6;
    input n10904;
    output \data_out[2][2] ;
    input n11245;
    input n11244;
    input n10902;
    output \data_out[2][5] ;
    input n11243;
    input n11242;
    input n11241;
    input n11240;
    output n10_adj_7;
    input n11239;
    input n11238;
    input n11237;
    input n11236;
    input n11235;
    input n11234;
    input n11233;
    input n11232;
    input n11231;
    input n11230;
    input n11229;
    input n11228;
    output \data_out[3][2] ;
    input VCC_net;
    output [7:0]rx_data;
    input n11227;
    input n11226;
    input n11225;
    input n11224;
    input n11223;
    input n11222;
    input n11221;
    input n11220;
    input n10901;
    input n11219;
    input n10900;
    input n11218;
    input n10899;
    input n11217;
    output n10705;
    input n10898;
    output \data_out[3][4] ;
    input n11216;
    input n11215;
    input n11214;
    input n11213;
    input n11212;
    output n31;
    input n11211;
    input n11210;
    input n11209;
    input n11208;
    input n11207;
    input n11206;
    input n11205;
    input n11204;
    output \data_out[3][5] ;
    input n11203;
    input n11202;
    input n11201;
    input n11200;
    input n11199;
    input n11198;
    input n11197;
    input n11196;
    input n11195;
    input n11194;
    input n11193;
    input n11192;
    input n11191;
    input n11190;
    input n11189;
    output tx2_active;
    input n11188;
    input n11187;
    input n11186;
    input n10897;
    input n10895;
    input n11185;
    output n488;
    output [7:0]\data_in_frame[6] ;
    input n11184;
    input n11183;
    input n11182;
    input n11181;
    input n11180;
    input n11179;
    input n11178;
    output data_out_10__7__N_110;
    output \data_out[10][0] ;
    output [0:0]n2698;
    input n11177;
    input n11176;
    input n11175;
    input n11174;
    input n11173;
    input n11172;
    input n11171;
    input n11170;
    input n11169;
    input n11168;
    input n11167;
    input n11166;
    input n11165;
    input n11164;
    input n11163;
    input n11162;
    input n11161;
    input n11160;
    input n11159;
    input n11158;
    input n11157;
    input n11156;
    input n11155;
    input n11154;
    input n11153;
    input n11152;
    input n11151;
    input n11150;
    input n11149;
    input n18286;
    input n18287;
    output n17392;
    output n4;
    input n11132;
    input n11131;
    output [7:0]\data_in[3] ;
    input n11130;
    input n11129;
    input n11128;
    input n11127;
    input n11126;
    input n11125;
    input n11124;
    input n11123;
    input n11121;
    input n11120;
    output n17075;
    output n9378;
    input n11119;
    input n11118;
    output n5_adj_8;
    output n17086;
    output n9;
    output n63;
    output n63_adj_9;
    output n63_adj_10;
    input n11117;
    input n11116;
    input n11115;
    output [7:0]\data_in[2] ;
    output n10_adj_11;
    input n11114;
    input n11113;
    input n11111;
    input n11110;
    input n11109;
    output n10088;
    input n11108;
    input n11107;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[1] ;
    input n11106;
    output n44;
    input n11105;
    output n10140;
    input n11104;
    input n11103;
    input n11102;
    input n11101;
    input n11100;
    input n11099;
    input n11098;
    input n11097;
    input n11096;
    input n11095;
    input n11094;
    input n11093;
    input n11092;
    input n11091;
    output n1_adj_12;
    output n10725;
    input n16618;
    input n13;
    input \rand_setpoint[0] ;
    output n9524;
    output n450;
    input \FRAME_MATCHER.state_31__N_1406[2] ;
    output n4_adj_13;
    output n4_adj_14;
    input n11033;
    input n11032;
    input n11028;
    input \rand_setpoint[25] ;
    input \rand_setpoint[17] ;
    input n11027;
    input n11025;
    input \rand_setpoint[18] ;
    input n11024;
    input n11023;
    input \rand_setpoint[19] ;
    input n11016;
    input \rand_setpoint[20] ;
    input \rand_setpoint[21] ;
    input \rand_setpoint[22] ;
    input \rand_setpoint[23] ;
    input \rand_setpoint[8] ;
    output n17327;
    output rx_data_ready;
    input \rand_setpoint[9] ;
    input \rand_setpoint[10] ;
    input \rand_setpoint[11] ;
    output n10969;
    output n10966;
    output n10963;
    output n10960;
    output n10957;
    output n10954;
    output n10951;
    output n10994;
    output \r_Bit_Index[2] ;
    input n16932;
    output [7:0]r_Tx_Data;
    input n16930;
    input n16928;
    input n16926;
    output \r_Bit_Index[1] ;
    input n10953;
    input n10956;
    input n10959;
    input n10962;
    input n10965;
    input n10968;
    input n10971;
    input n10974;
    input n16924;
    input n10996;
    input n16914;
    input n16902;
    input n18199;
    input n18073;
    output tx_o;
    output n9257;
    input n16912;
    output n5142;
    output n10972;
    output tx_enable;
    output \r_SM_Main_2__N_2031[1] ;
    output [2:0]r_SM_Main;
    output n4_adj_15;
    output [2:0]r_Bit_Index;
    input n18280;
    output n10674;
    input n10920;
    input n10923;
    input n10977;
    output n5266;
    output n17412;
    output n10976;
    output n3;
    output n8191;
    input n11039;
    input n11038;
    input n11037;
    output tx2_o;
    output tx2_enable;
    output [2:0]r_Bit_Index_adj_27;
    output n5244;
    output \r_SM_Main[1]_adj_21 ;
    output \r_SM_Main[2]_adj_22 ;
    output n17361;
    input n10983;
    input n11019;
    input n11031;
    output r_Rx_Data;
    input rx_i;
    input n11139;
    input n13744;
    input n11136;
    input n11135;
    output n1_adj_23;
    output n13116;
    input n11112;
    output n4_adj_24;
    input n11090;
    input n11089;
    input n11034;
    input n11026;
    input n10987;
    output n13692;
    output n11018;
    output n4_adj_25;
    output n9999;
    output n17708;
    output n17707;
    output n4_adj_26;
    output n10010;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n59, n65, n13662, n68, n17703, n5_c, n18172, n13146, 
        n4_c, n17404, n18281, n9334, n17697, n17696, n16096;
    wire [31:0]\FRAME_MATCHER.i ;   // coms.v(412[11:12])
    
    wire n18008, n16097;
    wire [7:0]\data_out_frame2[0] ;   // coms.v(380[12:27])
    wire [7:0]byte_transmit_counter2;   // coms.v(399[12:34])
    
    wire n17610;
    wire [31:0]\FRAME_MATCHER.i_31__N_1278 ;
    
    wire n16095;
    wire [31:0]\FRAME_MATCHER.i_31__N_1310 ;
    
    wire n276, n4_adj_2135, n18106, n18109;
    wire [31:0]\FRAME_MATCHER.state ;   // coms.v(409[11:16])
    
    wire n50;
    wire [7:0]\data_out_frame2[19] ;   // coms.v(380[12:27])
    
    wire n18274, n18277, n17764, n5_adj_2136, n18268, n10595;
    wire [7:0]\data_out[7] ;   // coms.v(21[11:19])
    
    wire n11146, n17676, n17675, n5_adj_2137, n18103, n18262, n6_c, 
        n17678, n18265, n6_adj_2138, n18067, n18061, n18256, n37, 
        n1034, n2_c, n18100, n6_adj_2139, n17761, n18259, n16740, 
        n48, n18202, n17686, n5815, n18253, n18049, n18043, n18244, 
        n6_adj_2140, n17586, n18247, n16094, n17671, n5_adj_2141, 
        n18166, n18025, n18019, n18238, n6_adj_2142, n17587, n18241, 
        n16093;
    wire [7:0]\data_out[9] ;   // coms.v(21[11:19])
    
    wire n8_c;
    wire [7:0]\data_out[10] ;   // coms.v(21[11:19])
    
    wire n17607, n18151, n18157, n18226;
    wire [7:0]\data_out[6] ;   // coms.v(21[11:19])
    
    wire n16882;
    wire [0:0]n2304;
    
    wire data_out_6__1__N_537, n12630, n6_adj_2143, n17603, n18229;
    wire [7:0]\data_out[8]_c ;   // coms.v(21[11:19])
    
    wire n2_adj_2145, n17701, n2_adj_2146, n4_adj_2147, n49, n47, 
        n16720, n4_adj_2150, n2_adj_2151, n4_adj_2152, n17747, n1_c, 
        n18220, n2_adj_2153, n4_adj_2154, n16824, n4_adj_2155, n2_adj_2156, 
        n18145, n18139, n18214, n8_adj_2157, n16092, n11002;
    wire [0:0]n2339;
    
    wire n18217;
    wire [13:0]n61;
    
    wire n10594;
    wire [13:0]delay_counter;   // coms.v(272[12:25])
    
    wire n11833, n17589, n11867, tx_active, tx_active_prev, n18208, 
        n30;
    wire [2:0]r_SM_Main_2__N_2034;
    
    wire n4650, n17568;
    wire [0:0]n1893;
    
    wire n17688, n18205, n16067;
    wire [13:0]n76;
    
    wire n16068;
    wire [0:0]n1928;
    wire [0:0]n1963;
    wire [0:0]n1998;
    wire [0:0]n2033;
    wire [0:0]n2068;
    wire [0:0]n2103;
    wire [0:0]n11;
    wire [0:0]n2173;
    wire [0:0]n2208;
    wire [0:0]n2243;
    wire [0:0]n2523;
    
    wire n18160, n17710;
    wire [0:0]n3118;
    wire [7:0]\data_out[1] ;   // coms.v(21[11:19])
    
    wire n17690, n18193, data_out_7__3__N_441, n17698, n5_adj_2159, 
        n18184;
    wire [0:0]n2374;
    
    wire n17612, n1_adj_2160;
    wire [0:0]n2409;
    
    wire n18127, n18121, n18178, n6_adj_2161, n17620, n18181, n17711;
    wire [0:0]n2444;
    
    wire n46;
    wire [0:0]n2479;
    
    wire n10815;
    wire [0:0]n2549;
    
    wire n15171, n16261;
    wire [0:0]n4334;
    
    wire n16066, n16091, n16116, n16115, n16114, n16090, n16089, 
        n445, n18163, n16088, n11079, n18094, n18097, n11084, 
        n15179, n16087, n16113, n16086, n16085, n16112, n45, n10910;
    wire [7:0]\data_out[0] ;   // coms.v(21[11:19])
    
    wire n3_c, n16084, n41, n10392, n17222, data_out_9__0__N_389, 
        n17581, n5_adj_2163, n18088, n10909, n17606, n16111, n16083, 
        n43, n2_adj_2164, n17622, n18154, n17367, n10139, n18076, 
        n17569, n26_adj_2165, n10170, n10_adj_2166, data_out_9__1__N_378, 
        n10018, n10166;
    wire [2:0]r_SM_Main_2__N_2034_adj_2405;
    wire [7:0]\data_out[5] ;   // coms.v(21[11:19])
    
    wire n56, n16, data_out_7__2__N_447, n51, n18148, n17174, n17138, 
        n17225, n22, n17200, n17201, n10316, data_out_9__4__N_344, 
        n24, n6_adj_2169, n17162, n17150, data_out_9__5__N_334, n17234, 
        n20, n17285, n17302, n10572, n10356, n16_adj_2170, n10204, 
        n10_adj_2172, n17141, n17219, n17, n17276, n17303, n17304, 
        n51_adj_2173;
    wire [7:0]\data_in_frame[0] ;   // coms.v(379[12:25])
    
    wire n2124, n18142, n10468, n10482, n10349, n17184, n15, n26_adj_2174, 
        n5817, n12491, n17490, n17255, n14, n17307, n17306, n17258, 
        n17095, n17291, n12, n4494, n17492, n17308, n10229, n6_adj_2175, 
        n17297, n14_adj_2176, n17110, n10196, n17147, n15_adj_2177, 
        n17123, n17231, n12_adj_2178, n10009, n3_adj_2179, n2120, 
        n17177, n17270, data_out_9__7__N_272, n16110, n10447, n17129, 
        n17252, n12_adj_2180, n16082, n17261, data_out_10__0__N_219, 
        n17294, n10428, n17295, n3_adj_2181, n6_adj_2182, n17156, 
        n10908, n8_adj_2183, n17243, n10440, n10346, n17165, n15_adj_2185, 
        n2_adj_2186, n4_adj_2187, n17240, n14_adj_2188, n17288, n17296, 
        n10395, n10_adj_2189, n10456, n17237, n17209, n10259, n16081, 
        n2122, n10223, n10334, n10_adj_2190, n17264, n10_adj_2191, 
        n65_adj_2192, n3_adj_2193;
    wire [7:0]\data_in_frame[2] ;   // coms.v(379[12:25])
    
    wire n10215, n20_adj_2195, n17180, n10_adj_2196, n17197, data_out_10__1__N_168, 
        n17712, n10179, data_out_10__2__N_157, n10903;
    wire [7:0]\data_out[2] ;   // coms.v(21[11:19])
    
    wire n6_adj_2197, data_out_10__3__N_146, n8_adj_2198, n2138;
    wire [7:0]\data_in_frame[1] ;   // coms.v(379[12:25])
    
    wire n23, n16080, n17309, n17315, n28_adj_2200, n18136, n22_adj_2201, 
        n27_adj_2202, n10513, n17153, n17168, n26_adj_2203, n17194, 
        n17216, n27_adj_2204, n16079, n10520, n25, n10183, data_out_10__4__N_135, 
        n16109, n10263, n15_adj_2205, n14_adj_2206, n17275, n2137, 
        n18, n16108, n17072;
    wire [7:0]\data_in_frame[3] ;   // coms.v(379[12:25])
    
    wire n11046, n10424, n10_adj_2207, data_out_10__5__N_124, n2128, 
        n26_adj_2210, n16078, n16077, n30_adj_2213, n16107, n17_adj_2214, 
        n6_adj_2215, n6_adj_2216, n17107, n17246, n5_adj_2217, n17300, 
        n30_adj_2218, n16076, n10188, data_out_10__6__N_113, n34, 
        n17116, n17171, n17132, n32, n17187, n17228, n17267, n33, 
        n16075, n10563, n31_c, n17301, n11047, n6_adj_2221, n17279, 
        n16106, n10548, n10530, n16074, n10504, n10492, n20_adj_2223, 
        data_out_10__7__N_101, n19_adj_2224, n17135, n21, n11048, 
        n17310, n2_adj_2225, n3_adj_2226, n3_adj_2227, n2126, n17206, 
        n6_adj_2228, n2_adj_2229, n3_adj_2230, n2_adj_2231, n3_adj_2232, 
        n2_adj_2233, n3_adj_2234, n2_adj_2235, n3_adj_2236, n2_adj_2237, 
        n3_adj_2238, n2_adj_2239, n3_adj_2240, n2_adj_2241, n3_adj_2242, 
        n2_adj_2243, n3_adj_2244, n2_adj_2245, n3_adj_2246, n2_adj_2247, 
        n3_adj_2248, n2_adj_2249, n3_adj_2250, n2_adj_2251, n3_adj_2252, 
        n2_adj_2253, n3_adj_2254, n16105, n16073, n17714, n15978, 
        tx2_transmit_N_1996, n2_adj_2256, n3_adj_2257, n2_adj_2258, 
        n3_adj_2259, n2_adj_2260, n3_adj_2261, n16104, n16072, n2_adj_2263, 
        n3_adj_2264, n2_adj_2265, n3_adj_2266, n2_adj_2267, n3_adj_2268, 
        n2_adj_2269, n3_adj_2270, n2_adj_2271, n3_adj_2272, n2_adj_2273, 
        n3_adj_2274, n2_adj_2275, n3_adj_2276, n2_adj_2277, n3_adj_2278, 
        n2_adj_2279, n3_adj_2280, n2_adj_2281, n3_adj_2282, n2_adj_2283, 
        n2_adj_2284, n2_adj_2285, n3_adj_2286, n2_adj_2287, n3_adj_2288, 
        n17312, n18064, n5_adj_2289, n10554, n18058, n18052, n18055, 
        n18046, n18040, n9157, n18034, n17440, n17439, n18037, 
        n18028, n18031, n18022, n5_adj_2290, n18016, n17713, n15977, 
        n15976, n15975, n15974, n18010, n15973, n18013, n15972, 
        n17659, n11049, n15_adj_2291, n17249, n14_adj_2292, n17290, 
        n18130, n18133, n16103, n13284, n16102, n10507, n16_adj_2293, 
        n17092, n17_adj_2294, n17282, n17313, n13628, n11050, n11051, 
        n9369, n16784, n7, n7_adj_2295, n10533, n14_adj_2296, n11052, 
        n17213, n10_adj_2297, n12_adj_2298, n17101, n39, n17076;
    wire [7:0]\data_in_frame[5] ;   // coms.v(379[12:25])
    
    wire n11043, n10_adj_2299, n10437, n17250, n7_adj_2300, n10472, 
        n18124, n10462, n10407, n16782, n16766, n10896;
    wire [7:0]\data_out[3] ;   // coms.v(21[11:19])
    
    wire n16780, n7_adj_2301, n13426, n7_adj_2302, n19_adj_2303, n17114, 
        n7_adj_2304, n7_adj_2305, n16768, n16101, n16764, n7_adj_2306, 
        n7_adj_2307, n10371, n14_adj_2308, n11053, n7_adj_2309, n16760, 
        n15_adj_2310, n16758, n7_adj_2311, n16756, n17098, n15_adj_2312, 
        n16754, n16752, n17203, n17284, n16750, n16071, n16070, 
        n16100, n16475, n5_adj_2315, n18_adj_2316, n11044, n10326, 
        n17126, n17373, n24_adj_2317, n17273, n6_adj_2318, n10359, 
        n16099, n10413, data_out_9__6__N_324, data_out_9__3__N_356, 
        n10459, n22_adj_2319, n16_adj_2320, n16700, n17_adj_2321, 
        n17274, n16744, n16698, n23_adj_2322, n21_adj_2323, n19_adj_2324, 
        n17215, n4_adj_2325, n2_adj_2326, n16746, n16658, n16748, 
        n16696, n16718, n16702, n16690, n16688, n13381, n16714, 
        n16686, n8_adj_2327, n8_adj_2328, n8_adj_2329, n16704, n16670, 
        n8_adj_2330, n8_adj_2331, n8_adj_2332, n16708, n8_adj_2333, 
        n16710, n16674, n16666, n16141, n8_adj_2334, n8_adj_2335, 
        n16716, n18285, n6_adj_2336, n16267, n9453, n5_adj_2337, 
        n10434, n6_adj_2339, n24_adj_2340, n11122, n15_adj_2341, n16069, 
        n5_adj_2343, n2_adj_2344, n4_adj_2345, n14_adj_2346, n17238, 
        n47_adj_2347, n17469, n18118, n17471, n17472, n17474, n17475, 
        n17477, n17489, n8_adj_2352, n5_adj_2353, n17102, n17214, 
        n16353, n9995, n17331, n10161, n12_adj_2355, n17410, n10133, 
        n10141, n6_adj_2356, n17406, n10027, n21_adj_2357, n17400, 
        n16474, n6_adj_2358, n8_adj_2359, n13450, n10136, n17388, 
        n18_adj_2360, n17487, n16_adj_2361, n17_adj_2362, n17402;
    wire [7:0]\data_out_frame2[20] ;   // coms.v(380[12:27])
    
    wire n22_adj_2363;
    wire [7:0]tx2_data;   // coms.v(402[13:21])
    
    wire n18115, n22_adj_2364, n22_adj_2365, n16_adj_2366, n16352, 
        n22_adj_2367, n26_adj_2368, n15164, n17_adj_2370, n22_adj_2371, 
        n22_adj_2372, n26_adj_2373, n42, n40, n28_adj_2374, n22_adj_2375, 
        n41_adj_2376, n39_adj_2377, n44_adj_2378, n48_adj_2379, n43_adj_2380, 
        n27_adj_2381, n29, n17281, n11076, n11075, n11074, n11073, 
        n11072, n11071, n11070, n11069, n11068, n11067, n11066, 
        n11065, n11064, n11063, n11062, n11061, n11060, n11059, 
        n11058, n11057, n11056, n11055, n11054, n13726, n453, 
        n11045, n11042, n16098, n11041, n11015, n11040, n11036, 
        n17069, n11035, n7_adj_2384, n17626, n15821, n17627, n17631, 
        n8_adj_2385, n17639, n17643, n17647, n17651, n18112, n17653, 
        n17574, n17583, n22_adj_2387, n18_adj_2388, n24_adj_2389, 
        n22_adj_2390, n26_adj_2391, n17585;
    
    SB_LUT4 i90_4_lut (.I0(tx_transmit_N_1947[3]), .I1(tx_transmit_N_1947[2]), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(\UART_TRANSMITTER.state[2] ), 
            .O(n59));   // coms.v(283[4] 369[11])
    defparam i90_4_lut.LUT_INIT = 16'h5350;
    SB_LUT4 i1_4_lut (.I0(tx_transmit_N_1947[3]), .I1(n59), .I2(n65), 
            .I3(n13662), .O(n68));   // coms.v(283[4] 369[11])
    defparam i1_4_lut.LUT_INIT = 16'h50dc;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15376 (.I0(byte_transmit_counter[1]), 
            .I1(n17703), .I2(n5_c), .I3(byte_transmit_counter[2]), .O(n18172));
    defparam byte_transmit_counter_1__bdd_4_lut_15376.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.i_31__N_1273 ), .I1(n3779), .I2(n13146), 
            .I3(GND_net), .O(n4_c));   // coms.v(416[12] 543[6])
    defparam i1_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i14627_4_lut (.I0(tx_transmit_N_1947[6]), .I1(tx_transmit_N_1947[5]), 
            .I2(n444), .I3(tx_transmit_N_1947[4]), .O(n17404));
    defparam i14627_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut (.I0(\UART_TRANSMITTER.state[0] ), .I1(n17404), .I2(tx_transmit_N_1947[7]), 
            .I3(n68), .O(n18281));   // coms.v(283[4] 369[11])
    defparam i3_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut (.I0(n2061), .I1(n13146), .I2(GND_net), .I3(GND_net), 
            .O(n9334));   // coms.v(443[6] 445[9])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 n18172_bdd_4_lut (.I0(n18172), .I1(n17697), .I2(n17696), .I3(byte_transmit_counter[2]), 
            .O(n18175));
    defparam n18172_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_977_20 (.CI(n16096), .I0(\FRAME_MATCHER.i [18]), .I1(n18008), 
            .CO(n16097));
    SB_LUT4 i15153_3_lut (.I0(\data_out_frame2[0] [7]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17610));
    defparam i15153_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 add_977_19_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [17]), .I1(\FRAME_MATCHER.i [17]), 
            .I2(n18008), .I3(n16095), .O(\FRAME_MATCHER.i_31__N_1278 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_19_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_4_lut_adj_404 (.I0(n276), .I1(n4408), .I2(\FRAME_MATCHER.i_31__N_1275 ), 
            .I3(n13146), .O(n4_adj_2135));
    defparam i1_4_lut_adj_404.LUT_INIT = 16'hbaaa;
    SB_LUT4 n18106_bdd_4_lut (.I0(n18106), .I1(\data_out_frame2[9] [5]), 
            .I2(\data_out_frame2[8] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n18109));
    defparam n18106_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i21_4_lut (.I0(\FRAME_MATCHER.state [13]), .I1(\FRAME_MATCHER.state [4]), 
            .I2(\FRAME_MATCHER.state [19]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n50));   // coms.v(494[5:21])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [4]), .I2(\data_out_frame2[19] [4]), 
            .I3(byte_transmit_counter2[1]), .O(n18274));
    defparam byte_transmit_counter2_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n18274_bdd_4_lut (.I0(n18274), .I1(\data_out_frame2[17] [4]), 
            .I2(\data_out_frame2[16] [4]), .I3(byte_transmit_counter2[1]), 
            .O(n18277));
    defparam n18274_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n17764), .I2(n5_adj_2136), .I3(byte_transmit_counter[2]), 
            .O(n18268));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_4_lut (.I0(n10595), .I1(n2593[0]), .I2(\rand_setpoint[15] ), 
            .I3(\data_out[7] [7]), .O(n11146));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 n18268_bdd_4_lut (.I0(n18268), .I1(n17676), .I2(n17675), .I3(byte_transmit_counter[2]), 
            .O(n18271));
    defparam n18268_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame2[6] [7]), 
            .I1(\data_out_frame2[7] [7]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2137));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut (.I0(byte_transmit_counter2[2]), 
            .I1(n18109), .I2(n18103), .I3(byte_transmit_counter2[3]), 
            .O(n18262));
    defparam byte_transmit_counter2_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n18262_bdd_4_lut (.I0(n18262), .I1(n6_c), .I2(n17678), .I3(byte_transmit_counter2[3]), 
            .O(n18265));
    defparam n18262_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut (.I0(\data_out_frame2[5] [7]), 
            .I1(n5_adj_2137), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2138));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15440 (.I0(byte_transmit_counter2[2]), 
            .I1(n18067), .I2(n18061), .I3(byte_transmit_counter2[3]), 
            .O(n18256));
    defparam byte_transmit_counter2_2__bdd_4_lut_15440.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_405 (.I0(n13146), .I1(\FRAME_MATCHER.i [0]), .I2(GND_net), 
            .I3(GND_net), .O(n37));
    defparam i1_2_lut_adj_405.LUT_INIT = 16'h8888;
    SB_LUT4 i10674_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [14]));   // coms.v(430[13] 433[7])
    defparam i10674_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_219_Select_0_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [0]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_c));
    defparam select_219_Select_0_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15311 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [5]), .I2(\data_out_frame2[15] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n18100));
    defparam byte_transmit_counter2_0__bdd_4_lut_15311.LUT_INIT = 16'he4aa;
    SB_LUT4 n18256_bdd_4_lut (.I0(n18256), .I1(n6_adj_2139), .I2(n17761), 
            .I3(byte_transmit_counter2[3]), .O(n18259));
    defparam n18256_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_406 (.I0(\FRAME_MATCHER.state [31]), .I1(n4_adj_2135), 
            .I2(GND_net), .I3(GND_net), .O(n16740));
    defparam i1_2_lut_adj_406.LUT_INIT = 16'h8888;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [16]), 
            .I2(\FRAME_MATCHER.state [21]), .I3(\FRAME_MATCHER.state [10]), 
            .O(n48));   // coms.v(494[5:21])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 n18250_bdd_4_lut (.I0(n18202), .I1(n17686), .I2(\data_out_frame2[0] [4]), 
            .I3(n5815), .O(n18253));
    defparam n18250_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_977_19 (.CI(n16095), .I0(\FRAME_MATCHER.i [17]), .I1(n18008), 
            .CO(n16096));
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15435 (.I0(byte_transmit_counter2[2]), 
            .I1(n18049), .I2(n18043), .I3(byte_transmit_counter2[3]), 
            .O(n18244));
    defparam byte_transmit_counter2_2__bdd_4_lut_15435.LUT_INIT = 16'he4aa;
    SB_LUT4 n18244_bdd_4_lut (.I0(n18244), .I1(n6_adj_2140), .I2(n17586), 
            .I3(byte_transmit_counter2[3]), .O(n18247));
    defparam n18244_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_977_18_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [16]), .I1(\FRAME_MATCHER.i [16]), 
            .I2(n18008), .I3(n16094), .O(\FRAME_MATCHER.i_31__N_1278 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_18_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15366 (.I0(byte_transmit_counter[1]), 
            .I1(n17671), .I2(n5_adj_2141), .I3(byte_transmit_counter[2]), 
            .O(n18166));
    defparam byte_transmit_counter_1__bdd_4_lut_15366.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15425 (.I0(byte_transmit_counter2[2]), 
            .I1(n18025), .I2(n18019), .I3(byte_transmit_counter2[3]), 
            .O(n18238));
    defparam byte_transmit_counter2_2__bdd_4_lut_15425.LUT_INIT = 16'he4aa;
    SB_CARRY add_977_18 (.CI(n16094), .I0(\FRAME_MATCHER.i [16]), .I1(n18008), 
            .CO(n16095));
    SB_LUT4 n18238_bdd_4_lut (.I0(n18238), .I1(n6_adj_2142), .I2(n17587), 
            .I3(byte_transmit_counter2[3]), .O(n18241));
    defparam n18238_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_407 (.I0(n13146), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [4]));
    defparam i1_2_lut_adj_407.LUT_INIT = 16'h8888;
    SB_LUT4 add_977_17_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [15]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(n18008), .I3(n16093), .O(\FRAME_MATCHER.i_31__N_1278 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_17_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i8_3_lut (.I0(\data_out[8] [7]), 
            .I1(\data_out[9] [7]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_c));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i10_4_lut (.I0(n8_c), .I1(\data_out[10] [7]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15018_2_lut (.I0(\data_out[1][7] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17607));
    defparam i15018_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15420 (.I0(byte_transmit_counter2[2]), 
            .I1(n18151), .I2(n18157), .I3(byte_transmit_counter2[3]), 
            .O(n18226));
    defparam byte_transmit_counter2_2__bdd_4_lut_15420.LUT_INIT = 16'he4aa;
    SB_LUT4 i11_4_lut (.I0(\rand_setpoint[16] ), .I1(\data_out[6] [0]), 
            .I2(n10596), .I3(n2593[0]), .O(n16882));
    defparam i11_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i10514_2_lut (.I0(\rand_setpoint[31] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2304[0]));   // coms.v(283[4] 369[11])
    defparam i10514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9952_3_lut (.I0(data_out_6__1__N_537), .I1(\data_out[7] [0]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n12630));   // coms.v(19[11:32])
    defparam i9952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n18100_bdd_4_lut (.I0(n18100), .I1(\data_out_frame2[13] [5]), 
            .I2(\data_out_frame2[12] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n18103));
    defparam n18100_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n18226_bdd_4_lut (.I0(n18226), .I1(n6_adj_2143), .I2(n17603), 
            .I3(byte_transmit_counter2[3]), .O(n18229));
    defparam n18226_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9896_3_lut (.I0(\data_out[8]_c [0]), .I1(\data_out[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n8));   // coms.v(19[11:32])
    defparam i9896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n18166_bdd_4_lut (.I0(n18166), .I1(n2_adj_2145), .I2(n17701), 
            .I3(byte_transmit_counter[2]), .O(n18169));
    defparam n18166_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSS byte_transmit_counter2_i5 (.Q(byte_transmit_counter2[5]), .C(CLK_c), 
            .D(n2_adj_2146), .S(n4_adj_2147));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i2_3_lut (.I0(\data_out[2][0] ), 
            .I1(\data_out[3][0] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20_4_lut (.I0(\FRAME_MATCHER.state [5]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(\FRAME_MATCHER.state [18]), 
            .O(n49));   // coms.v(494[5:21])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.state [28]), .I1(\FRAME_MATCHER.state [11]), 
            .I2(\FRAME_MATCHER.state [15]), .I3(\FRAME_MATCHER.state [24]), 
            .O(n47));   // coms.v(494[5:21])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9953_4_lut (.I0(\data_out[6] [0]), .I1(n12630), .I2(byte_transmit_counter[0]), 
            .I3(byte_transmit_counter[1]), .O(n6));   // coms.v(19[11:32])
    defparam i9953_4_lut.LUT_INIT = 16'hcac0;
    SB_DFFSS byte_transmit_counter2_i4 (.Q(byte_transmit_counter2[4]), .C(CLK_c), 
            .D(n16720), .S(n4_adj_2150));   // coms.v(416[12] 543[6])
    SB_DFFSS byte_transmit_counter2_i3 (.Q(byte_transmit_counter2[3]), .C(CLK_c), 
            .D(n2_adj_2151), .S(n4_adj_2152));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15445 (.I0(byte_transmit_counter[1]), 
            .I1(n17747), .I2(n1_c), .I3(byte_transmit_counter[2]), .O(n18220));
    defparam byte_transmit_counter_1__bdd_4_lut_15445.LUT_INIT = 16'he4aa;
    SB_DFFSS byte_transmit_counter2_i2 (.Q(byte_transmit_counter2[2]), .C(CLK_c), 
            .D(n2_adj_2153), .S(n4_adj_2154));   // coms.v(416[12] 543[6])
    SB_DFFSS byte_transmit_counter2_i1 (.Q(byte_transmit_counter2[1]), .C(CLK_c), 
            .D(n16824), .S(n4_adj_2155));   // coms.v(416[12] 543[6])
    SB_LUT4 n18220_bdd_4_lut (.I0(n18220), .I1(n2_adj_2156), .I2(n17607), 
            .I3(byte_transmit_counter[2]), .O(n18223));
    defparam n18220_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_977_17 (.CI(n16093), .I0(\FRAME_MATCHER.i [15]), .I1(n18008), 
            .CO(n16094));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i2_3_lut (.I0(\data_out[2][7] ), 
            .I1(\data_out[3][7] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2156));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15410 (.I0(byte_transmit_counter2[2]), 
            .I1(n18145), .I2(n18139), .I3(byte_transmit_counter2[3]), 
            .O(n18214));
    defparam byte_transmit_counter2_2__bdd_4_lut_15410.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i8_3_lut (.I0(\data_out[8][6] ), 
            .I1(\data_out[9] [6]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2157));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_977_16_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [14]), .I1(\FRAME_MATCHER.i [14]), 
            .I2(n18008), .I3(n16092), .O(\FRAME_MATCHER.i_31__N_1278 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_16_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_977_16 (.CI(n16092), .I0(\FRAME_MATCHER.i [14]), .I1(n18008), 
            .CO(n16093));
    SB_LUT4 i8316_4_lut_4_lut (.I0(n10595), .I1(n2593[0]), .I2(\rand_setpoint[12] ), 
            .I3(\data_out[7] [4]), .O(n11002));
    defparam i8316_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 i10513_2_lut (.I0(\rand_setpoint[30] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2339[0]));   // coms.v(283[4] 369[11])
    defparam i10513_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n18214_bdd_4_lut (.I0(n18214), .I1(n6_adj_2138), .I2(n17610), 
            .I3(byte_transmit_counter2[3]), .O(n18217));
    defparam n18214_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE delay_counter_2361__i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n10594), 
            .D(n61[0]));   // coms.v(305[16] 313[10])
    SB_LUT4 i1_2_lut_adj_408 (.I0(byte_transmit_counter2[1]), .I1(n11833), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2155));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_408.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i10_4_lut (.I0(n8_adj_2157), 
            .I1(\data_out[10] [6]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_3));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_409 (.I0(\FRAME_MATCHER.i_31__N_1272 ), .I1(n17589), 
            .I2(byte_transmit_counter2[1]), .I3(n11867), .O(n16824));
    defparam i1_4_lut_adj_409.LUT_INIT = 16'ha088;
    SB_DFF tx_active_prev_2167 (.Q(tx_active_prev), .C(CLK_c), .D(tx_active));   // coms.v(280[12] 370[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15450 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [4]), .I2(\data_out_frame2[11] [4]), 
            .I3(byte_transmit_counter2[1]), .O(n18208));
    defparam byte_transmit_counter2_0__bdd_4_lut_15450.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_410 (.I0(\FRAME_MATCHER.state [12]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(GND_net), .I3(GND_net), .O(n30));   // coms.v(494[5:21])
    defparam i1_2_lut_adj_410.LUT_INIT = 16'heeee;
    SB_DFFSR tx_transmit_2168 (.Q(r_SM_Main_2__N_2034[0]), .C(CLK_c), .D(n18281), 
            .R(n4650));   // coms.v(280[12] 370[6])
    SB_LUT4 n18208_bdd_4_lut (.I0(n18208), .I1(\data_out_frame2[9] [4]), 
            .I2(\data_out_frame2[8] [4]), .I3(byte_transmit_counter2[1]), 
            .O(n17568));
    defparam n18208_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \data_out_7[[3__2197  (.Q(\data_out[7] [3]), .C(CLK_c), .E(n10595), 
            .D(n1893[0]));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_adj_411 (.I0(n11833), .I1(byte_transmit_counter2[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2154));   // coms.v(409[11:16])
    defparam i1_2_lut_adj_411.LUT_INIT = 16'h8888;
    SB_LUT4 n18202_bdd_4_lut (.I0(n18202), .I1(n17688), .I2(\data_out_frame2[0] [3]), 
            .I3(n5815), .O(n18205));
    defparam n18202_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY delay_counter_2361_add_4_4 (.CI(n16067), .I0(GND_net), .I1(n76[2]), 
            .CO(n16068));
    SB_DFFE \data_out_7[[2__2198  (.Q(\data_out[7] [2]), .C(CLK_c), .E(n10595), 
            .D(n1928[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_7[[1__2199  (.Q(\data_out[7] [1]), .C(CLK_c), .E(n10595), 
            .D(n1963[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_7[[0__2200  (.Q(\data_out[7] [0]), .C(CLK_c), .E(n10595), 
            .D(n1998[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_6[[7__2201  (.Q(\data_out[6] [7]), .C(CLK_c), .E(n10596), 
            .D(n2033[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_6[[6__2202  (.Q(\data_out[6] [6]), .C(CLK_c), .E(n10596), 
            .D(n2068[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_6[[5__2203  (.Q(\data_out[6] [5]), .C(CLK_c), .E(n10596), 
            .D(n2103[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_6[[4__2204  (.Q(\data_out[6] [4]), .C(CLK_c), .E(n10596), 
            .D(n11[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_6[[3__2205  (.Q(\data_out[6] [3]), .C(CLK_c), .E(n10596), 
            .D(n2173[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_6[[2__2206  (.Q(\data_out[6] [2]), .C(CLK_c), .E(n10596), 
            .D(n2208[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_6[[1__2207  (.Q(\data_out[6] [1]), .C(CLK_c), .E(n10596), 
            .D(n2243[0]));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_5[[1__2215  (.Q(\data_out[5][1] ), .C(CLK_c), .E(n10596), 
            .D(n2523[0]));   // coms.v(280[12] 370[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15395 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [0]), .I2(\data_out_frame2[19] [0]), 
            .I3(byte_transmit_counter2[1]), .O(n18160));
    defparam byte_transmit_counter2_0__bdd_4_lut_15395.LUT_INIT = 16'he4aa;
    SB_LUT4 select_224_Select_2_i2_4_lut (.I0(byte_transmit_counter2[2]), 
            .I1(\FRAME_MATCHER.i_31__N_1272 ), .I2(n17710), .I3(n11867), 
            .O(n2_adj_2153));
    defparam select_224_Select_2_i2_4_lut.LUT_INIT = 16'h88c0;
    SB_DFFE \data_out_1[[1__2247  (.Q(\data_out[1] [1]), .C(CLK_c), .E(n10596), 
            .D(n3118[0]));   // coms.v(280[12] 370[6])
    SB_DFF \UART_TRANSMITTER.state__i1  (.Q(\UART_TRANSMITTER.state[0] ), 
           .C(CLK_c), .D(n16614));   // coms.v(280[12] 370[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(CLK_c), 
           .D(n16662));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_0[[0__2256  (.Q(\data_out[0][0] ), .C(CLK_c), .D(n10914));   // coms.v(280[12] 370[6])
    SB_LUT4 i5_3_lut (.I0(\data_out[6] [7]), .I1(\data_out[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_c));   // coms.v(19[11:32])
    defparam i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n18190_bdd_4_lut (.I0(n18202), .I1(n17690), .I2(\data_out_frame2[0] [2]), 
            .I3(n5815), .O(n18193));
    defparam n18190_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15148_2_lut (.I0(data_out_7__3__N_441), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17747));
    defparam i15148_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \data_out_0[[1__2255  (.Q(\data_out[0][1] ), .C(CLK_c), .D(n10913));   // coms.v(280[12] 370[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15405 (.I0(byte_transmit_counter[1]), 
            .I1(n17698), .I2(n5_adj_2159), .I3(byte_transmit_counter[2]), 
            .O(n18184));
    defparam byte_transmit_counter_1__bdd_4_lut_15405.LUT_INIT = 16'he4aa;
    SB_LUT4 i10508_2_lut (.I0(\rand_setpoint[29] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2374[0]));   // coms.v(283[4] 369[11])
    defparam i10508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n18184_bdd_4_lut (.I0(n18184), .I1(n17612), .I2(n1_adj_2160), 
            .I3(byte_transmit_counter[2]), .O(n18187));
    defparam n18184_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10505_2_lut (.I0(\rand_setpoint[28] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2409[0]));   // coms.v(283[4] 369[11])
    defparam i10505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_412 (.I0(n11833), .I1(byte_transmit_counter2[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2152));   // coms.v(409[11:16])
    defparam i1_2_lut_adj_412.LUT_INIT = 16'h8888;
    SB_DFF \data_out_0[[3__2253  (.Q(\data_out[0][3] ), .C(CLK_c), .D(n10912));   // coms.v(280[12] 370[6])
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15400 (.I0(byte_transmit_counter2[2]), 
            .I1(n18127), .I2(n18121), .I3(byte_transmit_counter2[3]), 
            .O(n18178));
    defparam byte_transmit_counter2_2__bdd_4_lut_15400.LUT_INIT = 16'he4aa;
    SB_LUT4 n18178_bdd_4_lut (.I0(n18178), .I1(n6_adj_2161), .I2(n17620), 
            .I3(byte_transmit_counter2[3]), .O(n18181));
    defparam n18178_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_224_Select_3_i2_4_lut (.I0(byte_transmit_counter2[3]), 
            .I1(\FRAME_MATCHER.i_31__N_1272 ), .I2(n17711), .I3(n11867), 
            .O(n2_adj_2151));
    defparam select_224_Select_3_i2_4_lut.LUT_INIT = 16'h88c0;
    SB_LUT4 i10472_2_lut (.I0(\rand_setpoint[27] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2444[0]));   // coms.v(283[4] 369[11])
    defparam i10472_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [25]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [26]), 
            .O(n46));   // coms.v(494[5:21])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10471_2_lut (.I0(\rand_setpoint[26] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2479[0]));   // coms.v(283[4] 369[11])
    defparam i10471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15194_2_lut (.I0(n10596), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n10815));
    defparam i15194_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i10561_2_lut (.I0(\rand_setpoint[24] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2549[0]));   // coms.v(283[4] 369[11])
    defparam i10561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_413 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [0]), 
            .I2(GND_net), .I3(GND_net), .O(n15171));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_413.LUT_INIT = 16'hbbbb;
    SB_LUT4 mux_1818_i1_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n16261), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(\FRAME_MATCHER.state[1] ), 
            .O(n4334[0]));   // coms.v(434[4] 542[11])
    defparam mux_1818_i1_4_lut.LUT_INIT = 16'h7570;
    SB_LUT4 delay_counter_2361_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[1]), .I3(n16066), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_977_15_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [13]), .I1(\FRAME_MATCHER.i [13]), 
            .I2(n18008), .I3(n16091), .O(\FRAME_MATCHER.i_31__N_1278 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_15_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_2506_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n16116), .O(tx_transmit_N_1947[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2506_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2506_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n16115), .O(tx_transmit_N_1947[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2506_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_977_15 (.CI(n16091), .I0(\FRAME_MATCHER.i [13]), .I1(n18008), 
            .CO(n16092));
    SB_CARRY delay_counter_2361_add_4_3 (.CI(n16066), .I0(GND_net), .I1(n76[1]), 
            .CO(n16067));
    SB_CARRY add_2506_8 (.CI(n16115), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n16116));
    SB_LUT4 add_2506_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n16114), .O(tx_transmit_N_1947[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2506_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_977_14_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [12]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(n18008), .I3(n16090), .O(\FRAME_MATCHER.i_31__N_1278 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_14_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_977_14 (.CI(n16090), .I0(\FRAME_MATCHER.i [12]), .I1(n18008), 
            .CO(n16091));
    SB_LUT4 add_977_13_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [11]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(n18008), .I3(n16089), .O(\FRAME_MATCHER.i_31__N_1278 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_13_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 delay_counter_2361_add_4_2_lut (.I0(GND_net), .I1(n445), .I2(n76[0]), 
            .I3(GND_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_977_13 (.CI(n16089), .I0(\FRAME_MATCHER.i [11]), .I1(n18008), 
            .CO(n16090));
    SB_LUT4 n18160_bdd_4_lut (.I0(n18160), .I1(\data_out_frame2[17] [0]), 
            .I2(\data_out_frame2[16] [0]), .I3(byte_transmit_counter2[1]), 
            .O(n18163));
    defparam n18160_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_977_12_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [10]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(n18008), .I3(n16088), .O(\FRAME_MATCHER.i_31__N_1278 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_12_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i8393_4_lut_4_lut (.I0(n10595), .I1(n2593[0]), .I2(\rand_setpoint[13] ), 
            .I3(\data_out[7] [5]), .O(n11079));
    defparam i8393_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15306 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [5]), .I2(\data_out_frame2[19] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n18094));
    defparam byte_transmit_counter2_0__bdd_4_lut_15306.LUT_INIT = 16'he4aa;
    SB_LUT4 n18094_bdd_4_lut (.I0(n18094), .I1(\data_out_frame2[17] [5]), 
            .I2(\data_out_frame2[16] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n18097));
    defparam n18094_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_414 (.I0(byte_transmit_counter2[4]), .I1(n11833), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2150));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_414.LUT_INIT = 16'h8888;
    SB_LUT4 i8398_4_lut_4_lut (.I0(n10595), .I1(n2593[0]), .I2(\rand_setpoint[14] ), 
            .I3(\data_out[7] [6]), .O(n11084));
    defparam i8398_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_CARRY delay_counter_2361_add_4_2 (.CI(GND_net), .I0(n445), .I1(n76[0]), 
            .CO(n16066));
    SB_LUT4 i1_2_lut_adj_415 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [0]), 
            .I2(GND_net), .I3(GND_net), .O(n15179));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_415.LUT_INIT = 16'heeee;
    SB_CARRY add_2506_7 (.CI(n16114), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n16115));
    SB_CARRY add_977_12 (.CI(n16088), .I0(\FRAME_MATCHER.i [10]), .I1(n18008), 
            .CO(n16089));
    SB_LUT4 add_977_11_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [9]), .I1(\FRAME_MATCHER.i [9]), 
            .I2(n18008), .I3(n16087), .O(\FRAME_MATCHER.i_31__N_1278 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_11_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_2506_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n16113), .O(tx_transmit_N_1947[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2506_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_977_11 (.CI(n16087), .I0(\FRAME_MATCHER.i [9]), .I1(n18008), 
            .CO(n16088));
    SB_LUT4 add_977_10_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [8]), .I1(\FRAME_MATCHER.i [8]), 
            .I2(n18008), .I3(n16086), .O(\FRAME_MATCHER.i_31__N_1278 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_10_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_2506_6 (.CI(n16113), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n16114));
    SB_CARRY add_977_10 (.CI(n16086), .I0(\FRAME_MATCHER.i [8]), .I1(n18008), 
            .CO(n16087));
    SB_LUT4 add_977_9_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [7]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(n18008), .I3(n16085), .O(\FRAME_MATCHER.i_31__N_1278 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_2506_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n16112), .O(tx_transmit_N_1947[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2506_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.state [23]), .I1(\FRAME_MATCHER.state [9]), 
            .I2(\FRAME_MATCHER.state [17]), .I3(\FRAME_MATCHER.state [29]), 
            .O(n45));   // coms.v(494[5:21])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \data_out_0[[5__2251  (.Q(\data_out[0][5] ), .C(CLK_c), .D(n10911));   // coms.v(280[12] 370[6])
    SB_DFF \data_out_0[[6__2250  (.Q(\data_out[0] [6]), .C(CLK_c), .D(n10910));   // coms.v(280[12] 370[6])
    SB_CARRY add_977_9 (.CI(n16085), .I0(\FRAME_MATCHER.i [7]), .I1(n18008), 
            .CO(n16086));
    SB_LUT4 add_977_8_lut (.I0(n41), .I1(\FRAME_MATCHER.i [6]), .I2(n18008), 
            .I3(n16084), .O(n3_c)) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_8_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_2506_5 (.CI(n16112), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n16113));
    SB_LUT4 i9889_3_lut (.I0(\data_out[6] [1]), .I1(\data_out[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5));   // coms.v(19[11:32])
    defparam i9889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_416 (.I0(\data_out[8][5] ), .I1(\data_out[6] [4]), 
            .I2(n10392), .I3(n17222), .O(data_out_9__0__N_389));   // coms.v(178[16:77])
    defparam i3_4_lut_adj_416.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15361 (.I0(byte_transmit_counter[1]), 
            .I1(n17581), .I2(n5_adj_2163), .I3(byte_transmit_counter[2]), 
            .O(n18088));
    defparam byte_transmit_counter_1__bdd_4_lut_15361.LUT_INIT = 16'he4aa;
    SB_DFF \data_out_1[[2__2246  (.Q(\data_out[1] [2]), .C(CLK_c), .D(n10909));   // coms.v(280[12] 370[6])
    SB_CARRY add_977_8 (.CI(n16084), .I0(\FRAME_MATCHER.i [6]), .I1(n18008), 
            .CO(n16085));
    SB_LUT4 i1_4_lut_adj_417 (.I0(\FRAME_MATCHER.i_31__N_1272 ), .I1(n17606), 
            .I2(byte_transmit_counter2[4]), .I3(n11867), .O(n16720));
    defparam i1_4_lut_adj_417.LUT_INIT = 16'ha088;
    SB_LUT4 add_2506_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n16111), .O(tx_transmit_N_1947[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2506_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_977_7_lut (.I0(n43), .I1(\FRAME_MATCHER.i [5]), .I2(n18008), 
            .I3(n16083), .O(\FRAME_MATCHER.i_31__N_1278 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_7_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 n18088_bdd_4_lut (.I0(n18088), .I1(n2_adj_2164), .I2(n17622), 
            .I3(byte_transmit_counter[2]), .O(n18091));
    defparam n18088_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15356 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [0]), .I2(\data_out_frame2[15] [0]), 
            .I3(byte_transmit_counter2[1]), .O(n18154));
    defparam byte_transmit_counter2_0__bdd_4_lut_15356.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_418 (.I0(\FRAME_MATCHER.i_31__N_1272 ), .I1(n17367), 
            .I2(\FRAME_MATCHER.state[1] ), .I3(\FRAME_MATCHER.state[2] ), 
            .O(n10139));
    defparam i1_4_lut_adj_418.LUT_INIT = 16'hbbba;
    SB_DFF byte_transmit_counter__i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
           .D(n16634));   // coms.v(280[12] 370[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15301 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [4]), .I2(\data_out_frame2[15] [4]), 
            .I3(byte_transmit_counter2[1]), .O(n18076));
    defparam byte_transmit_counter2_0__bdd_4_lut_15301.LUT_INIT = 16'he4aa;
    SB_DFF byte_transmit_counter__i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
           .D(n16632));   // coms.v(280[12] 370[6])
    SB_LUT4 n18076_bdd_4_lut (.I0(n18076), .I1(\data_out_frame2[13] [4]), 
            .I2(\data_out_frame2[12] [4]), .I3(byte_transmit_counter2[1]), 
            .O(n17569));
    defparam n18076_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF byte_transmit_counter__i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
           .D(n16630));   // coms.v(280[12] 370[6])
    SB_LUT4 i4_4_lut (.I0(n26_adj_2165), .I1(\data_out[6] [7]), .I2(n10170), 
            .I3(\data_out[6] [5]), .O(n10_adj_2166));   // coms.v(179[16:84])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_419 (.I0(\data_out[8][3] ), .I1(n10_adj_2166), 
            .I2(\data_out[8][4] ), .I3(GND_net), .O(data_out_9__1__N_378));   // coms.v(179[16:84])
    defparam i5_3_lut_adj_419.LUT_INIT = 16'h9696;
    SB_LUT4 n18154_bdd_4_lut (.I0(n18154), .I1(\data_out_frame2[13] [0]), 
            .I2(\data_out_frame2[12] [0]), .I3(byte_transmit_counter2[1]), 
            .O(n18157));
    defparam n18154_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_420 (.I0(n10018), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n10166));   // coms.v(494[5:21])
    defparam i1_2_lut_adj_420.LUT_INIT = 16'hbbbb;
    SB_DFFSR tx2_transmit_2261 (.Q(r_SM_Main_2__N_2034_adj_2405[0]), .C(CLK_c), 
            .D(n4334[0]), .R(n10018));   // coms.v(416[12] 543[6])
    SB_DFFESS \data_out_5[[0__2216  (.Q(data_out_6__1__N_537), .C(CLK_c), 
            .E(n10596), .D(n2549[0]), .S(n10815));   // coms.v(280[12] 370[6])
    SB_DFFESS \data_out_5[[2__2214  (.Q(\data_out[5] [2]), .C(CLK_c), .E(n10596), 
            .D(n2479[0]), .S(n10815));   // coms.v(280[12] 370[6])
    SB_DFFESS \data_out_5[[3__2213  (.Q(\data_out[5] [3]), .C(CLK_c), .E(n10596), 
            .D(n2444[0]), .S(n10815));   // coms.v(280[12] 370[6])
    SB_DFFESS \data_out_5[[4__2212  (.Q(\data_out[5] [4]), .C(CLK_c), .E(n10596), 
            .D(n2409[0]), .S(n10815));   // coms.v(280[12] 370[6])
    SB_DFF byte_transmit_counter__i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
           .D(n16628));   // coms.v(280[12] 370[6])
    SB_DFFESS \data_out_5[[5__2211  (.Q(\data_out[5] [5]), .C(CLK_c), .E(n10596), 
            .D(n2374[0]), .S(n10815));   // coms.v(280[12] 370[6])
    SB_LUT4 i27_4_lut (.I0(n47), .I1(n49), .I2(n48), .I3(n50), .O(n56));   // coms.v(494[5:21])
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut (.I0(\data_out_frame2[8] [2]), .I1(\data_out_frame2[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // coms.v(234[16:291])
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS \data_out_5[[6__2210  (.Q(data_out_7__2__N_447), .C(CLK_c), 
            .E(n10596), .D(n2339[0]), .S(n10815));   // coms.v(280[12] 370[6])
    SB_LUT4 i22_4_lut (.I0(\FRAME_MATCHER.state [6]), .I1(\FRAME_MATCHER.state [14]), 
            .I2(\FRAME_MATCHER.state [20]), .I3(n30), .O(n51));   // coms.v(494[5:21])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESS \data_out_5[[7__2209  (.Q(data_out_7__3__N_441), .C(CLK_c), 
            .E(n10596), .D(n2304[0]), .S(n10815));   // coms.v(280[12] 370[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15351 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [0]), .I2(\data_out_frame2[11] [0]), 
            .I3(byte_transmit_counter2[1]), .O(n18148));
    defparam byte_transmit_counter2_0__bdd_4_lut_15351.LUT_INIT = 16'he4aa;
    SB_LUT4 i9_4_lut (.I0(\data_out_frame2[9] [7]), .I1(n17174), .I2(n17138), 
            .I3(n17225), .O(n22));   // coms.v(234[16:291])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_421 (.I0(\data_out[8][6] ), .I1(\data_out[8] [7]), 
            .I2(\data_out[5] [3]), .I3(n17200), .O(n17201));   // coms.v(182[17:86])
    defparam i3_4_lut_adj_421.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i8_3_lut (.I0(\data_out[8][1] ), 
            .I1(\data_out[9] [1]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_4));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_1_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(\data_out[5] [2]), .I1(\data_out[7] [0]), .I2(n17201), 
            .I3(n10316), .O(data_out_9__4__N_344));   // coms.v(21[11:19])
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_422 (.I0(\data_out_frame2[15] [5]), .I1(n22), 
            .I2(n16), .I3(\data_out_frame2[9] [3]), .O(n24));   // coms.v(234[16:291])
    defparam i11_4_lut_adj_422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_423 (.I0(\data_out[10] [5]), .I1(\data_out[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2169));   // coms.v(182[17:86])
    defparam i1_2_lut_adj_423.LUT_INIT = 16'h6666;
    SB_CARRY add_2506_4 (.CI(n16111), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n16112));
    SB_CARRY add_977_7 (.CI(n16083), .I0(\FRAME_MATCHER.i [5]), .I1(n18008), 
            .CO(n16084));
    SB_LUT4 i4_4_lut_adj_424 (.I0(\data_out[9] [1]), .I1(n17162), .I2(n17150), 
            .I3(n6_adj_2169), .O(data_out_9__5__N_334));   // coms.v(182[17:86])
    defparam i4_4_lut_adj_424.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_425 (.I0(\data_out[9] [1]), .I1(\data_out[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17200));   // coms.v(182[17:86])
    defparam i1_2_lut_adj_425.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut (.I0(n17234), .I1(n24), .I2(n20), .I3(n17285), 
            .O(n17302));   // coms.v(234[16:291])
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame2[7] [5]), .I1(n10572), .I2(n10356), 
            .I3(\data_out_frame2[10] [0]), .O(n16_adj_2170));   // coms.v(233[16:291])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i1_3_lut (.I0(\data_out[0][1] ), 
            .I1(\data_out[1] [1]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n1));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_1_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n18148_bdd_4_lut (.I0(n18148), .I1(\data_out_frame2[9] [0]), 
            .I2(\data_out_frame2[8] [0]), .I3(byte_transmit_counter2[1]), 
            .O(n18151));
    defparam n18148_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_426 (.I0(n10204), .I1(\data_out[9] [3]), .I2(\data_out[10] [6]), 
            .I3(\data_out[7] [4]), .O(n10_adj_2172));   // coms.v(184[17:86])
    defparam i4_4_lut_adj_426.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(\data_out_frame2[16] [2]), .I1(n17141), .I2(\data_out_frame2[9] [2]), 
            .I3(n17219), .O(n17));   // coms.v(233[16:291])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_DFF \data_out_6[[0__2208  (.Q(\data_out[6] [0]), .C(CLK_c), .D(n16882));   // coms.v(280[12] 370[6])
    SB_LUT4 i9_4_lut_adj_427 (.I0(n17), .I1(n17276), .I2(n16_adj_2170), 
            .I3(n17303), .O(n17304));   // coms.v(233[16:291])
    defparam i9_4_lut_adj_427.LUT_INIT = 16'h6996;
    SB_DFF \data_out_7[[4__2196  (.Q(\data_out[7] [4]), .C(CLK_c), .D(n11002));   // coms.v(280[12] 370[6])
    SB_DFF byte_transmit_counter__i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
           .D(n16626));   // coms.v(280[12] 370[6])
    SB_LUT4 i28_4_lut (.I0(n51), .I1(n56), .I2(n45), .I3(n46), .O(n10018));   // coms.v(494[5:21])
    defparam i28_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_428 (.I0(\FRAME_MATCHER.state[1] ), .I1(n10018), 
            .I2(GND_net), .I3(GND_net), .O(n51_adj_2173));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_428.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_429 (.I0(\data_out_frame2[11] [0]), .I1(\data_out_frame2[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17276));   // coms.v(233[16:291])
    defparam i1_2_lut_adj_429.LUT_INIT = 16'h6666;
    SB_LUT4 i1012_2_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n2124));   // coms.v(67[15:26])
    defparam i1012_2_lut.LUT_INIT = 16'h6666;
    SB_DFF byte_transmit_counter__i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
           .D(n16624));   // coms.v(280[12] 370[6])
    SB_DFF byte_transmit_counter__i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
           .D(n16622));   // coms.v(280[12] 370[6])
    SB_DFF byte_transmit_counter__i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
           .D(n16620));   // coms.v(280[12] 370[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15346 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [7]), .I2(\data_out_frame2[11] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18142));
    defparam byte_transmit_counter2_0__bdd_4_lut_15346.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_430 (.I0(n10468), .I1(n10482), .I2(n10349), .I3(n17184), 
            .O(n15));   // coms.v(232[16:229])
    defparam i6_4_lut_adj_430.LUT_INIT = 16'h6996;
    SB_LUT4 i14713_4_lut (.I0(\data_out_frame2[0] [0]), .I1(n26_adj_2174), 
            .I2(n5817), .I3(n12491), .O(n17490));
    defparam i14713_4_lut.LUT_INIT = 16'hfa8a;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n17255), .I2(n14), .I3(n17276), 
            .O(n17307));   // coms.v(232[16:229])
    defparam i8_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_431 (.I0(\data_out_frame2[0] [3]), .I1(\data_out_frame2[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17306));   // coms.v(232[16:229])
    defparam i1_2_lut_adj_431.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame2[12] [4]), .I1(n17258), .I2(n17095), 
            .I3(n17291), .O(n12));   // coms.v(230[16:237])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14715_4_lut (.I0(n17490), .I1(n4494), .I2(n5815), .I3(n5817), 
            .O(n17492));
    defparam i14715_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i6_4_lut_adj_432 (.I0(n17306), .I1(n12), .I2(\data_out_frame2[16] [0]), 
            .I3(\data_out_frame2[11] [5]), .O(n17308));   // coms.v(230[16:237])
    defparam i6_4_lut_adj_432.LUT_INIT = 16'h6996;
    SB_LUT4 n18142_bdd_4_lut (.I0(n18142), .I1(\data_out_frame2[9] [7]), 
            .I2(\data_out_frame2[8] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n18145));
    defparam n18142_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_433 (.I0(\data_out_frame2[0] [2]), .I1(n10229), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2175));   // coms.v(230[16:237])
    defparam i1_2_lut_adj_433.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_434 (.I0(\data_out_frame2[14] [2]), .I1(\data_out_frame2[7] [2]), 
            .I2(\data_out_frame2[11] [4]), .I3(n6_adj_2175), .O(n17258));   // coms.v(230[16:237])
    defparam i4_4_lut_adj_434.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_435 (.I0(\data_out[7] [2]), .I1(\data_out[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10316));   // coms.v(182[17:86])
    defparam i1_2_lut_adj_435.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_436 (.I0(n17297), .I1(\data_out[9] [5]), .I2(data_out_7__2__N_447), 
            .I3(GND_net), .O(n14_adj_2176));   // coms.v(177[16:77])
    defparam i5_3_lut_adj_436.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_437 (.I0(n10316), .I1(n17110), .I2(n10196), .I3(n17147), 
            .O(n15_adj_2177));   // coms.v(177[16:77])
    defparam i6_4_lut_adj_437.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame2[9] [5]), .I1(\data_out_frame2[7] [6]), 
            .I2(\data_out_frame2[5] [7]), .I3(GND_net), .O(n17138));   // coms.v(234[16:291])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_438 (.I0(n17123), .I1(n17231), .I2(n17138), .I3(n17258), 
            .O(n12_adj_2178));   // coms.v(227[16:31])
    defparam i5_4_lut_adj_438.LUT_INIT = 16'h6996;
    SB_LUT4 select_219_Select_4_i3_2_lut_3_lut (.I0(n13146), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n10009), .I3(GND_net), .O(n3_adj_2179));
    defparam select_219_Select_4_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1008_2_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n2120));   // coms.v(65[15:26])
    defparam i1008_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_439 (.I0(n15_adj_2177), .I1(n17177), .I2(n14_adj_2176), 
            .I3(n17270), .O(data_out_9__7__N_272));   // coms.v(177[16:77])
    defparam i8_4_lut_adj_439.LUT_INIT = 16'h9669;
    SB_LUT4 add_2506_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n16110), .O(tx_transmit_N_1947[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2506_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut_adj_440 (.I0(n10447), .I1(n17129), .I2(\data_out[9] [3]), 
            .I3(n17252), .O(n12_adj_2180));   // coms.v(174[16:77])
    defparam i5_4_lut_adj_440.LUT_INIT = 16'h6996;
    SB_LUT4 add_977_6_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [4]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n18008), .I3(n16082), .O(\FRAME_MATCHER.i_31__N_1278 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i6_4_lut_adj_441 (.I0(n17261), .I1(n12_adj_2180), .I2(\data_out[7] [3]), 
            .I3(\data_out[7] [6]), .O(data_out_10__0__N_219));   // coms.v(174[16:77])
    defparam i6_4_lut_adj_441.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_442 (.I0(n17294), .I1(n12_adj_2178), .I2(n10428), 
            .I3(\data_out_frame2[15] [2]), .O(n17295));   // coms.v(227[16:31])
    defparam i6_4_lut_adj_442.LUT_INIT = 16'h6996;
    SB_CARRY add_977_6 (.CI(n16082), .I0(\FRAME_MATCHER.i [4]), .I1(n18008), 
            .CO(n16083));
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2_c), .S(n3_adj_2181));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i152 (.Q(\data_out_frame2[18] [7]), .C(CLK_c), 
           .D(n11260));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_adj_443 (.I0(\data_out[5] [4]), .I1(\data_out[9][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n10204));   // coms.v(184[17:86])
    defparam i1_2_lut_adj_443.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_444 (.I0(\data_out[9] [0]), .I1(\data_out[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17150));   // coms.v(181[17:93])
    defparam i1_2_lut_adj_444.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_445 (.I0(\data_out_frame2[11] [0]), .I1(\data_out_frame2[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2182));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_445.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i151 (.Q(\data_out_frame2[18] [6]), .C(CLK_c), 
           .D(n11259));   // coms.v(416[12] 543[6])
    SB_LUT4 i4_4_lut_adj_446 (.I0(\data_out_frame2[11] [3]), .I1(n17156), 
            .I2(\data_out_frame2[10] [7]), .I3(n6_adj_2182), .O(n10229));   // coms.v(227[16:31])
    defparam i4_4_lut_adj_446.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i150 (.Q(\data_out_frame2[18] [5]), .C(CLK_c), 
           .D(n11258));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i149 (.Q(\data_out_frame2[18] [4]), .C(CLK_c), 
           .D(n11257));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_1[[4__2244  (.Q(\data_out[1] [4]), .C(CLK_c), .D(n10908));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_adj_447 (.I0(\data_out_frame2[0] [1]), .I1(\data_out_frame2[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17294));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_447.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i148 (.Q(\data_out_frame2[18] [3]), .C(CLK_c), 
           .D(n11256));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i8_3_lut (.I0(\data_out[8][2] ), 
            .I1(\data_out[9][2] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2183));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i10_4_lut (.I0(n8_adj_2183), 
            .I1(\data_out[10] [2]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_5));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF data_out_frame2_0___i147 (.Q(\data_out_frame2[18] [2]), .C(CLK_c), 
           .D(n11255));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i146 (.Q(\data_out_frame2[18] [1]), .C(CLK_c), 
           .D(n11254));   // coms.v(416[12] 543[6])
    SB_LUT4 i2_3_lut_adj_448 (.I0(\data_out[10] [3]), .I1(n10196), .I2(\data_out[10] [7]), 
            .I3(GND_net), .O(n17243));   // coms.v(21[11:19])
    defparam i2_3_lut_adj_448.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_449 (.I0(\data_out[8][4] ), .I1(\data_out[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10392));   // coms.v(178[16:77])
    defparam i1_2_lut_adj_449.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_450 (.I0(n10440), .I1(n10229), .I2(n10346), .I3(n17165), 
            .O(n15_adj_2185));   // coms.v(228[16:596])
    defparam i6_4_lut_adj_450.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i145 (.Q(\data_out_frame2[18] [0]), .C(CLK_c), 
           .D(n11253));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i144 (.Q(\data_out_frame2[17] [7]), .C(CLK_c), 
           .D(n11252));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i143 (.Q(\data_out_frame2[17] [6]), .C(CLK_c), 
           .D(n11251));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i142 (.Q(\data_out_frame2[17] [5]), .C(CLK_c), 
           .D(n11250));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i141 (.Q(\data_out_frame2[17] [4]), .C(CLK_c), 
           .D(n11249));   // coms.v(416[12] 543[6])
    SB_DFFSS byte_transmit_counter2_i0 (.Q(byte_transmit_counter2[0]), .C(CLK_c), 
            .D(n2_adj_2186), .S(n4_adj_2187));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i140 (.Q(\data_out_frame2[17] [3]), .C(CLK_c), 
           .D(n11248));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i139 (.Q(\data_out_frame2[17] [2]), .C(CLK_c), 
           .D(n11247));   // coms.v(416[12] 543[6])
    SB_LUT4 i8_4_lut_adj_451 (.I0(n15_adj_2185), .I1(n17240), .I2(n14_adj_2188), 
            .I3(n17288), .O(n17296));   // coms.v(228[16:596])
    defparam i8_4_lut_adj_451.LUT_INIT = 16'h9669;
    SB_CARRY add_2506_3 (.CI(n16110), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n16111));
    SB_LUT4 i1_2_lut_adj_452 (.I0(\data_out[5][1] ), .I1(\data_out[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10395));   // coms.v(181[17:93])
    defparam i1_2_lut_adj_452.LUT_INIT = 16'h6666;
    SB_DFF \data_out_1[[6__2242  (.Q(\data_out[1][6] ), .C(CLK_c), .D(n10907));   // coms.v(280[12] 370[6])
    SB_LUT4 i4_4_lut_adj_453 (.I0(\data_out[10] [2]), .I1(n10395), .I2(n10392), 
            .I3(\data_out[7] [0]), .O(n10_adj_2189));   // coms.v(171[16:93])
    defparam i4_4_lut_adj_453.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_454 (.I0(n26_adj_2165), .I1(n10_adj_2189), .I2(\data_out[10] [6]), 
            .I3(GND_net), .O(data_out_9__2__N_367));   // coms.v(171[16:93])
    defparam i5_3_lut_adj_454.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_455 (.I0(\data_out[10][1] ), .I1(\data_out[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10170));   // coms.v(171[16:93])
    defparam i1_2_lut_adj_455.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i138 (.Q(\data_out_frame2[17] [1]), .C(CLK_c), 
           .D(n11246));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_1[[7__2241  (.Q(\data_out[1][7] ), .C(CLK_c), .D(n10906));   // coms.v(280[12] 370[6])
    SB_LUT4 i3_4_lut_adj_456 (.I0(\data_out_frame2[9] [2]), .I1(\data_out_frame2[7] [0]), 
            .I2(n10456), .I3(n17237), .O(n17165));   // coms.v(228[16:596])
    defparam i3_4_lut_adj_456.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_457 (.I0(n17209), .I1(n10170), .I2(data_out_9__2__N_367), 
            .I3(GND_net), .O(n17297));   // coms.v(178[16:77])
    defparam i2_3_lut_adj_457.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_458 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10259));   // coms.v(117[16:35])
    defparam i1_2_lut_adj_458.LUT_INIT = 16'h6666;
    SB_LUT4 add_977_5_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [3]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n18008), .I3(n16081), .O(\FRAME_MATCHER.i_31__N_1278 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1010_2_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n2122));   // coms.v(66[15:26])
    defparam i1010_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_459 (.I0(n10223), .I1(n10334), .I2(\data_out_frame2[5] [4]), 
            .I3(n17165), .O(n10_adj_2190));   // coms.v(228[16:596])
    defparam i4_4_lut_adj_459.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_460 (.I0(\data_out[5] [5]), .I1(\data_out[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17264));   // coms.v(184[17:86])
    defparam i1_2_lut_adj_460.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_461 (.I0(\data_out[9] [1]), .I1(n17222), .I2(\data_out[9] [7]), 
            .I3(n17243), .O(n10_adj_2191));   // coms.v(178[16:77])
    defparam i4_4_lut_adj_461.LUT_INIT = 16'h6996;
    SB_LUT4 add_2506_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(n65_adj_2192), .I3(GND_net), .O(tx_transmit_N_1947[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2506_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_462 (.I0(\data_out[6] [5]), .I1(n17264), .I2(n10_adj_2191), 
            .I3(n17297), .O(n17261));   // coms.v(171[16:355])
    defparam i1_4_lut_adj_462.LUT_INIT = 16'h6996;
    SB_CARRY add_977_5 (.CI(n16081), .I0(\FRAME_MATCHER.i [3]), .I1(n18008), 
            .CO(n16082));
    SB_DFF \data_out_2[[0__2240  (.Q(\data_out[2][0] ), .C(CLK_c), .D(n10905));   // coms.v(280[12] 370[6])
    SB_LUT4 i7_3_lut (.I0(\data_out[8][3] ), .I1(\data_out[9] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n3_adj_2193));   // coms.v(19[11:32])
    defparam i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_463 (.I0(n3_adj_2193), .I1(\data_out[10] [3]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_6));   // coms.v(19[11:32])
    defparam i8_4_lut_adj_463.LUT_INIT = 16'h0aca;
    SB_LUT4 i4_4_lut_adj_464 (.I0(\data_in_frame[2] [3]), .I1(n2122), .I2(n10215), 
            .I3(\data_in_frame[2] [5]), .O(n20_adj_2195));
    defparam i4_4_lut_adj_464.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_adj_465 (.I0(byte_transmit_counter2[5]), .I1(n11833), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2147));   // coms.v(409[11:16])
    defparam i1_2_lut_adj_465.LUT_INIT = 16'h8888;
    SB_DFF \data_out_2[[2__2238  (.Q(\data_out[2][2] ), .C(CLK_c), .D(n10904));   // coms.v(280[12] 370[6])
    SB_LUT4 i4_4_lut_adj_466 (.I0(\data_out[6] [2]), .I1(n17162), .I2(\data_out[9] [4]), 
            .I3(n17180), .O(n10_adj_2196));   // coms.v(171[16:355])
    defparam i4_4_lut_adj_466.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_467 (.I0(n17197), .I1(n10_adj_2196), .I2(n17261), 
            .I3(GND_net), .O(data_out_10__1__N_168));   // coms.v(171[16:355])
    defparam i5_3_lut_adj_467.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_468 (.I0(\data_out[6] [0]), .I1(data_out_7__2__N_447), 
            .I2(\data_out[7] [4]), .I3(GND_net), .O(n17197));   // coms.v(172[16:77])
    defparam i2_3_lut_adj_468.LUT_INIT = 16'h9696;
    SB_LUT4 select_224_Select_5_i2_4_lut (.I0(byte_transmit_counter2[5]), 
            .I1(\FRAME_MATCHER.i_31__N_1272 ), .I2(n17712), .I3(n11867), 
            .O(n2_adj_2146));
    defparam select_224_Select_5_i2_4_lut.LUT_INIT = 16'h88c0;
    SB_LUT4 i3_4_lut_adj_469 (.I0(\data_out[9] [6]), .I1(\data_out[9][2] ), 
            .I2(n10179), .I3(n17197), .O(data_out_10__2__N_157));   // coms.v(172[16:77])
    defparam i3_4_lut_adj_469.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i137 (.Q(\data_out_frame2[17] [0]), .C(CLK_c), 
           .D(n11245));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_2[[3__2237  (.Q(\data_out[2] [3]), .C(CLK_c), .D(n10903));   // coms.v(280[12] 370[6])
    SB_DFF data_out_frame2_0___i136 (.Q(\data_out_frame2[16] [7]), .C(CLK_c), 
           .D(n11244));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_2[[5__2235  (.Q(\data_out[2][5] ), .C(CLK_c), .D(n10902));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_adj_470 (.I0(\data_out_frame2[0] [0]), .I1(\data_out_frame2[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17240));
    defparam i1_2_lut_adj_470.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_471 (.I0(\data_out[7] [5]), .I1(\data_out[7] [6]), 
            .I2(\data_out[7] [7]), .I3(GND_net), .O(n10179));   // coms.v(172[16:77])
    defparam i2_3_lut_adj_471.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_472 (.I0(\data_out_frame2[10] [6]), .I1(\data_out_frame2[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17156));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_472.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i135 (.Q(\data_out_frame2[16] [6]), .C(CLK_c), 
           .D(n11243));   // coms.v(416[12] 543[6])
    SB_LUT4 i3_4_lut_adj_473 (.I0(data_out_7__3__N_441), .I1(\data_out[6] [1]), 
            .I2(\data_out[8]_c [0]), .I3(n10179), .O(n17147));   // coms.v(21[11:19])
    defparam i3_4_lut_adj_473.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i134 (.Q(\data_out_frame2[16] [5]), .C(CLK_c), 
           .D(n11242));   // coms.v(416[12] 543[6])
    SB_LUT4 i4_4_lut_adj_474 (.I0(\data_out_frame2[9] [3]), .I1(\data_out_frame2[16] [7]), 
            .I2(\data_out_frame2[15] [7]), .I3(n6_adj_2197), .O(n17123));
    defparam i4_4_lut_adj_474.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_475 (.I0(n17147), .I1(\data_out[9] [7]), .I2(\data_out[9] [3]), 
            .I3(GND_net), .O(data_out_10__3__N_146));   // coms.v(21[11:19])
    defparam i2_3_lut_adj_475.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_476 (.I0(\data_out_frame2[7] [5]), .I1(\data_out_frame2[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10346));   // coms.v(229[16:299])
    defparam i1_2_lut_adj_476.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i133 (.Q(\data_out_frame2[16] [4]), .C(CLK_c), 
           .D(n11241));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_adj_477 (.I0(\data_out_frame2[16] [1]), .I1(\data_out_frame2[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10468));   // coms.v(230[16:237])
    defparam i1_2_lut_adj_477.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_478 (.I0(\data_out_frame2[16] [3]), .I1(\data_out_frame2[6] [3]), 
            .I2(\data_out_frame2[13] [7]), .I3(GND_net), .O(n17285));   // coms.v(228[16:596])
    defparam i2_3_lut_adj_478.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_479 (.I0(\data_out[6] [2]), .I1(\data_out[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10447));   // coms.v(170[16:355])
    defparam i1_2_lut_adj_479.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i8_3_lut (.I0(\data_out[8][4] ), 
            .I1(\data_out[9] [4]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2198));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_4_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame2_0___i132 (.Q(\data_out_frame2[16] [3]), .C(CLK_c), 
           .D(n11240));   // coms.v(416[12] 543[6])
    SB_LUT4 i7_4_lut_adj_480 (.I0(\data_in_frame[0] [7]), .I1(n2138), .I2(\data_in_frame[1] [1]), 
            .I3(\data_in_frame[1] [7]), .O(n23));
    defparam i7_4_lut_adj_480.LUT_INIT = 16'hde7b;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i10_4_lut (.I0(n8_adj_2198), 
            .I1(\data_out[10] [4]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_7));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_4_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_977_4_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [2]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n18008), .I3(n16080), .O(\FRAME_MATCHER.i_31__N_1278 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i12_4_lut_adj_481 (.I0(n17291), .I1(n17309), .I2(n17303), 
            .I3(n17315), .O(n28_adj_2200));   // coms.v(228[16:596])
    defparam i12_4_lut_adj_481.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15341 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [7]), .I2(\data_out_frame2[15] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18136));
    defparam byte_transmit_counter2_0__bdd_4_lut_15341.LUT_INIT = 16'he4aa;
    SB_CARRY add_2506_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(n65_adj_2192), 
            .CO(n16110));
    SB_DFF data_out_frame2_0___i131 (.Q(\data_out_frame2[16] [2]), .C(CLK_c), 
           .D(n11239));   // coms.v(416[12] 543[6])
    SB_LUT4 i11_4_lut_adj_482 (.I0(\data_in_frame[1] [2]), .I1(n22_adj_2201), 
            .I2(\data_in_frame[2] [2]), .I3(n10259), .O(n27_adj_2202));
    defparam i11_4_lut_adj_482.LUT_INIT = 16'hdffd;
    SB_LUT4 i10_4_lut (.I0(n10513), .I1(n17153), .I2(\data_out_frame2[5] [7]), 
            .I3(n17168), .O(n26_adj_2203));   // coms.v(228[16:596])
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_483 (.I0(n17194), .I1(n17231), .I2(n17216), 
            .I3(n17285), .O(n27_adj_2204));   // coms.v(228[16:596])
    defparam i11_4_lut_adj_483.LUT_INIT = 16'h6996;
    SB_CARRY add_977_4 (.CI(n16080), .I0(\FRAME_MATCHER.i [2]), .I1(n18008), 
            .CO(n16081));
    SB_LUT4 add_977_3_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [1]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(n18008), .I3(n16079), .O(\FRAME_MATCHER.i_31__N_1278 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i9_4_lut_adj_484 (.I0(\data_out_frame2[5] [1]), .I1(\data_out_frame2[6] [7]), 
            .I2(n10520), .I3(\data_out_frame2[6] [0]), .O(n25));   // coms.v(228[16:596])
    defparam i9_4_lut_adj_484.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27_adj_2204), .I2(n26_adj_2203), 
            .I3(n28_adj_2200), .O(n10223));   // coms.v(228[16:596])
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_485 (.I0(n17177), .I1(\data_out[7] [6]), .I2(n10183), 
            .I3(GND_net), .O(data_out_10__4__N_135));   // coms.v(174[16:77])
    defparam i2_3_lut_adj_485.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame2_0___i130 (.Q(\data_out_frame2[16] [1]), .C(CLK_c), 
           .D(n11238));   // coms.v(416[12] 543[6])
    SB_LUT4 add_977_33_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [31]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n18008), .I3(n16109), .O(\FRAME_MATCHER.i_31__N_1278 [31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_33_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i6_4_lut_adj_486 (.I0(\data_out_frame2[12] [5]), .I1(n10263), 
            .I2(\data_out_frame2[12] [7]), .I3(n17123), .O(n15_adj_2205));
    defparam i6_4_lut_adj_486.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_487 (.I0(n15_adj_2205), .I1(n17156), .I2(n14_adj_2206), 
            .I3(n17240), .O(n17275));
    defparam i8_4_lut_adj_487.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame2_0___i129 (.Q(\data_out_frame2[16] [0]), .C(CLK_c), 
           .D(n11237));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i128 (.Q(\data_out_frame2[15] [7]), .C(CLK_c), 
           .D(n11236));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_adj_488 (.I0(\data_out_frame2[13] [4]), .I1(\data_out_frame2[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17315));   // coms.v(228[16:596])
    defparam i1_2_lut_adj_488.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_489 (.I0(\data_out[8]_c [0]), .I1(\data_out[8][1] ), 
            .I2(\data_out[7] [7]), .I3(GND_net), .O(n10183));   // coms.v(174[16:77])
    defparam i2_3_lut_adj_489.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_490 (.I0(\data_out[6] [3]), .I1(\data_out[6] [1]), 
            .I2(n10183), .I3(GND_net), .O(n17180));   // coms.v(175[16:77])
    defparam i2_3_lut_adj_490.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_491 (.I0(n2137), .I1(n2120), .I2(\data_in_frame[2] [1]), 
            .I3(\data_in_frame[2] [4]), .O(n18));
    defparam i2_4_lut_adj_491.LUT_INIT = 16'hb7ed;
    SB_LUT4 i15155_2_lut (.I0(\data_out[1] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17701));
    defparam i15155_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame2_0___i127 (.Q(\data_out_frame2[15] [6]), .C(CLK_c), 
           .D(n11235));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i126 (.Q(\data_out_frame2[15] [5]), .C(CLK_c), 
           .D(n11234));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i125 (.Q(\data_out_frame2[15] [4]), .C(CLK_c), 
           .D(n11233));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i124 (.Q(\data_out_frame2[15] [3]), .C(CLK_c), 
           .D(n11232));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i123 (.Q(\data_out_frame2[15] [2]), .C(CLK_c), 
           .D(n11231));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i122 (.Q(\data_out_frame2[15] [1]), .C(CLK_c), 
           .D(n11230));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i121 (.Q(\data_out_frame2[15] [0]), .C(CLK_c), 
           .D(n11229));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i120 (.Q(\data_out_frame2[14] [7]), .C(CLK_c), 
           .D(n11228));   // coms.v(416[12] 543[6])
    SB_DFFE delay_counter_2361__i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n10594), 
            .D(n61[13]));   // coms.v(305[16] 313[10])
    SB_LUT4 add_977_32_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [30]), .I1(\FRAME_MATCHER.i [30]), 
            .I2(n18008), .I3(n16108), .O(\FRAME_MATCHER.i_31__N_1278 [30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_32_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i2_3_lut (.I0(\data_out[2][2] ), 
            .I1(\data_out[3][2] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2145));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_977_3 (.CI(n16079), .I0(\FRAME_MATCHER.i [1]), .I1(n18008), 
            .CO(n16080));
    SB_LUT4 add_977_2_lut (.I0(n37), .I1(\FRAME_MATCHER.i [0]), .I2(n18008), 
            .I3(VCC_net), .O(\FRAME_MATCHER.i_31__N_1278 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i8360_3_lut_4_lut (.I0(n15171), .I1(n17072), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n11046));
    defparam i8360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15015_3_lut (.I0(\data_out_frame2[0] [0]), .I1(byte_transmit_counter2[1]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n17603));
    defparam i15015_3_lut.LUT_INIT = 16'h3232;
    SB_DFF data_out_frame2_0___i119 (.Q(\data_out_frame2[14] [6]), .C(CLK_c), 
           .D(n11227));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i118 (.Q(\data_out_frame2[14] [5]), .C(CLK_c), 
           .D(n11226));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i117 (.Q(\data_out_frame2[14] [4]), .C(CLK_c), 
           .D(n11225));   // coms.v(416[12] 543[6])
    SB_LUT4 i4_4_lut_adj_492 (.I0(\data_out_frame2[7] [6]), .I1(n10424), 
            .I2(\data_out_frame2[7] [3]), .I3(\data_out_frame2[9] [2]), 
            .O(n10_adj_2207));   // coms.v(230[16:237])
    defparam i4_4_lut_adj_492.LUT_INIT = 16'h6996;
    SB_DFFE delay_counter_2361__i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n10594), 
            .D(n61[12]));   // coms.v(305[16] 313[10])
    SB_DFFE delay_counter_2361__i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n10594), 
            .D(n61[11]));   // coms.v(305[16] 313[10])
    SB_DFF data_out_frame2_0___i116 (.Q(\data_out_frame2[14] [3]), .C(CLK_c), 
           .D(n11224));   // coms.v(416[12] 543[6])
    SB_DFFE delay_counter_2361__i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n10594), 
            .D(n61[10]));   // coms.v(305[16] 313[10])
    SB_DFFE delay_counter_2361__i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n10594), 
            .D(n61[9]));   // coms.v(305[16] 313[10])
    SB_DFFE delay_counter_2361__i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n10594), 
            .D(n61[8]));   // coms.v(305[16] 313[10])
    SB_CARRY add_977_2 (.CI(VCC_net), .I0(\FRAME_MATCHER.i [0]), .I1(n18008), 
            .CO(n16079));
    SB_DFFE delay_counter_2361__i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n10594), 
            .D(n61[7]));   // coms.v(305[16] 313[10])
    SB_LUT4 i2_3_lut_adj_493 (.I0(n17252), .I1(\data_out[10][1] ), .I2(\data_out[8][2] ), 
            .I3(GND_net), .O(data_out_10__5__N_124));   // coms.v(175[16:77])
    defparam i2_3_lut_adj_493.LUT_INIT = 16'h9696;
    SB_DFFE delay_counter_2361__i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n10594), 
            .D(n61[6]));   // coms.v(305[16] 313[10])
    SB_LUT4 i3_4_lut_adj_494 (.I0(\data_out_frame2[8] [0]), .I1(\data_out_frame2[7] [4]), 
            .I2(\data_out_frame2[15] [4]), .I3(n17174), .O(n10356));   // coms.v(234[16:291])
    defparam i3_4_lut_adj_494.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i115 (.Q(\data_out_frame2[14] [2]), .C(CLK_c), 
           .D(n11223));   // coms.v(416[12] 543[6])
    SB_DFFE delay_counter_2361__i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n10594), 
            .D(n61[5]));   // coms.v(305[16] 313[10])
    SB_LUT4 i10_4_lut_adj_495 (.I0(n2128), .I1(n20_adj_2195), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[1] [0]), .O(n26_adj_2210));
    defparam i10_4_lut_adj_495.LUT_INIT = 16'hefdf;
    SB_DFFE delay_counter_2361__i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n10594), 
            .D(n61[4]));   // coms.v(305[16] 313[10])
    SB_DFFE delay_counter_2361__i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n10594), 
            .D(n61[3]));   // coms.v(305[16] 313[10])
    SB_DFFE delay_counter_2361__i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n10594), 
            .D(n61[2]));   // coms.v(305[16] 313[10])
    SB_DFFE delay_counter_2361__i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n10594), 
            .D(n61[1]));   // coms.v(305[16] 313[10])
    SB_CARRY add_977_32 (.CI(n16108), .I0(\FRAME_MATCHER.i [30]), .I1(n18008), 
            .CO(n16109));
    SB_LUT4 delay_counter_2361_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[13]), .I3(n16078), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame2_0___i114 (.Q(\data_out_frame2[14] [1]), .C(CLK_c), 
           .D(n11222));   // coms.v(416[12] 543[6])
    SB_LUT4 delay_counter_2361_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[12]), .I3(n16077), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_496 (.I0(\data_out_frame2[5] [5]), .I1(\data_out_frame2[9] [3]), 
            .I2(n10356), .I3(GND_net), .O(n17184));   // coms.v(232[16:229])
    defparam i2_3_lut_adj_496.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut (.I0(n27_adj_2202), .I1(n23), .I2(\data_in_frame[1] [3]), 
            .I3(\data_in_frame[1] [4]), .O(n30_adj_2213));
    defparam i14_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_adj_497 (.I0(\data_out[9] [6]), .I1(\data_out[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17209));   // coms.v(176[16:77])
    defparam i1_2_lut_adj_497.LUT_INIT = 16'h6666;
    SB_LUT4 add_977_31_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [29]), .I1(\FRAME_MATCHER.i [29]), 
            .I2(n18008), .I3(n16107), .O(\FRAME_MATCHER.i_31__N_1278 [29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_31_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_4_lut_adj_498 (.I0(n2138), .I1(n2124), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[2] [6]), .O(n17_adj_2214));
    defparam i1_4_lut_adj_498.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_adj_499 (.I0(\data_out_frame2[0] [5]), .I1(\data_out_frame2[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17219));   // coms.v(380[12:27])
    defparam i1_2_lut_adj_499.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_500 (.I0(\data_out_frame2[0] [2]), .I1(\data_out_frame2[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2215));   // coms.v(380[12:27])
    defparam i1_2_lut_adj_500.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_501 (.I0(\data_out[8]_c [0]), .I1(\data_out[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2216));   // coms.v(176[16:77])
    defparam i1_2_lut_adj_501.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i113 (.Q(\data_out_frame2[14] [0]), .C(CLK_c), 
           .D(n11221));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i112 (.Q(\data_out_frame2[13] [7]), .C(CLK_c), 
           .D(n11220));   // coms.v(416[12] 543[6])
    SB_LUT4 i4_4_lut_adj_502 (.I0(\data_out_frame2[0] [1]), .I1(n17219), 
            .I2(n17107), .I3(n6_adj_2215), .O(n10263));   // coms.v(380[12:27])
    defparam i4_4_lut_adj_502.LUT_INIT = 16'h6996;
    SB_CARRY add_977_31 (.CI(n16107), .I0(\FRAME_MATCHER.i [29]), .I1(n18008), 
            .CO(n16108));
    SB_LUT4 i1_2_lut_adj_503 (.I0(\data_out_frame2[13] [0]), .I1(n10263), 
            .I2(GND_net), .I3(GND_net), .O(n17246));   // coms.v(228[16:596])
    defparam i1_2_lut_adj_503.LUT_INIT = 16'h6666;
    SB_CARRY delay_counter_2361_add_4_14 (.CI(n16077), .I0(GND_net), .I1(n76[12]), 
            .CO(n16078));
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame2[6] [0]), 
            .I1(\data_out_frame2[7] [0]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2217));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_504 (.I0(\data_out_frame2[15] [6]), .I1(\data_out_frame2[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17300));   // coms.v(230[16:237])
    defparam i1_2_lut_adj_504.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_505 (.I0(\data_out_frame2[5] [7]), .I1(\data_out_frame2[0] [0]), 
            .I2(\data_out_frame2[13] [6]), .I3(\data_out_frame2[13] [1]), 
            .O(n30_adj_2218));   // coms.v(230[16:237])
    defparam i11_4_lut_adj_505.LUT_INIT = 16'h6996;
    SB_DFF \data_out_2[[7__2233  (.Q(\data_out[2][7] ), .C(CLK_c), .D(n10901));   // coms.v(280[12] 370[6])
    SB_DFF data_out_frame2_0___i111 (.Q(\data_out_frame2[13] [6]), .C(CLK_c), 
           .D(n11219));   // coms.v(416[12] 543[6])
    SB_LUT4 delay_counter_2361_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[11]), .I3(n16076), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8217_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10596), .I3(\data_out[2] [3]), .O(n10903));
    defparam i8217_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_LUT4 i4_4_lut_adj_506 (.I0(\data_out[6] [2]), .I1(n17209), .I2(n10188), 
            .I3(n6_adj_2216), .O(data_out_10__6__N_113));   // coms.v(176[16:77])
    defparam i4_4_lut_adj_506.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_507 (.I0(n17300), .I1(n30_adj_2218), .I2(\data_out_frame2[10] [6]), 
            .I3(\data_out_frame2[5] [6]), .O(n34));   // coms.v(230[16:237])
    defparam i15_4_lut_adj_507.LUT_INIT = 16'h6996;
    SB_DFF \data_out_3[[0__2232  (.Q(\data_out[3][0] ), .C(CLK_c), .D(n10900));   // coms.v(280[12] 370[6])
    SB_DFF data_out_frame2_0___i110 (.Q(\data_out_frame2[13] [5]), .C(CLK_c), 
           .D(n11218));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_3[[2__2230  (.Q(\data_out[3][2] ), .C(CLK_c), .D(n10899));   // coms.v(280[12] 370[6])
    SB_DFF data_out_frame2_0___i109 (.Q(\data_out_frame2[13] [4]), .C(CLK_c), 
           .D(n11217));   // coms.v(416[12] 543[6])
    SB_LUT4 i13_4_lut (.I0(n17116), .I1(n17171), .I2(n17132), .I3(n17184), 
            .O(n32));   // coms.v(230[16:237])
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY delay_counter_2361_add_4_13 (.CI(n16076), .I0(GND_net), .I1(n76[11]), 
            .CO(n16077));
    SB_LUT4 i8222_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10596), .I3(\data_out[1] [4]), .O(n10908));
    defparam i8222_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_LUT4 i6_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(n10705));
    defparam i6_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i14_4_lut_adj_508 (.I0(n17187), .I1(n17246), .I2(n17228), 
            .I3(n17267), .O(n33));   // coms.v(230[16:237])
    defparam i14_4_lut_adj_508.LUT_INIT = 16'h6996;
    SB_LUT4 delay_counter_2361_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[10]), .I3(n16075), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF \data_out_3[[4__2228  (.Q(\data_out[3][4] ), .C(CLK_c), .D(n10898));   // coms.v(280[12] 370[6])
    SB_LUT4 i12_4_lut_adj_509 (.I0(\data_out_frame2[6] [6]), .I1(n10563), 
            .I2(\data_out_frame2[13] [5]), .I3(n17095), .O(n31_c));   // coms.v(230[16:237])
    defparam i12_4_lut_adj_509.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_510 (.I0(n31_c), .I1(n33), .I2(n32), .I3(n34), 
            .O(n17301));   // coms.v(230[16:237])
    defparam i18_4_lut_adj_510.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i108 (.Q(\data_out_frame2[13] [3]), .C(CLK_c), 
           .D(n11216));   // coms.v(416[12] 543[6])
    SB_LUT4 i8361_3_lut_4_lut (.I0(n15171), .I1(n17072), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n11047));
    defparam i8361_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame2_0___i107 (.Q(\data_out_frame2[13] [2]), .C(CLK_c), 
           .D(n11215));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_adj_511 (.I0(\data_out_frame2[5] [2]), .I1(\data_out_frame2[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10456));   // coms.v(228[16:596])
    defparam i1_2_lut_adj_511.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_512 (.I0(\data_out[6] [3]), .I1(\data_out[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2221));   // coms.v(179[16:84])
    defparam i1_2_lut_adj_512.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_513 (.I0(\data_out_frame2[11] [0]), .I1(\data_out_frame2[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17279));   // coms.v(228[16:596])
    defparam i1_2_lut_adj_513.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_514 (.I0(\data_out[6] [5]), .I1(\data_out[9] [7]), 
            .I2(n10188), .I3(n6_adj_2221), .O(n17110));   // coms.v(179[16:84])
    defparam i4_4_lut_adj_514.LUT_INIT = 16'h6996;
    SB_LUT4 add_977_30_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [28]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(n18008), .I3(n16106), .O(\FRAME_MATCHER.i_31__N_1278 [28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_30_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY delay_counter_2361_add_4_12 (.CI(n16075), .I0(GND_net), .I1(n76[10]), 
            .CO(n16076));
    SB_LUT4 i1_2_lut_adj_515 (.I0(\data_out_frame2[12] [3]), .I1(\data_out_frame2[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n10548));   // coms.v(241[17:248])
    defparam i1_2_lut_adj_515.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i106 (.Q(\data_out_frame2[13] [1]), .C(CLK_c), 
           .D(n11214));   // coms.v(416[12] 543[6])
    SB_LUT4 i8224_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10596), .I3(\data_out[0] [6]), .O(n10910));
    defparam i8224_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_DFF data_out_frame2_0___i105 (.Q(\data_out_frame2[13] [0]), .C(CLK_c), 
           .D(n11213));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i104 (.Q(\data_out_frame2[12] [7]), .C(CLK_c), 
           .D(n11212));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_adj_516 (.I0(\data_out_frame2[13] [6]), .I1(\data_out_frame2[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10530));   // coms.v(233[16:291])
    defparam i1_2_lut_adj_516.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut_adj_517 (.I0(n17_adj_2214), .I1(n30_adj_2213), .I2(n26_adj_2210), 
            .I3(n18), .O(n31));
    defparam i15_4_lut_adj_517.LUT_INIT = 16'hfffe;
    SB_LUT4 delay_counter_2361_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[9]), .I3(n16074), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut_adj_518 (.I0(n10456), .I1(n10504), .I2(\data_out_frame2[8] [4]), 
            .I3(n10492), .O(n20_adj_2223));   // coms.v(228[16:596])
    defparam i8_4_lut_adj_518.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_519 (.I0(\data_out[8][4] ), .I1(n17110), .I2(GND_net), 
            .I3(GND_net), .O(data_out_10__7__N_101));   // coms.v(179[16:84])
    defparam i1_2_lut_adj_519.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_520 (.I0(n10530), .I1(\data_out_frame2[7] [2]), 
            .I2(\data_out_frame2[9] [1]), .I3(n10548), .O(n19_adj_2224));   // coms.v(228[16:596])
    defparam i7_4_lut_adj_520.LUT_INIT = 16'h6996;
    SB_LUT4 n18136_bdd_4_lut (.I0(n18136), .I1(\data_out_frame2[13] [7]), 
            .I2(\data_out_frame2[12] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n18139));
    defparam n18136_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_521 (.I0(n17135), .I1(n17279), .I2(n17225), .I3(n17309), 
            .O(n21));   // coms.v(228[16:596])
    defparam i9_4_lut_adj_521.LUT_INIT = 16'h6996;
    SB_LUT4 i8362_3_lut_4_lut (.I0(n15171), .I1(n17072), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n11048));
    defparam i8362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame2[5] [0]), 
            .I1(n5_adj_2217), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2143));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i11_3_lut (.I0(n21), .I1(n19_adj_2224), .I2(n20_adj_2223), 
            .I3(GND_net), .O(n17310));   // coms.v(228[16:596])
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_CARRY add_977_30 (.CI(n16106), .I0(\FRAME_MATCHER.i [28]), .I1(n18008), 
            .CO(n16107));
    SB_CARRY delay_counter_2361_add_4_11 (.CI(n16074), .I0(GND_net), .I1(n76[9]), 
            .CO(n16075));
    SB_LUT4 i1_2_lut_adj_522 (.I0(\data_out_frame2[9] [0]), .I1(\data_out_frame2[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10504));   // coms.v(229[16:299])
    defparam i1_2_lut_adj_522.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_523 (.I0(\data_out_frame2[10] [5]), .I1(\data_out_frame2[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10428));   // coms.v(229[16:299])
    defparam i1_2_lut_adj_523.LUT_INIT = 16'h6666;
    SB_LUT4 i15202_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10596), .I3(GND_net), .O(n10595));
    defparam i15202_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_2225), .S(n3_adj_2226));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_3_i3_2_lut_3_lut (.I0(n13146), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n10009), .I3(GND_net), .O(n3_adj_2227));
    defparam select_219_Select_3_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i10673_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [15]));   // coms.v(430[13] 433[7])
    defparam i10673_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1014_2_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n2126));   // coms.v(68[15:26])
    defparam i1014_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_524 (.I0(\data_out_frame2[16] [4]), .I1(\data_out_frame2[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10572));   // coms.v(242[17:884])
    defparam i1_2_lut_adj_524.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_525 (.I0(\data_out_frame2[11] [7]), .I1(\data_out_frame2[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17141));   // coms.v(233[16:291])
    defparam i1_2_lut_adj_525.LUT_INIT = 16'h6666;
    SB_LUT4 i15074_3_lut (.I0(\data_out_frame2[0] [1]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17587));
    defparam i15074_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i3_4_lut_adj_526 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(n10215), .O(n17206));   // coms.v(76[16:62])
    defparam i3_4_lut_adj_526.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_527 (.I0(\data_out_frame2[8] [4]), .I1(\data_out_frame2[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2228));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_527.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i103 (.Q(\data_out_frame2[12] [6]), .C(CLK_c), 
           .D(n11211));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_2229), .S(n3_adj_2230));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_2231), .S(n3_adj_2232));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_2233), .S(n3_adj_2234));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_2235), .S(n3_adj_2236));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_2237), .S(n3_adj_2238));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_2239), .S(n3_adj_2240));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_2241), .S(n3_adj_2242));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_2243), .S(n3_adj_2244));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_2245), .S(n3_adj_2246));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_2247), .S(n3_adj_2248));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i102 (.Q(\data_out_frame2[12] [5]), .C(CLK_c), 
           .D(n11210));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i101 (.Q(\data_out_frame2[12] [4]), .C(CLK_c), 
           .D(n11209));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_2249), .S(n3_adj_2250));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_2251), .S(n3_adj_2252));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_2253), .S(n3_adj_2254));   // coms.v(416[12] 543[6])
    SB_LUT4 add_977_29_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [27]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(n18008), .I3(n16105), .O(\FRAME_MATCHER.i_31__N_1278 [27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_29_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i15122_2_lut (.I0(\data_out[0][5] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17622));
    defparam i15122_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 delay_counter_2361_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[8]), .I3(n16073), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2510_9_lut (.I0(tx2_transmit_N_1996), .I1(byte_transmit_counter2[7]), 
            .I2(GND_net), .I3(n15978), .O(n17714)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_9_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_2256), .S(n3_adj_2257));   // coms.v(416[12] 543[6])
    SB_CARRY delay_counter_2361_add_4_10 (.CI(n16073), .I0(GND_net), .I1(n76[8]), 
            .CO(n16074));
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_2258), .S(n3_adj_2259));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_2260), .S(n3_adj_2261));   // coms.v(416[12] 543[6])
    SB_CARRY add_977_29 (.CI(n16105), .I0(\FRAME_MATCHER.i [27]), .I1(n18008), 
            .CO(n16106));
    SB_LUT4 add_977_28_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [26]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(n18008), .I3(n16104), .O(\FRAME_MATCHER.i_31__N_1278 [26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_28_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 delay_counter_2361_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[7]), .I3(n16072), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_2263), .S(n3_adj_2264));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_2265), .S(n3_adj_2266));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_2267), .S(n3_adj_2268));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2_adj_2269), .S(n3_adj_2270));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_2271), .S(n3_adj_2272));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_2273), .S(n3_adj_2274));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_2275), .S(n3_adj_2276));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_2277), .S(n3_adj_2278));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_2279), .S(n3_adj_2280));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_2281), .S(n3_adj_2282));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_2283), .S(n3_adj_2179));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_2284), .S(n3_adj_2227));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_2285), .S(n3_adj_2286));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_2287), .S(n3_adj_2288));   // coms.v(416[12] 543[6])
    SB_LUT4 i4_4_lut_adj_528 (.I0(\data_out_frame2[5] [2]), .I1(n17312), 
            .I2(n10572), .I3(n6_adj_2228), .O(n17116));   // coms.v(227[16:31])
    defparam i4_4_lut_adj_528.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i100 (.Q(\data_out_frame2[12] [3]), .C(CLK_c), 
           .D(n11208));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15288 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [3]), .I2(\data_out_frame2[11] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n18064));
    defparam byte_transmit_counter2_0__bdd_4_lut_15288.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame2_0___i99 (.Q(\data_out_frame2[12] [2]), .C(CLK_c), 
           .D(n11207));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i98 (.Q(\data_out_frame2[12] [1]), .C(CLK_c), 
           .D(n11206));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i97 (.Q(\data_out_frame2[12] [0]), .C(CLK_c), 
           .D(n11205));   // coms.v(416[12] 543[6])
    SB_LUT4 n18064_bdd_4_lut (.I0(n18064), .I1(\data_out_frame2[9] [3]), 
            .I2(\data_out_frame2[8] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n18067));
    defparam n18064_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame2[6] [1]), 
            .I1(\data_out_frame2[7] [1]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2289));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_529 (.I0(\data_out_frame2[5] [0]), .I1(\data_out_frame2[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10554));   // coms.v(241[17:248])
    defparam i1_2_lut_adj_529.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15279 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [3]), .I2(\data_out_frame2[15] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n18058));
    defparam byte_transmit_counter2_0__bdd_4_lut_15279.LUT_INIT = 16'he4aa;
    SB_LUT4 n18058_bdd_4_lut (.I0(n18058), .I1(\data_out_frame2[13] [3]), 
            .I2(\data_out_frame2[12] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n18061));
    defparam n18058_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut (.I0(\data_out_frame2[5] [1]), 
            .I1(n5_adj_2289), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2142));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_DFF data_out_frame2_0___i96 (.Q(\data_out_frame2[11] [7]), .C(CLK_c), 
           .D(n11204));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i2_3_lut (.I0(\data_out[2][5] ), 
            .I1(\data_out[3][5] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2164));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_530 (.I0(\data_out_frame2[13] [5]), .I1(\data_out_frame2[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10520));   // coms.v(232[16:229])
    defparam i1_2_lut_adj_530.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15274 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [3]), .I2(\data_out_frame2[19] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n18052));
    defparam byte_transmit_counter2_0__bdd_4_lut_15274.LUT_INIT = 16'he4aa;
    SB_LUT4 n18052_bdd_4_lut (.I0(n18052), .I1(\data_out_frame2[17] [3]), 
            .I2(\data_out_frame2[16] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n18055));
    defparam n18052_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out[6] [2]), 
            .I1(\data_out[7] [2]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2141));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15269 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [2]), .I2(\data_out_frame2[11] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n18046));
    defparam byte_transmit_counter2_0__bdd_4_lut_15269.LUT_INIT = 16'he4aa;
    SB_LUT4 n18046_bdd_4_lut (.I0(n18046), .I1(\data_out_frame2[9] [2]), 
            .I2(\data_out_frame2[8] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n18049));
    defparam n18046_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame2_0___i95 (.Q(\data_out_frame2[11] [6]), .C(CLK_c), 
           .D(n11203));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i94 (.Q(\data_out_frame2[11] [5]), .C(CLK_c), 
           .D(n11202));   // coms.v(416[12] 543[6])
    SB_LUT4 i15088_2_lut (.I0(\data_out[5] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17671));
    defparam i15088_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10672_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [16]));   // coms.v(430[13] 433[7])
    defparam i10672_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15264 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [2]), .I2(\data_out_frame2[15] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n18040));
    defparam byte_transmit_counter2_0__bdd_4_lut_15264.LUT_INIT = 16'he4aa;
    SB_LUT4 n18040_bdd_4_lut (.I0(n18040), .I1(\data_out_frame2[13] [2]), 
            .I2(\data_out_frame2[12] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n18043));
    defparam n18040_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6489_2_lut (.I0(byte_transmit_counter2[0]), .I1(byte_transmit_counter2[1]), 
            .I2(GND_net), .I3(GND_net), .O(n9157));   // coms.v(403[36:58])
    defparam i6489_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15371 (.I0(byte_transmit_counter2[2]), 
            .I1(n17568), .I2(n17569), .I3(byte_transmit_counter2[3]), 
            .O(n18034));
    defparam byte_transmit_counter2_2__bdd_4_lut_15371.LUT_INIT = 16'he4aa;
    SB_LUT4 n18034_bdd_4_lut (.I0(n18034), .I1(n17440), .I2(n17439), .I3(byte_transmit_counter2[3]), 
            .O(n18037));
    defparam n18034_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_977_28 (.CI(n16104), .I0(\FRAME_MATCHER.i [26]), .I1(n18008), 
            .CO(n16105));
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15259 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [2]), .I2(\data_out_frame2[19] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n18028));
    defparam byte_transmit_counter2_0__bdd_4_lut_15259.LUT_INIT = 16'he4aa;
    SB_LUT4 n18028_bdd_4_lut (.I0(n18028), .I1(\data_out_frame2[17] [2]), 
            .I2(\data_out_frame2[16] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n18031));
    defparam n18028_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY delay_counter_2361_add_4_9 (.CI(n16072), .I0(GND_net), .I1(n76[7]), 
            .CO(n16073));
    SB_DFF data_out_frame2_0___i93 (.Q(\data_out_frame2[11] [4]), .C(CLK_c), 
           .D(n11201));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15250 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [1]), .I2(\data_out_frame2[11] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n18022));
    defparam byte_transmit_counter2_0__bdd_4_lut_15250.LUT_INIT = 16'he4aa;
    SB_LUT4 n18022_bdd_4_lut (.I0(n18022), .I1(\data_out_frame2[9] [1]), 
            .I2(\data_out_frame2[8] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n18025));
    defparam n18022_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame2[6] [2]), 
            .I1(\data_out_frame2[7] [2]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2290));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15245 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [1]), .I2(\data_out_frame2[15] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n18016));
    defparam byte_transmit_counter2_0__bdd_4_lut_15245.LUT_INIT = 16'he4aa;
    SB_LUT4 add_2510_8_lut (.I0(tx2_transmit_N_1996), .I1(byte_transmit_counter2[6]), 
            .I2(GND_net), .I3(n15977), .O(n17713)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n18016_bdd_4_lut (.I0(n18016), .I1(\data_out_frame2[13] [1]), 
            .I2(\data_out_frame2[12] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n18019));
    defparam n18016_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_2510_7_lut (.I0(tx2_transmit_N_1996), .I1(byte_transmit_counter2[5]), 
            .I2(GND_net), .I3(n15976), .O(n17712)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2510_7 (.CI(n15976), .I0(byte_transmit_counter2[5]), .I1(GND_net), 
            .CO(n15977));
    SB_CARRY add_2510_6 (.CI(n15975), .I0(byte_transmit_counter2[4]), .I1(GND_net), 
            .CO(n15976));
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame2[5] [2]), 
            .I1(n5_adj_2290), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2140));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 add_2510_5_lut (.I0(tx2_transmit_N_1996), .I1(byte_transmit_counter2[3]), 
            .I2(GND_net), .I3(n15974), .O(n17711)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15240 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [1]), .I2(\data_out_frame2[19] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n18010));
    defparam byte_transmit_counter2_0__bdd_4_lut_15240.LUT_INIT = 16'he4aa;
    SB_LUT4 add_2510_4_lut (.I0(tx2_transmit_N_1996), .I1(byte_transmit_counter2[2]), 
            .I2(GND_net), .I3(n15973), .O(n17710)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n18010_bdd_4_lut (.I0(n18010), .I1(\data_out_frame2[17] [1]), 
            .I2(\data_out_frame2[16] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n18013));
    defparam n18010_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame2_0___i92 (.Q(\data_out_frame2[11] [3]), .C(CLK_c), 
           .D(n11200));   // coms.v(416[12] 543[6])
    SB_CARRY add_2510_3 (.CI(n15972), .I0(byte_transmit_counter2[1]), .I1(GND_net), 
            .CO(n15973));
    SB_DFF data_out_frame2_0___i91 (.Q(\data_out_frame2[11] [2]), .C(CLK_c), 
           .D(n11199));   // coms.v(416[12] 543[6])
    SB_LUT4 add_2510_2_lut (.I0(tx2_transmit_N_1996), .I1(byte_transmit_counter2[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n17659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8363_3_lut_4_lut (.I0(n15171), .I1(n17072), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n11049));
    defparam i8363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_2510_8 (.CI(n15977), .I0(byte_transmit_counter2[6]), .I1(GND_net), 
            .CO(n15978));
    SB_LUT4 add_2510_6_lut (.I0(tx2_transmit_N_1996), .I1(byte_transmit_counter2[4]), 
            .I2(GND_net), .I3(n15975), .O(n17606)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2510_5 (.CI(n15974), .I0(byte_transmit_counter2[3]), .I1(GND_net), 
            .CO(n15975));
    SB_CARRY add_2510_4 (.CI(n15973), .I0(byte_transmit_counter2[2]), .I1(GND_net), 
            .CO(n15974));
    SB_DFF data_out_frame2_0___i90 (.Q(\data_out_frame2[11] [1]), .C(CLK_c), 
           .D(n11198));   // coms.v(416[12] 543[6])
    SB_LUT4 i6_4_lut_adj_531 (.I0(n10554), .I1(n17116), .I2(\data_out_frame2[8] [3]), 
            .I3(n17234), .O(n15_adj_2291));   // coms.v(227[16:31])
    defparam i6_4_lut_adj_531.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_532 (.I0(n15_adj_2291), .I1(n17249), .I2(n14_adj_2292), 
            .I3(n17255), .O(n17290));   // coms.v(227[16:31])
    defparam i8_4_lut_adj_532.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame2_0___i89 (.Q(\data_out_frame2[11] [0]), .C(CLK_c), 
           .D(n11197));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i88 (.Q(\data_out_frame2[10] [7]), .C(CLK_c), 
           .D(n11196));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i87 (.Q(\data_out_frame2[10] [6]), .C(CLK_c), 
           .D(n11195));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15336 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [7]), .I2(\data_out_frame2[19] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18130));
    defparam byte_transmit_counter2_0__bdd_4_lut_15336.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame2_0___i86 (.Q(\data_out_frame2[10] [5]), .C(CLK_c), 
           .D(n11194));   // coms.v(416[12] 543[6])
    SB_LUT4 n18130_bdd_4_lut (.I0(n18130), .I1(\data_out_frame2[17] [7]), 
            .I2(\data_out_frame2[16] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n18133));
    defparam n18130_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_533 (.I0(\data_out_frame2[16] [3]), .I1(\data_out_frame2[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n10482));   // coms.v(240[17:239])
    defparam i1_2_lut_adj_533.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i85 (.Q(\data_out_frame2[10] [4]), .C(CLK_c), 
           .D(n11193));   // coms.v(416[12] 543[6])
    SB_LUT4 add_977_27_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [25]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(n18008), .I3(n16103), .O(\FRAME_MATCHER.i_31__N_1278 [25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_27_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i10610_3_lut (.I0(byte_transmit_counter2[2]), .I1(byte_transmit_counter2[4]), 
            .I2(byte_transmit_counter2[3]), .I3(GND_net), .O(n13284));
    defparam i10610_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1016_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2128));   // coms.v(69[15:26])
    defparam i1016_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_977_27 (.CI(n16103), .I0(\FRAME_MATCHER.i [25]), .I1(n18008), 
            .CO(n16104));
    SB_DFF data_out_frame2_0___i84 (.Q(\data_out_frame2[10] [3]), .C(CLK_c), 
           .D(n11192));   // coms.v(416[12] 543[6])
    SB_LUT4 add_977_26_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [24]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(n18008), .I3(n16102), .O(\FRAME_MATCHER.i_31__N_1278 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_26_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i6_4_lut_adj_534 (.I0(n10507), .I1(\data_out_frame2[11] [6]), 
            .I2(\data_out_frame2[7] [0]), .I3(\data_out_frame2[14] [4]), 
            .O(n16_adj_2293));   // coms.v(239[17:230])
    defparam i6_4_lut_adj_534.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i83 (.Q(\data_out_frame2[10] [2]), .C(CLK_c), 
           .D(n11191));   // coms.v(416[12] 543[6])
    SB_LUT4 i7_4_lut_adj_535 (.I0(\data_out_frame2[13] [4]), .I1(n17135), 
            .I2(n17092), .I3(n17228), .O(n17_adj_2294));   // coms.v(239[17:230])
    defparam i7_4_lut_adj_535.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_536 (.I0(n17_adj_2294), .I1(n17282), .I2(n16_adj_2293), 
            .I3(n17312), .O(n17313));   // coms.v(239[17:230])
    defparam i9_4_lut_adj_536.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_537 (.I0(byte_transmit_counter2[6]), .I1(byte_transmit_counter2[7]), 
            .I2(byte_transmit_counter2[5]), .I3(n13284), .O(n13628));
    defparam i3_4_lut_adj_537.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame2_0___i82 (.Q(\data_out_frame2[10] [1]), .C(CLK_c), 
           .D(n11190));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i81 (.Q(\data_out_frame2[10] [0]), .C(CLK_c), 
           .D(n11189));   // coms.v(416[12] 543[6])
    SB_LUT4 i8364_3_lut_4_lut (.I0(n15171), .I1(n17072), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n11050));
    defparam i8364_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10493_2_lut (.I0(tx2_active), .I1(r_SM_Main_2__N_2034_adj_2405[0]), 
            .I2(GND_net), .I3(GND_net), .O(n11867));
    defparam i10493_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_538 (.I0(\data_out_frame2[12] [2]), .I1(\data_out_frame2[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17092));   // coms.v(228[16:596])
    defparam i1_2_lut_adj_538.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i80 (.Q(\data_out_frame2[9] [7]), .C(CLK_c), 
           .D(n11188));   // coms.v(416[12] 543[6])
    SB_CARRY add_977_26 (.CI(n16102), .I0(\FRAME_MATCHER.i [24]), .I1(n18008), 
            .CO(n16103));
    SB_LUT4 i8365_3_lut_4_lut (.I0(n15171), .I1(n17072), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n11051));
    defparam i8365_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_539 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10215));   // coms.v(76[16:62])
    defparam i1_2_lut_adj_539.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i79 (.Q(\data_out_frame2[9] [6]), .C(CLK_c), 
           .D(n11187));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [4]), .O(n16784));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_540 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [5]), .O(n7));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_540.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_541 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [6]), .O(n7_adj_2295));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_541.LUT_INIT = 16'hea00;
    SB_DFF data_out_frame2_0___i78 (.Q(\data_out_frame2[9] [5]), .C(CLK_c), 
           .D(n11186));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_3[[5__2227  (.Q(\data_out[3][5] ), .C(CLK_c), .D(n10897));   // coms.v(280[12] 370[6])
    SB_LUT4 i6_4_lut_adj_542 (.I0(n10533), .I1(n10334), .I2(n10507), .I3(\data_out_frame2[6] [3]), 
            .O(n14_adj_2296));   // coms.v(238[17:230])
    defparam i6_4_lut_adj_542.LUT_INIT = 16'h6996;
    SB_LUT4 i8366_3_lut_4_lut (.I0(n15171), .I1(n17072), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n11052));
    defparam i8366_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_543 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17213));   // coms.v(130[17:124])
    defparam i1_2_lut_adj_543.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_544 (.I0(\data_out_frame2[13] [3]), .I1(n14_adj_2296), 
            .I2(n10_adj_2297), .I3(\data_out_frame2[9] [7]), .O(n17171));   // coms.v(238[17:230])
    defparam i7_4_lut_adj_544.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_545 (.I0(\data_out_frame2[14] [3]), .I1(\data_out_frame2[8] [1]), 
            .I2(\data_out_frame2[8] [5]), .I3(n17171), .O(n12_adj_2298));   // coms.v(238[17:230])
    defparam i5_4_lut_adj_545.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_546 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17101));   // coms.v(505[9:81])
    defparam i1_2_lut_adj_546.LUT_INIT = 16'h6666;
    SB_LUT4 i8357_3_lut_4_lut (.I0(n39), .I1(n17076), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n11043));
    defparam i8357_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14591_2_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n10018), .I2(GND_net), 
            .I3(GND_net), .O(n17367));
    defparam i14591_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_547 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[0] [7]), .I3(n17101), .O(n10_adj_2299));   // coms.v(505[9:81])
    defparam i4_4_lut_adj_547.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_548 (.I0(n17249), .I1(n12_adj_2298), .I2(\data_out_frame2[6] [7]), 
            .I3(n10437), .O(n17250));   // coms.v(238[17:230])
    defparam i6_4_lut_adj_548.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_549 (.I0(\data_out_frame2[16] [0]), .I1(\data_out_frame2[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17168));   // coms.v(237[17:221])
    defparam i1_2_lut_adj_549.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_550 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [7]), .O(n7_adj_2300));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_550.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_adj_551 (.I0(\data_out_frame2[6] [6]), .I1(\data_out_frame2[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10472));   // coms.v(241[17:248])
    defparam i1_2_lut_adj_551.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_552 (.I0(n13146), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(GND_net), .O(n43));
    defparam i1_2_lut_adj_552.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15331 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [6]), .I2(\data_out_frame2[11] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n18124));
    defparam byte_transmit_counter2_0__bdd_4_lut_15331.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_553 (.I0(\data_out_frame2[10] [0]), .I1(\data_out_frame2[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10462));   // coms.v(239[17:230])
    defparam i1_2_lut_adj_553.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_554 (.I0(\data_in_frame[1] [3]), .I1(n10_adj_2299), 
            .I2(n17206), .I3(\data_in_frame[1] [2]), .O(n10407));   // coms.v(505[9:81])
    defparam i5_4_lut_adj_554.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_555 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [8]), .O(n16782));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_555.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_adj_556 (.I0(\data_out_frame2[16] [1]), .I1(\data_out_frame2[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10533));   // coms.v(238[17:230])
    defparam i1_2_lut_adj_556.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_557 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [9]), .O(n16766));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_557.LUT_INIT = 16'hea00;
    SB_DFF \data_out_3[[6__2226  (.Q(\data_out[3] [6]), .C(CLK_c), .D(n10896));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_4_lut_adj_558 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [10]), .O(n16780));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_558.LUT_INIT = 16'hea00;
    SB_DFF \data_out_3[[7__2225  (.Q(\data_out[3][7] ), .C(CLK_c), .D(n10895));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_4_lut_adj_559 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [11]), .O(n7_adj_2301));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_559.LUT_INIT = 16'hea00;
    SB_DFF data_out_frame2_0___i77 (.Q(\data_out_frame2[9] [4]), .C(CLK_c), 
           .D(n11185));   // coms.v(416[12] 543[6])
    SB_LUT4 i10750_2_lut_4_lut (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [12]), .O(n13426));   // coms.v(412[11:12])
    defparam i10750_2_lut_4_lut.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_560 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [13]), .O(n7_adj_2302));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_560.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_adj_561 (.I0(\FRAME_MATCHER.state[0] ), .I1(n488), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_2174));
    defparam i1_2_lut_adj_561.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_562 (.I0(n2124), .I1(n2120), .I2(\data_in_frame[3] [6]), 
            .I3(\data_in_frame[3] [4]), .O(n19_adj_2303));
    defparam i5_4_lut_adj_562.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_563 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [6]), 
            .I2(n10407), .I3(\data_in_frame[6] [1]), .O(n17114));   // coms.v(505[9:81])
    defparam i2_4_lut_adj_563.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out[6] [5]), 
            .I1(\data_out[7] [5]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2163));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_564 (.I0(\data_out_frame2[8] [1]), .I1(\data_out_frame2[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17132));   // coms.v(237[17:221])
    defparam i1_2_lut_adj_564.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_565 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [14]), .O(n7_adj_2304));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_565.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_566 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [15]), .O(n7_adj_2305));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_566.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_567 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [16]), .O(n16768));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_567.LUT_INIT = 16'hea00;
    SB_DFF data_out_frame2_0___i76 (.Q(\data_out_frame2[9] [3]), .C(CLK_c), 
           .D(n11184));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i75 (.Q(\data_out_frame2[9] [2]), .C(CLK_c), 
           .D(n11183));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i74 (.Q(\data_out_frame2[9] [1]), .C(CLK_c), 
           .D(n11182));   // coms.v(416[12] 543[6])
    SB_LUT4 i15104_2_lut (.I0(\data_out[5] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17581));
    defparam i15104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_977_25_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [23]), .I1(\FRAME_MATCHER.i [23]), 
            .I2(n18008), .I3(n16101), .O(\FRAME_MATCHER.i_31__N_1278 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_25_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_4_lut_adj_568 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [17]), .O(n16764));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_568.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_569 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [18]), .O(n7_adj_2306));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_569.LUT_INIT = 16'hea00;
    SB_DFF data_out_frame2_0___i73 (.Q(\data_out_frame2[9] [0]), .C(CLK_c), 
           .D(n11181));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_4_lut_adj_570 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [19]), .O(n7_adj_2307));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_570.LUT_INIT = 16'hea00;
    SB_LUT4 n18124_bdd_4_lut (.I0(n18124), .I1(\data_out_frame2[9] [6]), 
            .I2(\data_out_frame2[8] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n18127));
    defparam n18124_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_adj_571 (.I0(n17282), .I1(n10371), .I2(\data_out_frame2[14] [2]), 
            .I3(GND_net), .O(n14_adj_2308));   // coms.v(237[17:221])
    defparam i5_3_lut_adj_571.LUT_INIT = 16'h9696;
    SB_LUT4 i8367_3_lut_4_lut (.I0(n15171), .I1(n17072), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n11053));
    defparam i8367_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_572 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [20]), .O(n7_adj_2309));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_572.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_573 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [21]), .O(n16760));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_573.LUT_INIT = 16'hea00;
    SB_LUT4 i1_4_lut_adj_574 (.I0(n2137), .I1(\data_in_frame[3] [3]), .I2(\data_in_frame[3] [1]), 
            .I3(n10215), .O(n15_adj_2310));
    defparam i1_4_lut_adj_574.LUT_INIT = 16'hb7ed;
    SB_LUT4 i1_2_lut_4_lut_adj_575 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [22]), .O(n16758));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_575.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_576 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [23]), .O(n7_adj_2311));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_576.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_577 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [24]), .O(n16756));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_577.LUT_INIT = 16'hea00;
    SB_LUT4 i6_4_lut_adj_578 (.I0(n10533), .I1(n10462), .I2(n10472), .I3(n17098), 
            .O(n15_adj_2312));   // coms.v(237[17:221])
    defparam i6_4_lut_adj_578.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_579 (.I0(n13146), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(GND_net), .O(n41));
    defparam i1_2_lut_adj_579.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_580 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [25]), .O(n16754));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_580.LUT_INIT = 16'hea00;
    SB_DFF data_out_frame2_0___i72 (.Q(\data_out_frame2[8] [7]), .C(CLK_c), 
           .D(n11180));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_4_lut_adj_581 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [26]), .O(n16752));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_581.LUT_INIT = 16'hea00;
    SB_LUT4 i8_4_lut_adj_582 (.I0(n15_adj_2312), .I1(n17203), .I2(n14_adj_2308), 
            .I3(n17267), .O(n17284));   // coms.v(237[17:221])
    defparam i8_4_lut_adj_582.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_583 (.I0(n276), .I1(\FRAME_MATCHER.i_31__N_1275 ), 
            .I2(n9369), .I3(\FRAME_MATCHER.state [27]), .O(n16750));   // coms.v(412[11:12])
    defparam i1_2_lut_4_lut_adj_583.LUT_INIT = 16'hea00;
    SB_LUT4 delay_counter_2361_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[6]), .I3(n16071), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out[5] [3]), .I1(\data_out[5] [4]), 
            .I2(data_out_7__3__N_441), .I3(GND_net), .O(n17129));   // coms.v(115[16:67])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_CARRY add_977_25 (.CI(n16101), .I0(\FRAME_MATCHER.i [23]), .I1(n18008), 
            .CO(n16102));
    SB_CARRY delay_counter_2361_add_4_8 (.CI(n16071), .I0(GND_net), .I1(n76[6]), 
            .CO(n16072));
    SB_LUT4 add_2510_3_lut (.I0(tx2_transmit_N_1996), .I1(byte_transmit_counter2[1]), 
            .I2(GND_net), .I3(n15972), .O(n17589)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2510_2 (.CI(VCC_net), .I0(byte_transmit_counter2[0]), .I1(GND_net), 
            .CO(n15972));
    SB_LUT4 delay_counter_2361_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[5]), .I3(n16070), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_977_24_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [22]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(n18008), .I3(n16100), .O(\FRAME_MATCHER.i_31__N_1278 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_24_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_584 (.I0(\data_out_frame2[8] [4]), .I1(\data_out_frame2[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10513));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_584.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i71 (.Q(\data_out_frame2[8] [6]), .C(CLK_c), 
           .D(n11179));   // coms.v(416[12] 543[6])
    SB_LUT4 i2_3_lut_adj_585 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[5] [3]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n16475));   // coms.v(505[9:81])
    defparam i2_3_lut_adj_585.LUT_INIT = 16'h9696;
    SB_LUT4 select_219_Select_14_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [14]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2264));   // coms.v(430[13] 433[7])
    defparam select_219_Select_14_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i14662_3_lut (.I0(byte_transmit_counter2[0]), .I1(byte_transmit_counter2[1]), 
            .I2(\data_out_frame2[0] [4]), .I3(GND_net), .O(n17439));
    defparam i14662_3_lut.LUT_INIT = 16'h9898;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame2[6] [4]), 
            .I1(\data_out_frame2[7] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2315));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_586 (.I0(\data_out_frame2[9] [5]), .I1(\data_out_frame2[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17187));   // coms.v(234[16:291])
    defparam i1_2_lut_adj_586.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_587 (.I0(n2126), .I1(n2138), .I2(\data_in_frame[3] [7]), 
            .I3(\data_in_frame[3] [0]), .O(n18_adj_2316));
    defparam i4_4_lut_adj_587.LUT_INIT = 16'h7bde;
    SB_LUT4 i8358_3_lut_4_lut (.I0(n39), .I1(n17076), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n11044));
    defparam i8358_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame2_0___i70 (.Q(\data_out_frame2[8] [5]), .C(CLK_c), 
           .D(n11178));   // coms.v(416[12] 543[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out[5] [3]), .I1(\data_out[5] [4]), 
            .I2(data_out_7__2__N_447), .I3(n10326), .O(n17126));   // coms.v(115[16:67])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_219_Select_2_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2286));   // coms.v(430[13] 433[7])
    defparam select_219_Select_2_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_adj_588 (.I0(n13146), .I1(\FRAME_MATCHER.i [0]), 
            .I2(n10009), .I3(GND_net), .O(n3_adj_2181));
    defparam i1_2_lut_3_lut_adj_588.LUT_INIT = 16'h0808;
    SB_LUT4 i14663_4_lut (.I0(\data_out_frame2[5] [4]), .I1(n5_adj_2315), 
            .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n17440));
    defparam i14663_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i10_4_lut_adj_589 (.I0(n19_adj_2303), .I1(\data_in_frame[2] [3]), 
            .I2(n17373), .I3(\data_in_frame[2] [4]), .O(n24_adj_2317));
    defparam i10_4_lut_adj_589.LUT_INIT = 16'hbfff;
    SB_LUT4 select_219_Select_1_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2288));   // coms.v(430[13] 433[7])
    defparam select_219_Select_1_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_CARRY add_977_24 (.CI(n16100), .I0(\FRAME_MATCHER.i [22]), .I1(n18008), 
            .CO(n16101));
    SB_LUT4 i1_2_lut_adj_590 (.I0(\data_out_frame2[13] [1]), .I1(\data_out_frame2[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17273));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_590.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_591 (.I0(\data_out_frame2[16] [5]), .I1(\data_out_frame2[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2318));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_591.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_592 (.I0(n10359), .I1(n10349), .I2(\data_out_frame2[10] [3]), 
            .I3(n6_adj_2318), .O(n17216));   // coms.v(227[16:31])
    defparam i4_4_lut_adj_592.LUT_INIT = 16'h6996;
    SB_LUT4 add_977_23_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [21]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(n18008), .I3(n16099), .O(\FRAME_MATCHER.i_31__N_1278 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_23_lut.LUT_INIT = 16'hA3AC;
    SB_DFFE \data_out_10[[7__2169  (.Q(\data_out[10] [7]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__7__N_101));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_adj_593 (.I0(\data_out_frame2[12] [0]), .I1(\data_out_frame2[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10413));   // coms.v(238[17:230])
    defparam i1_2_lut_adj_593.LUT_INIT = 16'h6666;
    SB_CARRY delay_counter_2361_add_4_7 (.CI(n16070), .I0(GND_net), .I1(n76[5]), 
            .CO(n16071));
    SB_DFFE \data_out_10[[6__2170  (.Q(\data_out[10] [6]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__6__N_113));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_10[[5__2171  (.Q(\data_out[10] [5]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__5__N_124));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_10[[4__2172  (.Q(\data_out[10] [4]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__4__N_135));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_10[[3__2173  (.Q(\data_out[10] [3]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__3__N_146));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_10[[2__2174  (.Q(\data_out[10] [2]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__2__N_157));   // coms.v(280[12] 370[6])
    SB_LUT4 select_219_Select_31_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [31]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2226));   // coms.v(430[13] 433[7])
    defparam select_219_Select_31_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFFE \data_out_10[[1__2175  (.Q(\data_out[10][1] ), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__1__N_168));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_10[[0__2176  (.Q(\data_out[10][0] ), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__0__N_219));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_9[[7__2177  (.Q(\data_out[9] [7]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__7__N_272));   // coms.v(280[12] 370[6])
    SB_DFF data_out_frame2_0___i1 (.Q(\data_out_frame2[0] [0]), .C(CLK_c), 
           .D(n17492));   // coms.v(416[12] 543[6])
    SB_CARRY add_977_23 (.CI(n16099), .I0(\FRAME_MATCHER.i [21]), .I1(n18008), 
            .CO(n16100));
    SB_DFFE \data_out_9[[6__2178  (.Q(\data_out[9] [6]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__6__N_324));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_9[[5__2179  (.Q(\data_out[9] [5]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__5__N_334));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_9[[4__2180  (.Q(\data_out[9] [4]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__4__N_344));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_9[[3__2181  (.Q(\data_out[9] [3]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__3__N_356));   // coms.v(280[12] 370[6])
    SB_DFFE \data_out_9[[1__2183  (.Q(\data_out[9] [1]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__1__N_378));   // coms.v(280[12] 370[6])
    SB_LUT4 select_219_Select_30_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [30]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2230));   // coms.v(430[13] 433[7])
    defparam select_219_Select_30_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mux_1195_i1_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(n2698[0]));   // coms.v(283[4] 369[11])
    defparam mux_1195_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \data_out_9[[0__2184  (.Q(\data_out[9] [0]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__0__N_389));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_adj_594 (.I0(\data_out_frame2[16] [7]), .I1(n17194), 
            .I2(GND_net), .I3(GND_net), .O(n10459));   // coms.v(238[17:230])
    defparam i1_2_lut_adj_594.LUT_INIT = 16'h6666;
    SB_LUT4 select_219_Select_29_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [29]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2232));   // coms.v(430[13] 433[7])
    defparam select_219_Select_29_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i8_4_lut_adj_595 (.I0(n15_adj_2310), .I1(\data_in_frame[2] [6]), 
            .I2(n2138), .I3(\data_in_frame[2] [7]), .O(n22_adj_2319));
    defparam i8_4_lut_adj_595.LUT_INIT = 16'hfbbf;
    SB_DFF data_out_frame2_0___i69 (.Q(\data_out_frame2[8] [4]), .C(CLK_c), 
           .D(n11177));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i68 (.Q(\data_out_frame2[8] [3]), .C(CLK_c), 
           .D(n11176));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i67 (.Q(\data_out_frame2[8] [2]), .C(CLK_c), 
           .D(n11175));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i66 (.Q(\data_out_frame2[8] [1]), .C(CLK_c), 
           .D(n11174));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i65 (.Q(\data_out_frame2[8] [0]), .C(CLK_c), 
           .D(n11173));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i64 (.Q(\data_out_frame2[7] [7]), .C(CLK_c), 
           .D(n11172));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i63 (.Q(\data_out_frame2[7] [6]), .C(CLK_c), 
           .D(n11171));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i62 (.Q(\data_out_frame2[7] [5]), .C(CLK_c), 
           .D(n11170));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i61 (.Q(\data_out_frame2[7] [4]), .C(CLK_c), 
           .D(n11169));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i60 (.Q(\data_out_frame2[7] [3]), .C(CLK_c), 
           .D(n11168));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i59 (.Q(\data_out_frame2[7] [2]), .C(CLK_c), 
           .D(n11167));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i58 (.Q(\data_out_frame2[7] [1]), .C(CLK_c), 
           .D(n11166));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i57 (.Q(\data_out_frame2[7] [0]), .C(CLK_c), 
           .D(n11165));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i56 (.Q(\data_out_frame2[6] [7]), .C(CLK_c), 
           .D(n11164));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i55 (.Q(\data_out_frame2[6] [6]), .C(CLK_c), 
           .D(n11163));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i54 (.Q(\data_out_frame2[6] [5]), .C(CLK_c), 
           .D(n11162));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i53 (.Q(\data_out_frame2[6] [4]), .C(CLK_c), 
           .D(n11161));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i52 (.Q(\data_out_frame2[6] [3]), .C(CLK_c), 
           .D(n11160));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i51 (.Q(\data_out_frame2[6] [2]), .C(CLK_c), 
           .D(n11159));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i50 (.Q(\data_out_frame2[6] [1]), .C(CLK_c), 
           .D(n11158));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i49 (.Q(\data_out_frame2[6] [0]), .C(CLK_c), 
           .D(n11157));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i48 (.Q(\data_out_frame2[5] [7]), .C(CLK_c), 
           .D(n11156));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i47 (.Q(\data_out_frame2[5] [6]), .C(CLK_c), 
           .D(n11155));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i46 (.Q(\data_out_frame2[5] [5]), .C(CLK_c), 
           .D(n11154));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i45 (.Q(\data_out_frame2[5] [4]), .C(CLK_c), 
           .D(n11153));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i44 (.Q(\data_out_frame2[5] [3]), .C(CLK_c), 
           .D(n11152));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i43 (.Q(\data_out_frame2[5] [2]), .C(CLK_c), 
           .D(n11151));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i42 (.Q(\data_out_frame2[5] [1]), .C(CLK_c), 
           .D(n11150));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i41 (.Q(\data_out_frame2[5] [0]), .C(CLK_c), 
           .D(n11149));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_7[[5__2195  (.Q(\data_out[7] [5]), .C(CLK_c), .D(n11079));   // coms.v(280[12] 370[6])
    SB_DFF \data_out_7[[6__2194  (.Q(\data_out[7] [6]), .C(CLK_c), .D(n11084));   // coms.v(280[12] 370[6])
    SB_DFF \data_out_7[[7__2193  (.Q(\data_out[7] [7]), .C(CLK_c), .D(n11146));   // coms.v(280[12] 370[6])
    SB_LUT4 i6_4_lut_adj_596 (.I0(\data_out_frame2[0] [7]), .I1(\data_out_frame2[14] [1]), 
            .I2(n10563), .I3(\data_out_frame2[12] [1]), .O(n16_adj_2320));   // coms.v(227[16:31])
    defparam i6_4_lut_adj_596.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(CLK_c), 
            .D(n16740), .S(n16700));   // coms.v(416[12] 543[6])
    SB_LUT4 i7_4_lut_adj_597 (.I0(\data_out_frame2[16] [0]), .I1(\data_out_frame2[8] [3]), 
            .I2(n10459), .I3(n17098), .O(n17_adj_2321));   // coms.v(227[16:31])
    defparam i7_4_lut_adj_597.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_598 (.I0(n17_adj_2321), .I1(n17216), .I2(n16_adj_2320), 
            .I3(n17273), .O(n17274));   // coms.v(227[16:31])
    defparam i9_4_lut_adj_598.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_599 (.I0(\data_out_frame2[11] [6]), .I1(\data_out_frame2[11] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10437));   // coms.v(238[17:230])
    defparam i1_2_lut_adj_599.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(CLK_c), 
            .D(n16744), .S(n16698));   // coms.v(416[12] 543[6])
    SB_LUT4 i10681_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [7]));   // coms.v(430[13] 433[7])
    defparam i10681_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut_adj_600 (.I0(\data_in_frame[2] [2]), .I1(n18_adj_2316), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[2] [1]), .O(n23_adj_2322));
    defparam i9_4_lut_adj_600.LUT_INIT = 16'hdffd;
    SB_LUT4 i7_4_lut_adj_601 (.I0(n2122), .I1(\data_in_frame[3] [2]), .I2(\data_in_frame[3] [5]), 
            .I3(n10259), .O(n21_adj_2323));
    defparam i7_4_lut_adj_601.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_602 (.I0(n2128), .I1(n2126), .I2(\data_in_frame[5] [0]), 
            .I3(\data_in_frame[6] [7]), .O(n19_adj_2324));
    defparam i3_4_lut_adj_602.LUT_INIT = 16'h7bde;
    SB_LUT4 i13_4_lut_adj_603 (.I0(n21_adj_2323), .I1(n23_adj_2322), .I2(n22_adj_2319), 
            .I3(n24_adj_2317), .O(n4494));
    defparam i13_4_lut_adj_603.LUT_INIT = 16'hfffe;
    SB_LUT4 select_219_Select_28_i3_2_lut_3_lut (.I0(n13146), .I1(\FRAME_MATCHER.i [28]), 
            .I2(n10009), .I3(GND_net), .O(n3_adj_2234));
    defparam select_219_Select_28_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i15170_3_lut (.I0(\data_out_frame2[0] [3]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17761));
    defparam i15170_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i2_4_lut_adj_604 (.I0(n17213), .I1(\data_in_frame[6] [0]), .I2(\data_in_frame[1] [5]), 
            .I3(n10407), .O(n17215));   // coms.v(130[17:124])
    defparam i2_4_lut_adj_604.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_605 (.I0(byte_transmit_counter2[6]), .I1(n11833), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2325));   // coms.v(409[11:16])
    defparam i1_2_lut_adj_605.LUT_INIT = 16'h8888;
    SB_LUT4 select_219_Select_1_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [1]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2287));
    defparam select_219_Select_1_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10680_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [8]));   // coms.v(430[13] 433[7])
    defparam i10680_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_224_Select_6_i2_4_lut (.I0(byte_transmit_counter2[6]), 
            .I1(\FRAME_MATCHER.i_31__N_1272 ), .I2(n17713), .I3(n11867), 
            .O(n2_adj_2326));
    defparam select_224_Select_6_i2_4_lut.LUT_INIT = 16'h88c0;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(CLK_c), 
            .D(n16746), .S(n16658));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(CLK_c), 
            .D(n16748), .S(n16696));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(CLK_c), 
            .D(n16750), .S(n16718));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(CLK_c), 
            .D(n16752), .S(n16702));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(CLK_c), 
            .D(n16754), .S(n16690));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(CLK_c), 
            .D(n16756), .S(n16688));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(CLK_c), 
            .D(n7_adj_2311), .S(n13381));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(CLK_c), 
            .D(n16758), .S(n16714));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(CLK_c), 
            .D(n16760), .S(n16686));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(CLK_c), 
            .D(n7_adj_2309), .S(n8_adj_2327));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(CLK_c), 
            .D(n7_adj_2307), .S(n8_adj_2328));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(CLK_c), 
            .D(n7_adj_2306), .S(n8_adj_2329));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(CLK_c), 
            .D(n16764), .S(n16704));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(CLK_c), 
            .D(n16768), .S(n16670));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(CLK_c), 
            .D(n7_adj_2305), .S(n8_adj_2330));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(CLK_c), 
            .D(n7_adj_2304), .S(n8_adj_2331));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(CLK_c), 
            .D(n7_adj_2302), .S(n8_adj_2332));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(CLK_c), 
            .D(n13426), .S(n16708));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(CLK_c), 
            .D(n7_adj_2301), .S(n8_adj_2333));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(CLK_c), 
            .D(n16780), .S(n16710));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(CLK_c), 
            .D(n16766), .S(n16674));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(CLK_c), 
            .D(n16782), .S(n16666));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(CLK_c), 
            .D(n7_adj_2300), .S(n16141));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(CLK_c), 
            .D(n7_adj_2295), .S(n8_adj_2334));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(CLK_c), 
            .D(n7), .S(n8_adj_2335));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(CLK_c), 
            .D(n16784), .S(n16716));   // coms.v(416[12] 543[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(CLK_c), 
            .D(n18285), .S(n6_adj_2336));   // coms.v(416[12] 543[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state[1] ), .C(CLK_c), 
           .D(n18286));   // coms.v(416[12] 543[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state[2] ), .C(CLK_c), 
           .D(n18287));   // coms.v(416[12] 543[6])
    SB_LUT4 i10679_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [9]));   // coms.v(430[13] 433[7])
    defparam i10679_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14615_2_lut_4_lut (.I0(n444), .I1(n16267), .I2(n9453), .I3(\UART_TRANSMITTER.state[2] ), 
            .O(n17392));
    defparam i14615_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame2[6] [3]), 
            .I1(\data_out_frame2[7] [3]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2337));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10678_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [10]));   // coms.v(430[13] 433[7])
    defparam i10678_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame2[5] [3]), 
            .I1(n5_adj_2337), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2139));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_adj_606 (.I0(\data_out_frame2[12] [0]), .I1(\data_out_frame2[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10434));   // coms.v(234[16:291])
    defparam i1_2_lut_adj_606.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_607 (.I0(n444), .I1(n16267), .I2(n9453), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n4));
    defparam i1_2_lut_4_lut_adj_607.LUT_INIT = 16'h00fb;
    SB_LUT4 i15151_3_lut (.I0(\data_out_frame2[0] [5]), .I1(byte_transmit_counter2[1]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n17678));
    defparam i15151_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i10677_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [11]));   // coms.v(430[13] 433[7])
    defparam i10677_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_608 (.I0(\data_out_frame2[16] [6]), .I1(\data_out_frame2[15] [6]), 
            .I2(\data_out_frame2[14] [0]), .I3(GND_net), .O(n17237));   // coms.v(235[16:291])
    defparam i2_3_lut_adj_608.LUT_INIT = 16'h9696;
    SB_DFF \data_out_8[[2__2190  (.Q(\data_out[8][2] ), .C(CLK_c), .D(n11132));   // coms.v(280[12] 370[6])
    SB_LUT4 i2_3_lut_adj_609 (.I0(\data_out_frame2[10] [2]), .I1(\data_out_frame2[16] [4]), 
            .I2(\data_out_frame2[12] [1]), .I3(GND_net), .O(n10492));   // coms.v(241[17:248])
    defparam i2_3_lut_adj_609.LUT_INIT = 16'h9696;
    SB_LUT4 select_219_Select_2_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [2]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2285));
    defparam select_219_Select_2_i2_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \data_in_3[[7__2262  (.Q(\data_in[3] [7]), .C(CLK_c), .D(n11131));   // coms.v(416[12] 543[6])
    SB_DFF \data_out_8[[3__2189  (.Q(\data_out[8][3] ), .C(CLK_c), .D(n11130));   // coms.v(280[12] 370[6])
    SB_LUT4 i10676_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [12]));   // coms.v(430[13] 433[7])
    defparam i10676_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \data_out_8[[4__2188  (.Q(\data_out[8][4] ), .C(CLK_c), .D(n11129));   // coms.v(280[12] 370[6])
    SB_LUT4 i4_4_lut_adj_610 (.I0(\data_out_frame2[10] [0]), .I1(\data_out_frame2[8] [2]), 
            .I2(n10492), .I3(n6_adj_2339), .O(n17153));   // coms.v(228[16:596])
    defparam i4_4_lut_adj_610.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_611 (.I0(\data_in_frame[5] [6]), .I1(n17215), .I2(\data_in_frame[1] [4]), 
            .I3(\data_in_frame[1] [5]), .O(n24_adj_2340));
    defparam i8_4_lut_adj_611.LUT_INIT = 16'hb77b;
    SB_DFF \data_out_8[[5__2187  (.Q(\data_out[8][5] ), .C(CLK_c), .D(n11128));   // coms.v(280[12] 370[6])
    SB_DFF \data_out_8[[6__2186  (.Q(\data_out[8][6] ), .C(CLK_c), .D(n11127));   // coms.v(280[12] 370[6])
    SB_DFF \data_out_8[[7__2185  (.Q(\data_out[8] [7]), .C(CLK_c), .D(n11126));   // coms.v(280[12] 370[6])
    SB_DFF \data_in_3[[6__2263  (.Q(\data_in[3] [6]), .C(CLK_c), .D(n11125));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_adj_612 (.I0(\data_out_frame2[0] [7]), .I1(\data_out_frame2[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17107));   // coms.v(380[12:27])
    defparam i1_2_lut_adj_612.LUT_INIT = 16'h6666;
    SB_DFF \data_out_9[[2__2182  (.Q(\data_out[9][2] ), .C(CLK_c), .D(n11124));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_adj_613 (.I0(\data_out_frame2[15] [7]), .I1(\data_out_frame2[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10563));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_613.LUT_INIT = 16'h6666;
    SB_DFF \data_out_8[[1__2191  (.Q(\data_out[8][1] ), .C(CLK_c), .D(n11123));   // coms.v(280[12] 370[6])
    SB_LUT4 i3_4_lut_adj_614 (.I0(\data_out_frame2[9] [4]), .I1(\data_out_frame2[6] [0]), 
            .I2(\data_out_frame2[7] [7]), .I3(\data_out_frame2[9] [6]), 
            .O(n10424));   // coms.v(231[16:291])
    defparam i3_4_lut_adj_614.LUT_INIT = 16'h6996;
    SB_DFF \data_out_8[[0__2192  (.Q(\data_out[8]_c [0]), .C(CLK_c), .D(n11122));   // coms.v(280[12] 370[6])
    SB_DFF \data_in_3[[5__2264  (.Q(\data_in[3] [5]), .C(CLK_c), .D(n11121));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_3[[4__2265  (.Q(\data_in[3] [4]), .C(CLK_c), .D(n11120));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_27_i3_2_lut_3_lut (.I0(n13146), .I1(\FRAME_MATCHER.i [27]), 
            .I2(n10009), .I3(GND_net), .O(n3_adj_2236));
    defparam select_219_Select_27_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i10675_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [13]));   // coms.v(430[13] 433[7])
    defparam i10675_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_219_Select_26_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [26]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2238));   // coms.v(430[13] 433[7])
    defparam select_219_Select_26_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_25_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [25]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2240));   // coms.v(430[13] 433[7])
    defparam select_219_Select_25_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i6_4_lut_adj_615 (.I0(\data_out_frame2[11] [7]), .I1(n10424), 
            .I2(n10563), .I3(\data_out_frame2[13] [0]), .O(n15_adj_2341));   // coms.v(235[16:291])
    defparam i6_4_lut_adj_615.LUT_INIT = 16'h6996;
    SB_LUT4 i15080_3_lut (.I0(\data_out_frame2[0] [6]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17620));
    defparam i15080_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 delay_counter_2361_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[4]), .I3(n16069), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame2[6] [6]), 
            .I1(\data_out_frame2[7] [6]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2343));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS byte_transmit_counter2_i7 (.Q(byte_transmit_counter2[7]), .C(CLK_c), 
            .D(n2_adj_2344), .S(n4_adj_2345));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_24_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [24]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2242));   // coms.v(430[13] 433[7])
    defparam select_219_Select_24_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut (.I0(\data_out_frame2[5] [6]), 
            .I1(n5_adj_2343), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2161));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i2_3_lut_adj_616 (.I0(n17072), .I1(\FRAME_MATCHER.i [2]), .I2(\FRAME_MATCHER.i [0]), 
            .I3(GND_net), .O(n17075));
    defparam i2_3_lut_adj_616.LUT_INIT = 16'hfbfb;
    SB_LUT4 i8_4_lut_adj_617 (.I0(n15_adj_2341), .I1(n17107), .I2(n14_adj_2346), 
            .I3(n17153), .O(n17238));   // coms.v(235[16:291])
    defparam i8_4_lut_adj_617.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_618 (.I0(n1034), .I1(n10139), .I2(n9378), 
            .I3(GND_net), .O(n47_adj_2347));
    defparam i1_2_lut_3_lut_adj_618.LUT_INIT = 16'h1010;
    SB_LUT4 i14692_4_lut (.I0(\data_out_frame2[0] [7]), .I1(n26_adj_2174), 
            .I2(n5817), .I3(n12491), .O(n17469));
    defparam i14692_4_lut.LUT_INIT = 16'hfa8a;
    SB_LUT4 select_219_Select_23_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [23]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2244));   // coms.v(430[13] 433[7])
    defparam select_219_Select_23_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15326 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [6]), .I2(\data_out_frame2[15] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n18118));
    defparam byte_transmit_counter2_0__bdd_4_lut_15326.LUT_INIT = 16'he4aa;
    SB_LUT4 select_219_Select_22_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [22]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2246));   // coms.v(430[13] 433[7])
    defparam select_219_Select_22_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i15059_3_lut_4_lut (.I0(\data_out_frame2[0] [4]), .I1(n12491), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n488), .O(n17686));
    defparam i15059_3_lut_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 n18118_bdd_4_lut (.I0(n18118), .I1(\data_out_frame2[13] [6]), 
            .I2(\data_out_frame2[12] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n18121));
    defparam n18118_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \data_in_3[[3__2266  (.Q(\data_in[3] [3]), .C(CLK_c), .D(n11119));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_3[[2__2267  (.Q(\data_in[3] [2]), .C(CLK_c), .D(n11118));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(n5_adj_8), 
            .I2(n17086), .I3(n9), .O(n10009));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'hf2f7;
    SB_LUT4 i15063_3_lut_4_lut (.I0(\data_out_frame2[0] [3]), .I1(n12491), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n488), .O(n17688));
    defparam i15063_3_lut_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i14694_4_lut (.I0(n17469), .I1(n4494), .I2(n5815), .I3(n5817), 
            .O(n17471));
    defparam i14694_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_219_Select_3_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [3]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2284));
    defparam select_219_Select_3_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut (.I0(n63), .I1(n4408), .I2(n63_adj_9), .I3(n63_adj_10), 
            .O(n9369));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i14695_4_lut (.I0(\data_out_frame2[0] [6]), .I1(n26_adj_2174), 
            .I2(n5817), .I3(n12491), .O(n17472));
    defparam i14695_4_lut.LUT_INIT = 16'hfa8a;
    SB_LUT4 i14697_4_lut (.I0(n17472), .I1(n4494), .I2(n5815), .I3(n5817), 
            .O(n17474));
    defparam i14697_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_219_Select_17_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [17]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2257));   // coms.v(430[13] 433[7])
    defparam select_219_Select_17_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_21_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [21]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2248));   // coms.v(430[13] 433[7])
    defparam select_219_Select_21_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_4_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [4]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2283));
    defparam select_219_Select_4_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15186_2_lut_3_lut (.I0(n16267), .I1(tx_active), .I2(r_SM_Main_2__N_2034[0]), 
            .I3(GND_net), .O(n445));   // coms.v(305[16] 313[10])
    defparam i15186_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i1_3_lut (.I0(\data_out[0] [6]), 
            .I1(\data_out[1][6] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n1_adj_2160));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15119_2_lut (.I0(\data_out[3] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17612));
    defparam i15119_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14698_4_lut (.I0(\data_out_frame2[0] [5]), .I1(n26_adj_2174), 
            .I2(n5817), .I3(n12491), .O(n17475));
    defparam i14698_4_lut.LUT_INIT = 16'hfa8a;
    SB_DFF \data_in_3[[1__2268  (.Q(\data_in[3] [1]), .C(CLK_c), .D(n11117));   // coms.v(416[12] 543[6])
    SB_LUT4 i14700_4_lut (.I0(n17475), .I1(n4494), .I2(n5815), .I3(n5817), 
            .O(n17477));
    defparam i14700_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_219_Select_20_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [20]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2250));   // coms.v(430[13] 433[7])
    defparam select_219_Select_20_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_5_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [5]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2281));
    defparam select_219_Select_5_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1026_2_lut_3_lut_4_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(n17206), .I3(\data_in_frame[0] [0]), .O(n2138));   // coms.v(76[16:69])
    defparam i1026_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i2 (.Q(\data_out_frame2[0] [1]), .C(CLK_c), 
           .D(n17489));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_3[[0__2269  (.Q(\data_in[3] [0]), .C(CLK_c), .D(n11116));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_2[[7__2270  (.Q(\data_in[2] [7]), .C(CLK_c), .D(n11115));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i8_3_lut (.I0(\data_out[8][5] ), 
            .I1(\data_out[9] [5]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2352));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame2[6] [5]), 
            .I1(\data_out_frame2[7] [5]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2353));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i10_4_lut (.I0(n8_adj_2352), 
            .I1(\data_out[10] [5]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_11));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_619 (.I0(n1034), .I1(n3_c), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_2279));   // coms.v(373[7:20])
    defparam i1_2_lut_adj_619.LUT_INIT = 16'h8888;
    SB_DFF \data_in_2[[6__2271  (.Q(\data_in[2] [6]), .C(CLK_c), .D(n11114));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out[6] [6]), 
            .I1(\data_out[7] [6]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2159));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n10018), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state[1] ), 
            .O(\FRAME_MATCHER.i_31__N_1272 ));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 select_219_Select_7_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [7]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2277));
    defparam select_219_Select_7_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_620 (.I0(\FRAME_MATCHER.state[2] ), .I1(n10018), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state[1] ), 
            .O(\FRAME_MATCHER.i_31__N_1273 ));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_3_lut_4_lut_adj_620.LUT_INIT = 16'h0020;
    SB_LUT4 i15149_2_lut (.I0(data_out_7__2__N_447), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17698));
    defparam i15149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_219_Select_19_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [19]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2252));   // coms.v(430[13] 433[7])
    defparam select_219_Select_19_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_18_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [18]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2254));   // coms.v(430[13] 433[7])
    defparam select_219_Select_18_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_13_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [13]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2266));   // coms.v(430[13] 433[7])
    defparam select_219_Select_13_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut (.I0(\data_out_frame2[5] [5]), 
            .I1(n5_adj_2353), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_c));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 select_219_Select_12_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [12]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2268));   // coms.v(430[13] 433[7])
    defparam select_219_Select_12_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF \data_in_2[[5__2272  (.Q(\data_in[2] [5]), .C(CLK_c), .D(n11113));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_3_lut_adj_621 (.I0(\data_out_frame2[8] [3]), .I1(\data_out_frame2[6] [4]), 
            .I2(\data_out_frame2[7] [6]), .I3(GND_net), .O(n6_adj_2339));   // coms.v(239[17:230])
    defparam i1_2_lut_3_lut_adj_621.LUT_INIT = 16'h9696;
    SB_DFF \data_in_2[[4__2273  (.Q(\data_in[2] [4]), .C(CLK_c), .D(n11111));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_8_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [8]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2275));
    defparam select_219_Select_8_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15103_2_lut (.I0(\data_out[1] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17675));
    defparam i15103_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF \data_in_2[[3__2274  (.Q(\data_in[2] [3]), .C(CLK_c), .D(n11110));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_2[[2__2275  (.Q(\data_in[2] [2]), .C(CLK_c), .D(n11109));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_11_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [11]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2270));   // coms.v(430[13] 433[7])
    defparam select_219_Select_11_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_3_lut_adj_622 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n17102));   // coms.v(505[9:81])
    defparam i1_3_lut_adj_622.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_623 (.I0(\data_in_frame[1] [6]), .I1(n10407), .I2(\data_in_frame[5] [7]), 
            .I3(n17213), .O(n17214));   // coms.v(130[17:124])
    defparam i3_4_lut_adj_623.LUT_INIT = 16'h6996;
    SB_LUT4 select_219_Select_9_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [9]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2273));
    defparam select_219_Select_9_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15208_4_lut_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(n10596));
    defparam i15208_4_lut_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 select_219_Select_10_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [10]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2271));
    defparam select_219_Select_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10566_2_lut (.I0(\UART_TRANSMITTER.state[0] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n2593[0]));   // coms.v(283[4] 369[11])
    defparam i10566_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_624 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[6] [2]), .O(n16353));
    defparam i2_3_lut_4_lut_adj_624.LUT_INIT = 16'h6996;
    SB_LUT4 select_219_Select_11_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [11]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2269));
    defparam select_219_Select_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4980_2_lut (.I0(n63_adj_9), .I1(n63_adj_10), .I2(GND_net), 
            .I3(GND_net), .O(n10088));   // coms.v(427[13] 433[7])
    defparam i4980_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15100_2_lut (.I0(\data_out[3][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17676));
    defparam i15100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out[6] [4]), 
            .I1(\data_out[7] [4]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2136));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15173_2_lut (.I0(\data_out[5] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17764));
    defparam i15173_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \data_in_2[[1__2276  (.Q(\data_in[2] [1]), .C(CLK_c), .D(n11108));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_2[[0__2277  (.Q(\data_in[2] [0]), .C(CLK_c), .D(n11107));   // coms.v(416[12] 543[6])
    SB_LUT4 i10579_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n9995), .I2(\FRAME_MATCHER.i [31]), 
            .I3(GND_net), .O(n4408));   // coms.v(523[9:58])
    defparam i10579_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 select_219_Select_12_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [12]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2267));
    defparam select_219_Select_12_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14556_2_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n17331));
    defparam i14556_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10589_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n10161), .I3(\FRAME_MATCHER.i [0]), .O(n2061));   // coms.v(443[9:60])
    defparam i10589_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i5_4_lut_adj_625 (.I0(\data_in[2] [4]), .I1(\data_in[3] [3]), 
            .I2(\data_in[2] [6]), .I3(\data_in[2] [1]), .O(n12_adj_2355));   // coms.v(430[16:93])
    defparam i5_4_lut_adj_625.LUT_INIT = 16'hfffe;
    SB_LUT4 i14633_4_lut (.I0(\data_in[1] [5]), .I1(\data_in[0] [4]), .I2(\data_in[1] [0]), 
            .I3(n17331), .O(n17410));
    defparam i14633_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_adj_626 (.I0(\FRAME_MATCHER.state[1] ), .I1(n5_adj_8), 
            .I2(n17086), .I3(GND_net), .O(n1034));
    defparam i1_2_lut_3_lut_adj_626.LUT_INIT = 16'hf2f2;
    SB_LUT4 i6_4_lut_adj_627 (.I0(n17410), .I1(n12_adj_2355), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n10133));   // coms.v(430[16:93])
    defparam i6_4_lut_adj_627.LUT_INIT = 16'hfffd;
    SB_DFF \data_in_1[[7__2278  (.Q(\data_in[1] [7]), .C(CLK_c), .D(n11106));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_13_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [13]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2265));
    defparam select_219_Select_13_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_628 (.I0(\data_in[1] [2]), .I1(\data_in[1] [1]), 
            .I2(\data_in[3] [6]), .I3(GND_net), .O(n10141));   // coms.v(427[16:89])
    defparam i2_3_lut_adj_628.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_adj_629 (.I0(\FRAME_MATCHER.state[1] ), .I1(n5_adj_8), 
            .I2(GND_net), .I3(GND_net), .O(n44));
    defparam i1_2_lut_adj_629.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_630 (.I0(\FRAME_MATCHER.i_31__N_1273 ), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n5_adj_8), .I3(GND_net), .O(n17086));
    defparam i1_2_lut_3_lut_adj_630.LUT_INIT = 16'habab;
    SB_LUT4 i1_2_lut_adj_631 (.I0(\data_in[0] [6]), .I1(n10133), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_2356));
    defparam i1_2_lut_adj_631.LUT_INIT = 16'heeee;
    SB_LUT4 i14629_4_lut (.I0(\data_in[3] [0]), .I1(\data_in[3] [4]), .I2(\data_in[3] [2]), 
            .I3(\data_in[0] [5]), .O(n17406));
    defparam i14629_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15230_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(n10594));
    defparam i15230_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_DFF \data_in_1[[6__2279  (.Q(\data_in[1] [6]), .C(CLK_c), .D(n11105));   // coms.v(416[12] 543[6])
    SB_LUT4 i4_4_lut_adj_632 (.I0(\data_in[1] [4]), .I1(n17406), .I2(\data_in[2] [3]), 
            .I3(n6_adj_2356), .O(n10027));
    defparam i4_4_lut_adj_632.LUT_INIT = 16'hfffb;
    SB_LUT4 i5_4_lut_adj_633 (.I0(\data_in_frame[5] [4]), .I1(n17102), .I2(\data_in_frame[1] [3]), 
            .I3(\data_in_frame[1] [2]), .O(n21_adj_2357));
    defparam i5_4_lut_adj_633.LUT_INIT = 16'hedde;
    SB_LUT4 select_219_Select_14_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [14]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2263));
    defparam select_219_Select_14_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14623_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[2] [5]), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n17400));
    defparam i14623_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_adj_634 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[5] [5]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n16474));   // coms.v(505[9:81])
    defparam i2_3_lut_adj_634.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_635 (.I0(\data_in[3] [7]), .I1(\data_in[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2358));   // coms.v(430[16:93])
    defparam i1_2_lut_adj_635.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_636 (.I0(\FRAME_MATCHER.state[2] ), .I1(n10018), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n5_adj_8));
    defparam i1_2_lut_3_lut_adj_636.LUT_INIT = 16'hefef;
    SB_LUT4 i3_4_lut_adj_637 (.I0(\data_in[2] [2]), .I1(n6_adj_2358), .I2(n17400), 
            .I3(\data_in[2] [0]), .O(n8_adj_2359));   // coms.v(430[16:93])
    defparam i3_4_lut_adj_637.LUT_INIT = 16'hdfff;
    SB_LUT4 i1_2_lut_3_lut_adj_638 (.I0(n63), .I1(n63_adj_9), .I2(n63_adj_10), 
            .I3(GND_net), .O(n9378));
    defparam i1_2_lut_3_lut_adj_638.LUT_INIT = 16'h8080;
    SB_LUT4 select_219_Select_15_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [15]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2260));
    defparam select_219_Select_15_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_639 (.I0(\FRAME_MATCHER.i [2]), .I1(n9995), .I2(GND_net), 
            .I3(GND_net), .O(n10161));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_639.LUT_INIT = 16'heeee;
    SB_LUT4 i10774_2_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n13450));
    defparam i10774_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_640 (.I0(\data_in[1] [6]), .I1(n13450), .I2(n8_adj_2359), 
            .I3(\data_in[3] [5]), .O(n10136));   // coms.v(430[16:93])
    defparam i1_4_lut_adj_640.LUT_INIT = 16'hfffb;
    SB_LUT4 i14611_2_lut (.I0(\data_in[1] [2]), .I1(\data_in[3] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n17388));
    defparam i14611_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_641 (.I0(\FRAME_MATCHER.state[1] ), .I1(n5_adj_8), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1275 ));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_641.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_642 (.I0(n10136), .I1(n10027), .I2(\data_in[1] [1]), 
            .I3(n17388), .O(n63));
    defparam i3_4_lut_adj_642.LUT_INIT = 16'hfeff;
    SB_LUT4 select_219_Select_10_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [10]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2272));   // coms.v(430[13] 433[7])
    defparam select_219_Select_10_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i15212_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(data_out_10__7__N_110));
    defparam i15212_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2_4_lut_adj_643 (.I0(n17114), .I1(\data_in_frame[1] [0]), .I2(\data_in_frame[5] [1]), 
            .I3(\data_in_frame[0] [7]), .O(n18_adj_2360));
    defparam i2_4_lut_adj_643.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_2_lut_adj_644 (.I0(n1034), .I1(n10139), .I2(GND_net), .I3(GND_net), 
            .O(n10140));
    defparam i1_2_lut_adj_644.LUT_INIT = 16'heeee;
    SB_LUT4 i14710_4_lut (.I0(\data_out_frame2[0] [1]), .I1(n26_adj_2174), 
            .I2(n5817), .I3(n12491), .O(n17487));
    defparam i14710_4_lut.LUT_INIT = 16'hfa8a;
    SB_LUT4 i6_4_lut_adj_645 (.I0(n10136), .I1(\data_in[1] [4]), .I2(\data_in[3] [0]), 
            .I3(\data_in[3] [2]), .O(n16_adj_2361));
    defparam i6_4_lut_adj_645.LUT_INIT = 16'hfffb;
    SB_LUT4 i7_4_lut_adj_646 (.I0(\data_in[3] [4]), .I1(\data_in[0] [5]), 
            .I2(\data_in[0] [6]), .I3(n10133), .O(n17_adj_2362));
    defparam i7_4_lut_adj_646.LUT_INIT = 16'hffef;
    SB_LUT4 i9_4_lut_adj_647 (.I0(n17_adj_2362), .I1(n10141), .I2(n16_adj_2361), 
            .I3(\data_in[2] [3]), .O(n63_adj_10));
    defparam i9_4_lut_adj_647.LUT_INIT = 16'hfeff;
    SB_LUT4 i14625_4_lut (.I0(\data_in[3] [5]), .I1(\data_in[1] [6]), .I2(\data_in[3] [7]), 
            .I3(\data_in[0] [0]), .O(n17402));
    defparam i14625_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i14712_4_lut (.I0(n17487), .I1(n4494), .I2(n5815), .I3(n5817), 
            .O(n17489));
    defparam i14712_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF \data_in_1[[5__2280  (.Q(\data_in[1] [5]), .C(CLK_c), .D(n11104));   // coms.v(416[12] 543[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame2[11] [2]), .I1(n10359), 
            .I2(n10434), .I3(n17237), .O(n14_adj_2346));   // coms.v(235[16:291])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF \data_in_1[[4__2281  (.Q(\data_in[1] [4]), .C(CLK_c), .D(n11103));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_3_lut_adj_648 (.I0(\data_out_frame2[11] [2]), .I1(n10359), 
            .I2(\data_out_frame2[11] [1]), .I3(GND_net), .O(n17174));   // coms.v(235[16:291])
    defparam i1_2_lut_3_lut_adj_648.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut (.I0(n18133), .I1(\data_out_frame2[20] [7]), 
            .I2(byte_transmit_counter2[2]), .I3(n9157), .O(n22_adj_2363));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i31_4_lut (.I0(n18217), .I1(n22_adj_2363), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[7]));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_219_Select_16_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [16]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2258));
    defparam select_219_Select_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15061_3_lut_4_lut (.I0(\data_out_frame2[0] [2]), .I1(n12491), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n488), .O(n17690));
    defparam i15061_3_lut_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut (.I0(n18115), .I1(\data_out_frame2[20] [6]), 
            .I2(byte_transmit_counter2[2]), .I3(n9157), .O(n22_adj_2364));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF \data_in_1[[3__2282  (.Q(\data_in[1] [3]), .C(CLK_c), .D(n11102));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_1[[2__2283  (.Q(\data_in[1] [2]), .C(CLK_c), .D(n11101));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i31_4_lut (.I0(n18181), .I1(n22_adj_2364), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[6]));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_219_Select_9_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [9]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2274));   // coms.v(430[13] 433[7])
    defparam select_219_Select_9_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_17_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [17]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2256));
    defparam select_219_Select_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10953_1_lut (.I0(n13628), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(tx2_transmit_N_1996));
    defparam i10953_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 select_219_Select_8_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [8]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2276));   // coms.v(430[13] 433[7])
    defparam select_219_Select_8_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF \data_in_1[[1__2284  (.Q(\data_in[1] [1]), .C(CLK_c), .D(n11100));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut (.I0(n18097), .I1(\data_out_frame2[20] [5]), 
            .I2(byte_transmit_counter2[2]), .I3(n9157), .O(n22_adj_2365));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i6_4_lut_adj_649 (.I0(\data_in[2] [7]), .I1(n10141), .I2(\data_in[2] [2]), 
            .I3(n10027), .O(n16_adj_2366));   // coms.v(427[16:89])
    defparam i6_4_lut_adj_649.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_650 (.I0(\data_out_frame2[8] [3]), .I1(\data_out_frame2[6] [4]), 
            .I2(\data_out_frame2[10] [0]), .I3(\data_out_frame2[10] [2]), 
            .O(n17228));   // coms.v(239[17:230])
    defparam i1_2_lut_3_lut_4_lut_adj_650.LUT_INIT = 16'h6996;
    SB_DFF \data_in_1[[0__2285  (.Q(\data_in[1] [0]), .C(CLK_c), .D(n11099));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_0[[7__2286  (.Q(\data_in[0] [7]), .C(CLK_c), .D(n11098));   // coms.v(416[12] 543[6])
    SB_LUT4 i10670_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [18]));   // coms.v(430[13] 433[7])
    defparam i10670_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \data_in_0[[6__2287  (.Q(\data_in[0] [6]), .C(CLK_c), .D(n11097));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_7_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [7]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2278));   // coms.v(430[13] 433[7])
    defparam select_219_Select_7_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i2_3_lut_4_lut_adj_651 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[6] [3]), .O(n16352));
    defparam i2_3_lut_4_lut_adj_651.LUT_INIT = 16'h6996;
    SB_DFF \data_in_0[[5__2288  (.Q(\data_in[0] [5]), .C(CLK_c), .D(n11096));   // coms.v(416[12] 543[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i31_4_lut (.I0(n18265), .I1(n22_adj_2365), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[5]));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF \data_in_0[[4__2289  (.Q(\data_in[0] [4]), .C(CLK_c), .D(n11095));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_3_lut_adj_652 (.I0(n13146), .I1(\FRAME_MATCHER.i [6]), 
            .I2(n10009), .I3(GND_net), .O(n3_adj_2280));
    defparam i1_2_lut_3_lut_adj_652.LUT_INIT = 16'h0808;
    SB_LUT4 i2_3_lut_4_lut_adj_653 (.I0(\data_out_frame2[12] [1]), .I1(\data_out_frame2[12] [3]), 
            .I2(n10413), .I3(\data_out_frame2[10] [4]), .O(n17282));   // coms.v(239[17:230])
    defparam i2_3_lut_4_lut_adj_653.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut (.I0(n18277), .I1(\data_out_frame2[20] [4]), 
            .I2(byte_transmit_counter2[2]), .I3(n9157), .O(n22_adj_2367));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_219_Select_18_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [18]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2253));
    defparam select_219_Select_18_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10_4_lut_adj_654 (.I0(n19_adj_2324), .I1(n16475), .I2(n2120), 
            .I3(\data_in_frame[6] [4]), .O(n26_adj_2368));
    defparam i10_4_lut_adj_654.LUT_INIT = 16'heffe;
    SB_LUT4 i10669_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [19]));   // coms.v(430[13] 433[7])
    defparam i10669_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \data_in_0[[3__2290  (.Q(\data_in[0] [3]), .C(CLK_c), .D(n11094));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_0[[2__2291  (.Q(\data_in[0] [2]), .C(CLK_c), .D(n11093));   // coms.v(416[12] 543[6])
    SB_DFF \data_in_0[[1__2292  (.Q(\data_in[0] [1]), .C(CLK_c), .D(n11092));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_3_lut_adj_655 (.I0(\data_out_frame2[12] [1]), .I1(\data_out_frame2[12] [3]), 
            .I2(\data_out_frame2[10] [3]), .I3(GND_net), .O(n17249));   // coms.v(239[17:230])
    defparam i1_2_lut_3_lut_adj_655.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i31_4_lut (.I0(n18037), .I1(n22_adj_2367), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[4]));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF \data_in_0[[0__2293  (.Q(\data_in[0] [0]), .C(CLK_c), .D(n11091));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(n31), .I1(n9), .I2(\FRAME_MATCHER.state[1] ), 
            .I3(GND_net), .O(n1_adj_12));   // coms.v(449[9:87])
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i3_4_lut_4_lut (.I0(n31), .I1(n51_adj_2173), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(\FRAME_MATCHER.state[2] ), .O(n10725));   // coms.v(449[9:87])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i2_3_lut_adj_656 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n15164));   // coms.v(416[12] 543[6])
    defparam i2_3_lut_adj_656.LUT_INIT = 16'hfefe;
    SB_LUT4 select_219_Select_19_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [19]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2251));
    defparam select_219_Select_19_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_657 (.I0(\data_in[2] [5]), .I1(\data_in[2] [0]), 
            .I2(\data_in[0] [1]), .I3(\data_in[0] [3]), .O(n17_adj_2370));   // coms.v(427[16:89])
    defparam i7_4_lut_adj_657.LUT_INIT = 16'hfffe;
    SB_DFF \UART_TRANSMITTER.state__i2  (.Q(\UART_TRANSMITTER.state[1] ), 
           .C(CLK_c), .D(n16618));   // coms.v(280[12] 370[6])
    SB_LUT4 i1_2_lut_adj_658 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i1_2_lut_adj_658.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut (.I0(n18055), .I1(\data_out_frame2[20] [3]), 
            .I2(byte_transmit_counter2[2]), .I3(n9157), .O(n22_adj_2371));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i31_4_lut (.I0(n18259), .I1(n22_adj_2371), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[3]));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n5817_bdd_4_lut_15430_4_lut (.I0(n31), .I1(n5815), .I2(n4494), 
            .I3(n5817), .O(n18202));   // coms.v(449[9:87])
    defparam n5817_bdd_4_lut_15430_4_lut.LUT_INIT = 16'h77c0;
    SB_LUT4 i8223_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10596), .I3(\data_out[1] [2]), .O(n10909));   // coms.v(283[4] 369[11])
    defparam i8223_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut (.I0(n18031), .I1(\data_out_frame2[20] [2]), 
            .I2(byte_transmit_counter2[2]), .I3(n9157), .O(n22_adj_2372));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_659 (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_2373));   // coms.v(440[7:23])
    defparam i1_2_lut_adj_659.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_660 (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [20]), .I3(\FRAME_MATCHER.i [23]), .O(n42));   // coms.v(440[7:23])
    defparam i17_4_lut_adj_660.LUT_INIT = 16'hfffe;
    SB_LUT4 i10668_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [20]));   // coms.v(430[13] 433[7])
    defparam i10668_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8210_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10596), .I3(\data_out[3] [6]), .O(n10896));   // coms.v(283[4] 369[11])
    defparam i8210_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i31_4_lut (.I0(n18247), .I1(n22_adj_2372), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[2]));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15_4_lut_adj_661 (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(\FRAME_MATCHER.i [25]), .I3(\FRAME_MATCHER.i [30]), .O(n40));   // coms.v(440[7:23])
    defparam i15_4_lut_adj_661.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_662 (.I0(n16352), .I1(n24_adj_2340), .I2(n2122), 
            .I3(\data_in_frame[6] [5]), .O(n28_adj_2374));
    defparam i12_4_lut_adj_662.LUT_INIT = 16'hdffd;
    SB_LUT4 i1_2_lut_3_lut_adj_663 (.I0(n13146), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n10009), .I3(GND_net), .O(n3_adj_2282));
    defparam i1_2_lut_3_lut_adj_663.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_20_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [20]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2249));
    defparam select_219_Select_20_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_664 (.I0(\data_out_frame2[15] [2]), .I1(\data_out_frame2[16] [2]), 
            .I2(\data_out_frame2[15] [3]), .I3(GND_net), .O(n17291));   // coms.v(228[16:596])
    defparam i1_2_lut_3_lut_adj_664.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut (.I0(n18013), .I1(\data_out_frame2[20] [1]), 
            .I2(byte_transmit_counter2[2]), .I3(n9157), .O(n22_adj_2375));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i31_4_lut (.I0(n18241), .I1(n22_adj_2375), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[1]));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i2_3_lut_4_lut_adj_665 (.I0(\data_out_frame2[15] [2]), .I1(\data_out_frame2[16] [2]), 
            .I2(\data_out_frame2[5] [0]), .I3(\data_out_frame2[8] [2]), 
            .O(n10507));   // coms.v(228[16:596])
    defparam i2_3_lut_4_lut_adj_665.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_666 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [14]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [16]), .O(n41_adj_2376));   // coms.v(440[7:23])
    defparam i16_4_lut_adj_666.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_667 (.I0(\data_out_frame2[5] [1]), .I1(\data_out_frame2[12] [4]), 
            .I2(\data_out_frame2[12] [5]), .I3(\data_out_frame2[10] [6]), 
            .O(n17135));   // coms.v(239[17:230])
    defparam i2_3_lut_4_lut_adj_667.LUT_INIT = 16'h6996;
    SB_LUT4 i10667_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [21]));   // coms.v(430[13] 433[7])
    defparam i10667_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14_4_lut_adj_668 (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [27]), .I3(\FRAME_MATCHER.i [22]), .O(n39_adj_2377));   // coms.v(440[7:23])
    defparam i14_4_lut_adj_668.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_669 (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n26_adj_2373), .O(n44_adj_2378));   // coms.v(440[7:23])
    defparam i19_4_lut_adj_669.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_670 (.I0(n17_adj_2370), .I1(\data_in[1] [7]), .I2(n16_adj_2366), 
            .I3(n17402), .O(n63_adj_9));   // coms.v(427[16:89])
    defparam i9_4_lut_adj_670.LUT_INIT = 16'hfeff;
    SB_LUT4 i23_4_lut (.I0(n39_adj_2377), .I1(n41_adj_2376), .I2(n40), 
            .I3(n42), .O(n48_adj_2379));   // coms.v(440[7:23])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \UART_TRANSMITTER.state__i3  (.Q(\UART_TRANSMITTER.state[2] ), 
           .C(CLK_c), .D(n13));   // coms.v(280[12] 370[6])
    SB_LUT4 i5_3_lut_4_lut_adj_671 (.I0(\data_out_frame2[5] [1]), .I1(\data_out_frame2[12] [4]), 
            .I2(\data_out_frame2[12] [0]), .I3(n17288), .O(n14_adj_2292));   // coms.v(239[17:230])
    defparam i5_3_lut_4_lut_adj_671.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i3 (.Q(\data_out_frame2[0] [2]), .C(CLK_c), 
           .D(n18193));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_4_lut_adj_672 (.I0(\data_out_frame2[11] [3]), .I1(\data_out_frame2[11] [4]), 
            .I2(\data_out_frame2[11] [6]), .I3(\data_out_frame2[11] [5]), 
            .O(n10359));   // coms.v(237[17:221])
    defparam i1_2_lut_4_lut_adj_672.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_673 (.I0(n63_adj_9), .I1(n63_adj_10), .I2(n63), 
            .I3(GND_net), .O(n13146));   // coms.v(443[6] 445[9])
    defparam i2_3_lut_adj_673.LUT_INIT = 16'h8080;
    SB_LUT4 i18_4_lut_adj_674 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [7]), .I3(\FRAME_MATCHER.i [13]), .O(n43_adj_2380));   // coms.v(440[7:23])
    defparam i18_4_lut_adj_674.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_675 (.I0(n43_adj_2380), .I1(n15164), .I2(n48_adj_2379), 
            .I3(n44_adj_2378), .O(n9995));   // coms.v(440[7:23])
    defparam i1_4_lut_adj_675.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_676 (.I0(n21_adj_2357), .I1(n17214), .I2(n2124), 
            .I3(\data_in_frame[6] [6]), .O(n27_adj_2381));
    defparam i11_4_lut_adj_676.LUT_INIT = 16'hbffb;
    SB_LUT4 i1_3_lut_4_lut_adj_677 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n10018), .I3(\FRAME_MATCHER.state[2] ), .O(n5817));   // coms.v(409[11:16])
    defparam i1_3_lut_4_lut_adj_677.LUT_INIT = 16'h0c04;
    SB_LUT4 select_219_Select_16_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [16]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2259));   // coms.v(430[13] 433[7])
    defparam select_219_Select_16_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_219_Select_21_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [21]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2247));
    defparam select_219_Select_21_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10671_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [17]));   // coms.v(430[13] 433[7])
    defparam i10671_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_678 (.I0(n16353), .I1(n26_adj_2368), .I2(n18_adj_2360), 
            .I3(n16474), .O(n29));
    defparam i13_4_lut_adj_678.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_679 (.I0(byte_transmit_counter2[7]), .I1(n11833), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2345));   // coms.v(409[11:16])
    defparam i1_2_lut_adj_679.LUT_INIT = 16'h8888;
    SB_LUT4 select_224_Select_7_i2_4_lut (.I0(byte_transmit_counter2[7]), 
            .I1(\FRAME_MATCHER.i_31__N_1272 ), .I2(n17714), .I3(n11867), 
            .O(n2_adj_2344));
    defparam select_224_Select_7_i2_4_lut.LUT_INIT = 16'h88c0;
    SB_LUT4 i15075_2_lut (.I0(\data_out[0][3] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17696));
    defparam i15075_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10584_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n9995), .I3(n39), .O(n3779));   // coms.v(499[9:54])
    defparam i10584_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_3_lut_adj_680 (.I0(\data_out_frame2[11] [4]), .I1(\data_out_frame2[11] [6]), 
            .I2(\data_out_frame2[11] [5]), .I3(GND_net), .O(n17203));   // coms.v(237[17:221])
    defparam i1_2_lut_3_lut_adj_680.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame2_0___i4 (.Q(\data_out_frame2[0] [3]), .C(CLK_c), 
           .D(n18205));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i5 (.Q(\data_out_frame2[0] [4]), .C(CLK_c), 
           .D(n18253));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i6 (.Q(\data_out_frame2[0] [5]), .C(CLK_c), 
           .D(n17477));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i7 (.Q(\data_out_frame2[0] [6]), .C(CLK_c), 
           .D(n17474));   // coms.v(416[12] 543[6])
    SB_DFF data_out_frame2_0___i8 (.Q(\data_out_frame2[0] [7]), .C(CLK_c), 
           .D(n17471));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i153 (.Q(\data_out_frame2[19] [0]), .C(CLK_c), 
            .E(n10725), .D(n17238));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i154 (.Q(\data_out_frame2[19] [1]), .C(CLK_c), 
            .E(n10725), .D(n17274));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i155 (.Q(\data_out_frame2[19] [2]), .C(CLK_c), 
            .E(n10725), .D(n17284));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i156 (.Q(\data_out_frame2[19] [3]), .C(CLK_c), 
            .E(n10725), .D(n17250));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i157 (.Q(\data_out_frame2[19] [4]), .C(CLK_c), 
            .E(n10725), .D(n17313));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i158 (.Q(\data_out_frame2[19] [5]), .C(CLK_c), 
            .E(n10725), .D(n17290));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i159 (.Q(\data_out_frame2[19] [6]), .C(CLK_c), 
            .E(n10725), .D(n17310));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i160 (.Q(\data_out_frame2[19] [7]), .C(CLK_c), 
            .E(n10725), .D(n17301));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i161 (.Q(\data_out_frame2[20] [0]), .C(CLK_c), 
            .E(n10725), .D(n17275));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i162 (.Q(\data_out_frame2[20] [1]), .C(CLK_c), 
            .E(n10725), .D(n17281));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i163 (.Q(\data_out_frame2[20] [2]), .C(CLK_c), 
            .E(n10725), .D(n17296));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i164 (.Q(\data_out_frame2[20] [3]), .C(CLK_c), 
            .E(n10725), .D(n17295));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i165 (.Q(\data_out_frame2[20] [4]), .C(CLK_c), 
            .E(n10725), .D(n17308));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i166 (.Q(\data_out_frame2[20] [5]), .C(CLK_c), 
            .E(n10725), .D(n17307));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i167 (.Q(\data_out_frame2[20] [6]), .C(CLK_c), 
            .E(n10725), .D(n17304));   // coms.v(416[12] 543[6])
    SB_DFFE data_out_frame2_0___i168 (.Q(\data_out_frame2[20] [7]), .C(CLK_c), 
            .E(n10725), .D(n17302));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n11076));   // coms.v(416[12] 543[6])
    SB_LUT4 i10666_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [22]));   // coms.v(430[13] 433[7])
    defparam i10666_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_681 (.I0(\data_out_frame2[12] [2]), .I1(\data_out_frame2[8] [4]), 
            .I2(\data_out_frame2[8] [0]), .I3(GND_net), .O(n17098));   // coms.v(227[16:31])
    defparam i1_2_lut_3_lut_adj_681.LUT_INIT = 16'h9696;
    SB_LUT4 i9895_3_lut (.I0(\data_out[8]_c [0]), .I1(\rand_setpoint[0] ), 
            .I2(data_out_10__7__N_110), .I3(GND_net), .O(n11122));   // coms.v(21[11:19])
    defparam i9895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_219_Select_22_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [22]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2245));
    defparam select_219_Select_22_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_219_Select_15_i3_2_lut_3_lut (.I0(\FRAME_MATCHER.i [15]), 
            .I1(n13146), .I2(n10009), .I3(GND_net), .O(n3_adj_2261));   // coms.v(430[13] 433[7])
    defparam select_219_Select_15_i3_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i10665_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [23]));   // coms.v(430[13] 433[7])
    defparam i10665_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_682 (.I0(\data_out_frame2[10] [1]), .I1(\data_out_frame2[12] [0]), 
            .I2(\data_out_frame2[11] [7]), .I3(GND_net), .O(n17194));   // coms.v(238[17:230])
    defparam i1_2_lut_3_lut_adj_682.LUT_INIT = 16'h9696;
    SB_LUT4 select_219_Select_23_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [23]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2243));
    defparam select_219_Select_23_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10664_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [24]));   // coms.v(430[13] 433[7])
    defparam i10664_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_683 (.I0(\data_out_frame2[9] [5]), .I1(\data_out_frame2[6] [1]), 
            .I2(\data_out_frame2[7] [7]), .I3(\data_out_frame2[9] [7]), 
            .O(n10349));   // coms.v(234[16:291])
    defparam i2_3_lut_4_lut_adj_683.LUT_INIT = 16'h6996;
    SB_LUT4 select_219_Select_24_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [24]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2241));
    defparam select_219_Select_24_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10663_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [25]));   // coms.v(430[13] 433[7])
    defparam i10663_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_684 (.I0(\data_out_frame2[16] [6]), .I1(\data_out_frame2[15] [0]), 
            .I2(\data_out_frame2[16] [0]), .I3(\data_out_frame2[13] [2]), 
            .O(n17267));   // coms.v(237[17:221])
    defparam i1_2_lut_4_lut_adj_684.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_685 (.I0(\data_out_frame2[9] [6]), .I1(\data_out_frame2[8] [1]), 
            .I2(\data_out_frame2[6] [2]), .I3(GND_net), .O(n10371));   // coms.v(237[17:221])
    defparam i1_2_lut_3_lut_adj_685.LUT_INIT = 16'h9696;
    SB_LUT4 select_219_Select_25_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [25]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2239));
    defparam select_219_Select_25_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10662_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [26]));   // coms.v(430[13] 433[7])
    defparam i10662_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14597_3_lut_4_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[2] [0]), .O(n17373));
    defparam i14597_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 select_219_Select_26_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [26]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2237));
    defparam select_219_Select_26_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_686 (.I0(n13146), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [27]));
    defparam i1_2_lut_adj_686.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_687 (.I0(tx2_active), .I1(r_SM_Main_2__N_2034_adj_2405[0]), 
            .I2(n13628), .I3(GND_net), .O(n488));
    defparam i1_2_lut_3_lut_adj_687.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_4_lut_adj_688 (.I0(\data_out[8][3] ), .I1(\data_out[8][2] ), 
            .I2(\data_out[10] [4]), .I3(\data_out[10][0] ), .O(n17222));   // coms.v(176[16:77])
    defparam i2_3_lut_4_lut_adj_688.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n11075));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n11074));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n11073));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n11072));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n11071));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_27_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [27]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2235));
    defparam select_219_Select_27_i2_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n11070));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n11069));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n11068));   // coms.v(416[12] 543[6])
    SB_LUT4 i15101_2_lut (.I0(\data_out[2] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17697));
    defparam i15101_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n11067));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_3_lut_adj_689 (.I0(\data_out[8][3] ), .I1(\data_out[8][2] ), 
            .I2(\data_out[8][1] ), .I3(GND_net), .O(n10188));   // coms.v(176[16:77])
    defparam i1_2_lut_3_lut_adj_689.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n11066));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n11065));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n11064));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n11063));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n11062));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n11061));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n11060));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n11059));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n11058));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n11057));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n11056));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n11055));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n11054));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n11053));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n11052));   // coms.v(416[12] 543[6])
    SB_LUT4 i5_3_lut_4_lut_adj_690 (.I0(\data_out_frame2[9] [4]), .I1(\data_out_frame2[5] [6]), 
            .I2(\data_out_frame2[8] [6]), .I3(n17294), .O(n14_adj_2188));   // coms.v(229[16:299])
    defparam i5_3_lut_4_lut_adj_690.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n11051));   // coms.v(416[12] 543[6])
    SB_LUT4 i2_3_lut_4_lut_adj_691 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n10018), .I3(\FRAME_MATCHER.state[2] ), .O(n5815));
    defparam i2_3_lut_4_lut_adj_691.LUT_INIT = 16'h0102;
    SB_LUT4 i2_3_lut_4_lut_adj_692 (.I0(\data_out_frame2[9] [4]), .I1(\data_out_frame2[5] [6]), 
            .I2(n10371), .I3(n10530), .O(n17303));   // coms.v(229[16:299])
    defparam i2_3_lut_4_lut_adj_692.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n11050));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n11049));   // coms.v(416[12] 543[6])
    SB_LUT4 i2_3_lut_4_lut_adj_693 (.I0(\data_out[8][5] ), .I1(\data_out[8][6] ), 
            .I2(n10395), .I3(n17243), .O(data_out_9__3__N_356));   // coms.v(21[11:19])
    defparam i2_3_lut_4_lut_adj_693.LUT_INIT = 16'h9669;
    SB_LUT4 i11047_2_lut (.I0(n13662), .I1(tx_transmit_N_1947[2]), .I2(GND_net), 
            .I3(GND_net), .O(n13726));
    defparam i11047_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_694 (.I0(\data_out[8][5] ), .I1(\data_out[8][6] ), 
            .I2(data_out_6__1__N_537), .I3(GND_net), .O(n26_adj_2165));   // coms.v(21[11:19])
    defparam i1_2_lut_3_lut_adj_694.LUT_INIT = 16'h9696;
    SB_LUT4 i146_4_lut (.I0(n13726), .I1(n444), .I2(n9524), .I3(tx_transmit_N_1947[3]), 
            .O(n450));   // coms.v(335[6] 342[9])
    defparam i146_4_lut.LUT_INIT = 16'hcdcf;
    SB_LUT4 i1_2_lut_3_lut_adj_695 (.I0(\data_out_frame2[15] [0]), .I1(\data_out_frame2[16] [0]), 
            .I2(\data_out_frame2[13] [2]), .I3(GND_net), .O(n10440));   // coms.v(237[17:221])
    defparam i1_2_lut_3_lut_adj_695.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_696 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(n17206), .I3(GND_net), .O(n2137));   // coms.v(76[16:62])
    defparam i1_2_lut_3_lut_adj_696.LUT_INIT = 16'h9696;
    SB_LUT4 i149_3_lut (.I0(tx_transmit_N_1947[3]), .I1(n444), .I2(n9524), 
            .I3(GND_net), .O(n453));   // coms.v(360[6] 367[9])
    defparam i149_3_lut.LUT_INIT = 16'hcdcd;
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n11048));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n11047));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_28_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [28]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2233));
    defparam select_219_Select_28_i2_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n11046));   // coms.v(416[12] 543[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n11045));   // coms.v(416[12] 543[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame2[16] [7]), .I1(n17194), 
            .I2(\data_out_frame2[10] [5]), .I3(GND_net), .O(n10_adj_2297));   // coms.v(238[17:230])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n11044));   // coms.v(416[12] 543[6])
    SB_LUT4 select_217_Select_2_i4_3_lut (.I0(\FRAME_MATCHER.state_31__N_1406[2] ), 
            .I1(\FRAME_MATCHER.i_31__N_1273 ), .I2(n3779), .I3(GND_net), 
            .O(n4_adj_13));
    defparam select_217_Select_2_i4_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_697 (.I0(\UART_TRANSMITTER.state[1] ), .I1(n453), 
            .I2(n450), .I3(\UART_TRANSMITTER.state[0] ), .O(n4_adj_14));
    defparam i1_4_lut_adj_697.LUT_INIT = 16'h88d8;
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n11043));   // coms.v(416[12] 543[6])
    SB_LUT4 select_219_Select_29_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [29]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2231));
    defparam select_219_Select_29_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_698 (.I0(\FRAME_MATCHER.state[1] ), .I1(n9), 
            .I2(n10139), .I3(n31), .O(n11833));   // coms.v(416[12] 543[6])
    defparam i1_3_lut_4_lut_adj_698.LUT_INIT = 16'h2f0f;
    SB_LUT4 i1_2_lut_3_lut_adj_699 (.I0(\data_out_frame2[12] [4]), .I1(\data_out_frame2[12] [2]), 
            .I2(\data_out_frame2[8] [6]), .I3(GND_net), .O(n10334));   // coms.v(228[16:596])
    defparam i1_2_lut_3_lut_adj_699.LUT_INIT = 16'h9696;
    SB_LUT4 select_219_Select_30_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [30]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2229));
    defparam select_219_Select_30_i2_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n11042));   // coms.v(416[12] 543[6])
    SB_LUT4 add_977_22_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [20]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(n18008), .I3(n16098), .O(\FRAME_MATCHER.i_31__N_1278 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_22_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n11041));   // coms.v(416[12] 543[6])
    SB_LUT4 i8329_3_lut_4_lut (.I0(n15179), .I1(n17076), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n11015));
    defparam i8329_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n11040));   // coms.v(416[12] 543[6])
    SB_LUT4 i10541_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[2]), .O(n76[2]));
    defparam i10541_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 select_219_Select_31_i2_2_lut (.I0(\FRAME_MATCHER.i_31__N_1278 [31]), 
            .I1(n1034), .I2(GND_net), .I3(GND_net), .O(n2_adj_2225));
    defparam select_219_Select_31_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10543_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[1]), .O(n76[1]));
    defparam i10543_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_CARRY add_977_22 (.CI(n16098), .I0(\FRAME_MATCHER.i [20]), .I1(n18008), 
            .CO(n16099));
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n11036));   // coms.v(416[12] 543[6])
    SB_LUT4 i1_2_lut_adj_700 (.I0(\FRAME_MATCHER.state [3]), .I1(n17069), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2336));
    defparam i1_2_lut_adj_700.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n11035));   // coms.v(416[12] 543[6])
    SB_LUT4 add_977_21_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [19]), .I1(\FRAME_MATCHER.i [19]), 
            .I2(n18008), .I3(n16097), .O(\FRAME_MATCHER.i_31__N_1278 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_21_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_701 (.I0(n13146), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [28]));
    defparam i1_2_lut_adj_701.LUT_INIT = 16'h8888;
    SB_LUT4 i8384_3_lut_4_lut (.I0(n15179), .I1(n17076), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n11070));
    defparam i8384_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_3_lut_4_lut (.I0(n488), .I1(n13146), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(n9369), .O(n7_adj_2384));
    defparam i18_3_lut_4_lut.LUT_INIT = 16'h8f80;
    SB_CARRY add_977_21 (.CI(n16097), .I0(\FRAME_MATCHER.i [19]), .I1(n18008), 
            .CO(n16098));
    SB_LUT4 i1_4_lut_adj_702 (.I0(\FRAME_MATCHER.state[0] ), .I1(n29), .I2(n27_adj_2381), 
            .I3(n28_adj_2374), .O(n12491));   // coms.v(416[12] 543[6])
    defparam i1_4_lut_adj_702.LUT_INIT = 16'h5554;
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n11033));   // coms.v(416[12] 543[6])
    SB_LUT4 i10454_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[0]), .O(n76[0]));
    defparam i10454_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n11032));   // coms.v(416[12] 543[6])
    SB_LUT4 i3_4_lut_adj_703 (.I0(n10166), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n7_adj_2384), .O(n18285));
    defparam i3_4_lut_adj_703.LUT_INIT = 16'h4000;
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n11028));   // coms.v(416[12] 543[6])
    SB_CARRY delay_counter_2361_add_4_6 (.CI(n16069), .I0(GND_net), .I1(n76[4]), 
            .CO(n16070));
    SB_LUT4 mux_1507_i1_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(n3118[0]));   // coms.v(283[4] 369[11])
    defparam mux_1507_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i8385_3_lut_4_lut (.I0(n15179), .I1(n17076), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n11071));
    defparam i8385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1065_i1_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\rand_setpoint[25] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(\UART_TRANSMITTER.state[0] ), 
            .O(n2523[0]));   // coms.v(283[4] 369[11])
    defparam mux_1065_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i15053_2_lut (.I0(\rand_setpoint[17] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17626));   // coms.v(283[4] 369[11])
    defparam i15053_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_857_i1_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(n17626), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(data_out_6__1__N_537), 
            .O(n2243[0]));   // coms.v(283[4] 369[11])
    defparam mux_857_i1_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i8386_3_lut_4_lut (.I0(n15179), .I1(n17076), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n11072));
    defparam i8386_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_704 (.I0(\FRAME_MATCHER.state [5]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2335));
    defparam i1_2_lut_adj_704.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n11027));   // coms.v(416[12] 543[6])
    SB_LUT4 i8387_3_lut_4_lut (.I0(n15179), .I1(n17076), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n11073));
    defparam i8387_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15033_3_lut (.I0(\data_out[5][1] ), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(data_out_6__1__N_537), .I3(GND_net), .O(n17627));   // coms.v(283[4] 369[11])
    defparam i15033_3_lut.LUT_INIT = 16'h4848;
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n11025));   // coms.v(416[12] 543[6])
    SB_LUT4 mux_831_i1_4_lut (.I0(n17627), .I1(\rand_setpoint[18] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2208[0]));   // coms.v(283[4] 369[11])
    defparam mux_831_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i10522_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[13]), .O(n76[13]));
    defparam i10522_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 i1_2_lut_adj_705 (.I0(\FRAME_MATCHER.state [6]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2334));
    defparam i1_2_lut_adj_705.LUT_INIT = 16'h8888;
    SB_LUT4 i10527_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[12]), .O(n76[12]));
    defparam i10527_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n11024));   // coms.v(416[12] 543[6])
    SB_LUT4 i14999_3_lut (.I0(\data_out[5] [2]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5][1] ), .I3(GND_net), .O(n17631));   // coms.v(283[4] 369[11])
    defparam i14999_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i1_2_lut_3_lut_adj_706 (.I0(\data_out_frame2[8] [7]), .I1(\data_out_frame2[16] [3]), 
            .I2(\data_out_frame2[15] [3]), .I3(GND_net), .O(n17312));   // coms.v(239[17:230])
    defparam i1_2_lut_3_lut_adj_706.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n11023));   // coms.v(416[12] 543[6])
    SB_LUT4 i13368_2_lut (.I0(\FRAME_MATCHER.state [7]), .I1(n15821), .I2(GND_net), 
            .I3(GND_net), .O(n16141));   // coms.v(412[11:12])
    defparam i13368_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10659_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [29]));   // coms.v(430[13] 433[7])
    defparam i10659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10528_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[11]), .O(n76[11]));
    defparam i10528_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 i10531_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[10]), .O(n76[10]));
    defparam i10531_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 i10532_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[9]), .O(n76[9]));
    defparam i10532_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 i1_2_lut_adj_707 (.I0(\FRAME_MATCHER.state [8]), .I1(n8_adj_2385), 
            .I2(GND_net), .I3(GND_net), .O(n16666));
    defparam i1_2_lut_adj_707.LUT_INIT = 16'h8888;
    SB_LUT4 mux_805_i1_4_lut (.I0(n17631), .I1(\rand_setpoint[19] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2173[0]));   // coms.v(283[4] 369[11])
    defparam mux_805_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i10533_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[8]), .O(n76[8]));
    defparam i10533_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 i1_2_lut_adj_708 (.I0(\FRAME_MATCHER.state [9]), .I1(n8_adj_2385), 
            .I2(GND_net), .I3(GND_net), .O(n16674));
    defparam i1_2_lut_adj_708.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n11016));   // coms.v(416[12] 543[6])
    SB_LUT4 i10535_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[7]), .O(n76[7]));
    defparam i10535_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 i15145_3_lut (.I0(\data_out[5] [3]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [2]), .I3(GND_net), .O(n17639));   // coms.v(283[4] 369[11])
    defparam i15145_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i8388_3_lut_4_lut (.I0(n15179), .I1(n17076), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n11074));
    defparam i8388_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10658_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [30]));   // coms.v(430[13] 433[7])
    defparam i10658_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 delay_counter_2361_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[3]), .I3(n16068), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_779_i1_4_lut (.I0(n17639), .I1(\rand_setpoint[20] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n11[0]));   // coms.v(283[4] 369[11])
    defparam mux_779_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i10536_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[6]), .O(n76[6]));
    defparam i10536_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 i1_2_lut_adj_709 (.I0(\FRAME_MATCHER.state [11]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2333));
    defparam i1_2_lut_adj_709.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_710 (.I0(\data_out_frame2[10] [5]), .I1(\data_out_frame2[7] [1]), 
            .I2(\data_out_frame2[9] [0]), .I3(\data_out_frame2[12] [2]), 
            .O(n17288));   // coms.v(228[16:596])
    defparam i1_2_lut_4_lut_adj_710.LUT_INIT = 16'h6996;
    SB_LUT4 i15001_3_lut (.I0(\data_out[5] [4]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [3]), .I3(GND_net), .O(n17643));   // coms.v(283[4] 369[11])
    defparam i15001_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i1_2_lut_adj_711 (.I0(\FRAME_MATCHER.state [12]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n16708));
    defparam i1_2_lut_adj_711.LUT_INIT = 16'h8888;
    SB_LUT4 i10537_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[5]), .O(n76[5]));
    defparam i10537_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 mux_753_i1_4_lut (.I0(n17643), .I1(\rand_setpoint[21] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2103[0]));   // coms.v(283[4] 369[11])
    defparam mux_753_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i8389_3_lut_4_lut (.I0(n15179), .I1(n17076), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n11075));
    defparam i8389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_712 (.I0(\FRAME_MATCHER.state [13]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2332));
    defparam i1_2_lut_adj_712.LUT_INIT = 16'h8888;
    SB_LUT4 i15002_3_lut (.I0(\data_out[5] [5]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [4]), .I3(GND_net), .O(n17647));   // coms.v(283[4] 369[11])
    defparam i15002_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i10657_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [31]));   // coms.v(430[13] 433[7])
    defparam i10657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15004_2_lut_3_lut (.I0(\data_out_frame2[0] [2]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17586));
    defparam i15004_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 mux_727_i1_4_lut (.I0(n17647), .I1(\rand_setpoint[22] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2068[0]));   // coms.v(283[4] 369[11])
    defparam mux_727_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i15003_3_lut (.I0(data_out_7__3__N_441), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(n17126), .I3(GND_net), .O(n17651));   // coms.v(283[4] 369[11])
    defparam i15003_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 i1_2_lut_adj_713 (.I0(\FRAME_MATCHER.state [14]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2331));
    defparam i1_2_lut_adj_713.LUT_INIT = 16'h8888;
    SB_LUT4 i8390_3_lut_4_lut (.I0(n15179), .I1(n17076), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n11076));
    defparam i8390_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10687_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [1]));   // coms.v(430[13] 433[7])
    defparam i10687_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_714 (.I0(\data_out_frame2[12] [5]), .I1(\data_out_frame2[13] [5]), 
            .I2(\data_out_frame2[10] [7]), .I3(GND_net), .O(n17255));   // coms.v(232[16:229])
    defparam i1_2_lut_3_lut_adj_714.LUT_INIT = 16'h9696;
    SB_LUT4 mux_701_i1_4_lut (.I0(n17651), .I1(\rand_setpoint[23] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2033[0]));   // coms.v(283[4] 369[11])
    defparam mux_701_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i10686_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n13146), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [2]));   // coms.v(430[13] 433[7])
    defparam i10686_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_715 (.I0(\FRAME_MATCHER.state [15]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2330));
    defparam i1_2_lut_adj_715.LUT_INIT = 16'h8888;
    SB_LUT4 i10538_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[4]), .O(n76[4]));
    defparam i10538_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15321 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [6]), .I2(\data_out_frame2[19] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n18112));
    defparam byte_transmit_counter2_0__bdd_4_lut_15321.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_716 (.I0(\FRAME_MATCHER.state [16]), .I1(n8_adj_2385), 
            .I2(GND_net), .I3(GND_net), .O(n16670));
    defparam i1_2_lut_adj_716.LUT_INIT = 16'h8888;
    SB_LUT4 i10539_2_lut_3_lut_4_lut (.I0(n9453), .I1(n16267), .I2(n444), 
            .I3(delay_counter[3]), .O(n76[3]));
    defparam i10539_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_LUT4 i260_2_lut_3_lut (.I0(n488), .I1(n13146), .I2(\FRAME_MATCHER.i_31__N_1272 ), 
            .I3(GND_net), .O(n276));
    defparam i260_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i15044_4_lut (.I0(n17129), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [5]), .I3(n10326), .O(n17653));   // coms.v(283[4] 369[11])
    defparam i15044_4_lut.LUT_INIT = 16'h4884;
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n11015));   // coms.v(416[12] 543[6])
    SB_LUT4 mux_675_i1_4_lut (.I0(n17653), .I1(\rand_setpoint[8] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n1998[0]));   // coms.v(283[4] 369[11])
    defparam mux_675_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_3_lut_adj_717 (.I0(\data_out_frame2[10] [1]), .I1(\data_out_frame2[11] [7]), 
            .I2(\data_out_frame2[14] [5]), .I3(GND_net), .O(n17234));   // coms.v(227[16:31])
    defparam i1_2_lut_3_lut_adj_717.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_718 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [4]), .O(n16716));
    defparam i1_2_lut_4_lut_adj_718.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_adj_719 (.I0(\FRAME_MATCHER.state [18]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2329));   // coms.v(416[12] 543[6])
    defparam i1_2_lut_adj_719.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_720 (.I0(\data_out[5] [2]), .I1(\data_out[5][1] ), 
            .I2(data_out_6__1__N_537), .I3(GND_net), .O(n10326));   // coms.v(130[17:68])
    defparam i2_3_lut_adj_720.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_721 (.I0(\data_out_frame2[12] [7]), .I1(\data_out_frame2[16] [5]), 
            .I2(\data_out_frame2[12] [0]), .I3(\data_out_frame2[14] [6]), 
            .O(n17225));   // coms.v(228[16:596])
    defparam i2_3_lut_4_lut_adj_721.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_722 (.I0(\data_out_frame2[5] [0]), .I1(\data_out_frame2[15] [4]), 
            .I2(\data_out_frame2[6] [6]), .I3(\data_out_frame2[8] [5]), 
            .O(n17309));   // coms.v(228[16:596])
    defparam i1_2_lut_4_lut_adj_722.LUT_INIT = 16'h6996;
    SB_LUT4 i15142_3_lut (.I0(n17126), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [5]), .I3(GND_net), .O(n17574));   // coms.v(283[4] 369[11])
    defparam i15142_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i14552_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[1] ), .I1(n13662), 
            .I2(tx_transmit_N_1947[2]), .I3(GND_net), .O(n17327));
    defparam i14552_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_723 (.I0(\FRAME_MATCHER.state [19]), .I1(n15821), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2328));
    defparam i1_2_lut_adj_723.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_724 (.I0(\data_out_frame2[5] [4]), .I1(n10_adj_2207), 
            .I2(\data_out_frame2[13] [4]), .I3(\data_out_frame2[9] [0]), 
            .O(n17095));   // coms.v(230[16:237])
    defparam i5_3_lut_4_lut_adj_724.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_725 (.I0(n15821), .I1(\FRAME_MATCHER.state [20]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2327));
    defparam i1_2_lut_adj_725.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_726 (.I0(n1034), .I1(rx_data_ready), .I2(\FRAME_MATCHER.i [1]), 
            .I3(n15164), .O(n17072));
    defparam i1_3_lut_4_lut_adj_726.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_4_lut_adj_727 (.I0(\data_out[9] [5]), .I1(\data_out[6] [3]), 
            .I2(\data_out[6] [1]), .I3(n10183), .O(n17252));   // coms.v(175[16:77])
    defparam i1_2_lut_4_lut_adj_727.LUT_INIT = 16'h6996;
    SB_LUT4 add_977_20_lut (.I0(\FRAME_MATCHER.i_31__N_1310 [18]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(n18008), .I3(n16096), .O(\FRAME_MATCHER.i_31__N_1278 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_977_20_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mux_649_i1_4_lut (.I0(n17574), .I1(\rand_setpoint[9] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n1963[0]));   // coms.v(283[4] 369[11])
    defparam mux_649_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_adj_728 (.I0(\FRAME_MATCHER.state [21]), .I1(n8_adj_2385), 
            .I2(GND_net), .I3(GND_net), .O(n16686));
    defparam i1_2_lut_adj_728.LUT_INIT = 16'h8888;
    SB_LUT4 i14993_2_lut (.I0(\rand_setpoint[10] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17583));   // coms.v(283[4] 369[11])
    defparam i14993_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_729 (.I0(\data_out_frame2[13] [1]), .I1(\data_out_frame2[15] [0]), 
            .I2(\data_out_frame2[5] [5]), .I3(n10223), .O(n14_adj_2206));
    defparam i5_3_lut_4_lut_adj_729.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_730 (.I0(n1034), .I1(rx_data_ready), .I2(\FRAME_MATCHER.i [1]), 
            .I3(n15164), .O(n17076));
    defparam i1_3_lut_4_lut_adj_730.LUT_INIT = 16'hfff7;
    SB_LUT4 mux_623_i1_4_lut (.I0(data_out_7__2__N_447), .I1(n17583), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n1928[0]));   // coms.v(283[4] 369[11])
    defparam mux_623_i1_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i2_3_lut_4_lut_adj_731 (.I0(\data_out[9] [4]), .I1(\data_out[10][0] ), 
            .I2(\data_out[6] [2]), .I3(\data_out[6] [0]), .O(n17177));   // coms.v(174[16:77])
    defparam i2_3_lut_4_lut_adj_731.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_732 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [31]), .O(n16700));
    defparam i1_2_lut_4_lut_adj_732.LUT_INIT = 16'hf400;
    SB_LUT4 i3_4_lut_adj_733 (.I0(tx_transmit_N_1947[6]), .I1(tx_transmit_N_1947[4]), 
            .I2(tx_transmit_N_1947[5]), .I3(tx_transmit_N_1947[7]), .O(n9524));   // coms.v(336[10:53])
    defparam i3_4_lut_adj_733.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_734 (.I0(\data_out_frame2[16] [1]), .I1(\data_out_frame2[9] [1]), 
            .I2(\data_out_frame2[13] [3]), .I3(n10346), .O(n17231));   // coms.v(227[16:31])
    defparam i2_3_lut_4_lut_adj_734.LUT_INIT = 16'h6996;
    SB_LUT4 i8376_3_lut_4_lut (.I0(n15171), .I1(n17076), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n11062));
    defparam i8376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_735 (.I0(\data_out_frame2[8] [7]), .I1(\data_out_frame2[12] [3]), 
            .I2(\data_out_frame2[5] [3]), .I3(GND_net), .O(n6_adj_2197));
    defparam i1_2_lut_3_lut_adj_735.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_736 (.I0(n9524), .I1(tx_transmit_N_1947[2]), .I2(tx_transmit_N_1947[3]), 
            .I3(n13662), .O(n16267));
    defparam i2_4_lut_adj_736.LUT_INIT = 16'hfefa;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut (.I0(n18163), .I1(\data_out_frame2[20] [0]), 
            .I2(byte_transmit_counter2[2]), .I3(n9157), .O(n22_adj_2387));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_737 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [10]), .O(n16710));
    defparam i1_2_lut_4_lut_adj_737.LUT_INIT = 16'hf400;
    SB_LUT4 i8377_3_lut_4_lut (.I0(n15171), .I1(n17076), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n11063));
    defparam i8377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[2] [7]), .O(n22_adj_2201));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h9f6f;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i31_4_lut (.I0(n18229), .I1(n22_adj_2387), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[0]));   // coms.v(403[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out[6] [3]), 
            .I1(\data_out[7] [3]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_c));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10706_2_lut (.I0(\FRAME_MATCHER.state [23]), .I1(n15821), .I2(GND_net), 
            .I3(GND_net), .O(n13381));
    defparam i10706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_738 (.I0(\data_out[7] [3]), .I1(\data_out[5] [3]), 
            .I2(\data_out[5] [4]), .I3(\data_out[9][2] ), .O(n17162));   // coms.v(171[16:355])
    defparam i1_2_lut_4_lut_adj_738.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_739 (.I0(n44), .I1(n9334), .I2(n4_c), .I3(n47_adj_2347), 
            .O(n15821));
    defparam i1_3_lut_4_lut_adj_739.LUT_INIT = 16'hfff4;
    SB_LUT4 i8349_3_lut_4_lut (.I0(n39), .I1(n17076), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n11035));
    defparam i8349_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8378_3_lut_4_lut (.I0(n15171), .I1(n17076), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n11064));
    defparam i8378_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8379_3_lut_4_lut (.I0(n15171), .I1(n17076), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n11065));
    defparam i8379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8380_3_lut_4_lut (.I0(n15171), .I1(n17076), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n11066));
    defparam i8380_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_2_lut (.I0(delay_counter[8]), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_2388));   // coms.v(306[11:30])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_3_lut_4_lut_adj_740 (.I0(\data_out_frame2[13] [0]), .I1(n10263), 
            .I2(n10_adj_2190), .I3(n17279), .O(n17281));   // coms.v(228[16:596])
    defparam i5_3_lut_4_lut_adj_740.LUT_INIT = 16'h6996;
    SB_LUT4 i8381_3_lut_4_lut (.I0(n15171), .I1(n17076), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n11067));
    defparam i8381_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_741 (.I0(delay_counter[7]), .I1(delay_counter[12]), 
            .I2(delay_counter[11]), .I3(delay_counter[4]), .O(n24_adj_2389));   // coms.v(306[11:30])
    defparam i10_4_lut_adj_741.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_742 (.I0(\data_out[9] [0]), .I1(\data_out[7] [1]), 
            .I2(\data_out[5] [2]), .I3(\data_out[6] [7]), .O(n10196));   // coms.v(181[17:93])
    defparam i2_3_lut_4_lut_adj_742.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_743 (.I0(delay_counter[6]), .I1(delay_counter[0]), 
            .I2(delay_counter[10]), .I3(delay_counter[13]), .O(n22_adj_2390));   // coms.v(306[11:30])
    defparam i8_4_lut_adj_743.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_744 (.I0(delay_counter[2]), .I1(n24_adj_2389), 
            .I2(n18_adj_2388), .I3(delay_counter[5]), .O(n26_adj_2391));   // coms.v(306[11:30])
    defparam i12_4_lut_adj_744.LUT_INIT = 16'hfffe;
    SB_LUT4 n18112_bdd_4_lut (.I0(n18112), .I1(\data_out_frame2[17] [6]), 
            .I2(\data_out_frame2[16] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n18115));
    defparam n18112_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8382_3_lut_4_lut (.I0(n15171), .I1(n17076), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n11068));
    defparam i8382_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_745 (.I0(\data_out[5] [3]), .I1(\data_out[5] [4]), 
            .I2(\data_out[9][2] ), .I3(GND_net), .O(n17270));   // coms.v(177[16:77])
    defparam i1_2_lut_3_lut_adj_745.LUT_INIT = 16'h9696;
    SB_LUT4 i8383_3_lut_4_lut (.I0(n15171), .I1(n17076), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n11069));
    defparam i8383_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15108_2_lut (.I0(\data_out[5] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17703));
    defparam i15108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_746 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [17]), .O(n16704));
    defparam i1_2_lut_4_lut_adj_746.LUT_INIT = 16'hf400;
    SB_LUT4 i5_3_lut_4_lut_adj_747 (.I0(\data_out_frame2[0] [3]), .I1(\data_out_frame2[14] [3]), 
            .I2(\data_out_frame2[7] [3]), .I3(\data_out_frame2[0] [4]), 
            .O(n14));   // coms.v(232[16:229])
    defparam i5_3_lut_4_lut_adj_747.LUT_INIT = 16'h6996;
    SB_LUT4 i8350_3_lut_4_lut (.I0(n39), .I1(n17076), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n11036));
    defparam i8350_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13_4_lut_adj_748 (.I0(delay_counter[1]), .I1(n26_adj_2391), 
            .I2(n22_adj_2390), .I3(delay_counter[9]), .O(n9453));   // coms.v(306[11:30])
    defparam i13_4_lut_adj_748.LUT_INIT = 16'hfffe;
    SB_LUT4 i8368_3_lut_4_lut (.I0(n15179), .I1(n17072), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n11054));
    defparam i8368_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_749 (.I0(\data_out[9] [1]), .I1(\data_out[9] [0]), 
            .I2(n10_adj_2172), .I3(n17264), .O(data_out_9__6__N_324));   // coms.v(184[17:86])
    defparam i5_3_lut_4_lut_adj_749.LUT_INIT = 16'h9669;
    SB_LUT4 i8354_3_lut_4_lut (.I0(n39), .I1(n17076), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n11040));
    defparam i8354_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8369_3_lut_4_lut (.I0(n15179), .I1(n17072), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n11055));
    defparam i8369_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8370_3_lut_4_lut (.I0(n15179), .I1(n17072), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n11056));
    defparam i8370_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_750 (.I0(n13146), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1310 [3]));
    defparam i1_2_lut_adj_750.LUT_INIT = 16'h8888;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_out_frame2[15] [6]), .I1(\data_out_frame2[7] [5]), 
            .I2(\data_out_frame2[0] [5]), .I3(\data_out_frame2[8] [1]), 
            .O(n20));   // coms.v(234[16:291])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8371_3_lut_4_lut (.I0(n15179), .I1(n17072), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n11057));
    defparam i8371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_751 (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n10018), .I3(GND_net), .O(n9));
    defparam i1_2_lut_3_lut_adj_751.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_752 (.I0(\FRAME_MATCHER.state [28]), .I1(n4_adj_2135), 
            .I2(GND_net), .I3(GND_net), .O(n16748));
    defparam i1_2_lut_adj_752.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_753 (.I0(n5_adj_8), .I1(n17069), .I2(\FRAME_MATCHER.state[1] ), 
            .I3(n9334), .O(n8_adj_2385));
    defparam i1_4_lut_adj_753.LUT_INIT = 16'hcdcc;
    SB_LUT4 i1_2_lut_adj_754 (.I0(\FRAME_MATCHER.state [29]), .I1(n8_adj_2385), 
            .I2(GND_net), .I3(GND_net), .O(n16658));
    defparam i1_2_lut_adj_754.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15316 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [5]), .I2(\data_out_frame2[11] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n18106));
    defparam byte_transmit_counter2_0__bdd_4_lut_15316.LUT_INIT = 16'he4aa;
    SB_LUT4 i8372_3_lut_4_lut (.I0(n15179), .I1(n17072), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n11058));
    defparam i8372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_755 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [22]), .O(n16714));
    defparam i1_2_lut_4_lut_adj_755.LUT_INIT = 16'hf400;
    SB_LUT4 i2_3_lut_4_lut_adj_756 (.I0(n13628), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(tx2_active), .I3(r_SM_Main_2__N_2034_adj_2405[0]), .O(n16261));   // coms.v(434[4] 542[11])
    defparam i2_3_lut_4_lut_adj_756.LUT_INIT = 16'hfffb;
    SB_LUT4 i8359_3_lut_4_lut (.I0(n39), .I1(n17076), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n11045));
    defparam i8359_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_757 (.I0(\FRAME_MATCHER.state [29]), .I1(n4_adj_2135), 
            .I2(GND_net), .I3(GND_net), .O(n16746));
    defparam i1_2_lut_adj_757.LUT_INIT = 16'h8888;
    SB_LUT4 i8373_3_lut_4_lut (.I0(n15179), .I1(n17072), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n11059));
    defparam i8373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8355_3_lut_4_lut (.I0(n39), .I1(n17076), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n11041));
    defparam i8355_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_758 (.I0(\FRAME_MATCHER.state [30]), .I1(n4_adj_2135), 
            .I2(GND_net), .I3(GND_net), .O(n16744));
    defparam i1_2_lut_adj_758.LUT_INIT = 16'h8888;
    SB_LUT4 i8374_3_lut_4_lut (.I0(n15179), .I1(n17072), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n11060));
    defparam i8374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_759 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [24]), .O(n16688));
    defparam i1_2_lut_4_lut_adj_759.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_4_lut_adj_760 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [25]), .O(n16690));
    defparam i1_2_lut_4_lut_adj_760.LUT_INIT = 16'hf400;
    SB_CARRY delay_counter_2361_add_4_5 (.CI(n16068), .I0(GND_net), .I1(n76[3]), 
            .CO(n16069));
    SB_LUT4 i8375_3_lut_4_lut (.I0(n15179), .I1(n17072), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n11061));
    defparam i8375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14998_2_lut (.I0(\rand_setpoint[11] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17585));   // coms.v(283[4] 369[11])
    defparam i14998_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_761 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [26]), .O(n16702));
    defparam i1_2_lut_4_lut_adj_761.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_4_lut_adj_762 (.I0(\FRAME_MATCHER.i_31__N_1273 ), .I1(n3779), 
            .I2(n13146), .I3(n47_adj_2347), .O(n17069));
    defparam i1_2_lut_4_lut_adj_762.LUT_INIT = 16'hff20;
    SB_LUT4 mux_597_i1_4_lut (.I0(data_out_7__3__N_441), .I1(n17585), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n1893[0]));   // coms.v(283[4] 369[11])
    defparam mux_597_i1_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1_2_lut_adj_763 (.I0(n11833), .I1(byte_transmit_counter2[0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2187));   // coms.v(409[11:16])
    defparam i1_2_lut_adj_763.LUT_INIT = 16'h8888;
    SB_LUT4 i8356_3_lut_4_lut (.I0(n39), .I1(n17076), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n11042));
    defparam i8356_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_224_Select_0_i2_4_lut (.I0(byte_transmit_counter2[0]), 
            .I1(\FRAME_MATCHER.i_31__N_1272 ), .I2(n17659), .I3(n11867), 
            .O(n2_adj_2186));
    defparam select_224_Select_0_i2_4_lut.LUT_INIT = 16'h88c0;
    SB_LUT4 i1_2_lut_4_lut_adj_764 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [27]), .O(n16718));
    defparam i1_2_lut_4_lut_adj_764.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_4_lut_adj_765 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [28]), .O(n16696));
    defparam i1_2_lut_4_lut_adj_765.LUT_INIT = 16'hf400;
    SB_DFFSS byte_transmit_counter2_i6 (.Q(byte_transmit_counter2[6]), .C(CLK_c), 
            .D(n2_adj_2326), .S(n4_adj_2325));   // coms.v(416[12] 543[6])
    SB_LUT4 i10986_2_lut (.I0(tx_transmit_N_1947[0]), .I1(tx_transmit_N_1947[1]), 
            .I2(GND_net), .I3(GND_net), .O(n13662));
    defparam i10986_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_766 (.I0(\UART_TRANSMITTER.state[0] ), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(n4650));
    defparam i2_3_lut_adj_766.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut_adj_767 (.I0(n44), .I1(n9334), .I2(n17069), 
            .I3(\FRAME_MATCHER.state [30]), .O(n16698));
    defparam i1_2_lut_4_lut_adj_767.LUT_INIT = 16'hf400;
    SB_LUT4 i1_3_lut_adj_768 (.I0(\UART_TRANSMITTER.state[1] ), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(tx_transmit_N_1947[2]), .I3(GND_net), .O(n65));   // coms.v(283[4] 369[11])
    defparam i1_3_lut_adj_768.LUT_INIT = 16'hcece;
    SB_LUT4 delay_counter_2361_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n76[2]), .I3(n16067), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2361_add_4_4_lut.LUT_INIT = 16'hC33C;
    uart_tx tx (.n10969(n10969), .n10966(n10966), .n10963(n10963), .n10960(n10960), 
            .n10957(n10957), .GND_net(GND_net), .n10954(n10954), .n10951(n10951), 
            .n10994(n10994), .VCC_net(VCC_net), .\r_Bit_Index[2] (\r_Bit_Index[2] ), 
            .n16932(n16932), .r_Tx_Data({r_Tx_Data}), .CLK_c(CLK_c), .n16930(n16930), 
            .n16928(n16928), .n16926(n16926), .\r_Bit_Index[1] (\r_Bit_Index[1] ), 
            .n10953(n10953), .n10956(n10956), .n10959(n10959), .n10962(n10962), 
            .n10965(n10965), .n10968(n10968), .n10971(n10971), .n10974(n10974), 
            .n16924(n16924), .n10996(n10996), .\r_SM_Main_2__N_2034[0] (r_SM_Main_2__N_2034[0]), 
            .n16914(n16914), .n16902(n16902), .n18199(n18199), .n18073(n18073), 
            .tx_o(tx_o), .tx_active(tx_active), .n9257(n9257), .n16912(n16912), 
            .n5142(n5142), .tx_active_prev(tx_active_prev), .n65(n65_adj_2192), 
            .n10972(n10972), .tx_enable(tx_enable), .n444(n444)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(259[10:70])
    uart_tx_U0 tx2 (.\r_SM_Main_2__N_2031[1] (\r_SM_Main_2__N_2031[1] ), .r_SM_Main({r_SM_Main}), 
            .\r_SM_Main_2__N_2034[0] (r_SM_Main_2__N_2034_adj_2405[0]), .n4(n4_adj_15), 
            .GND_net(GND_net), .r_Bit_Index({r_Bit_Index}), .n18280(n18280), 
            .CLK_c(CLK_c), .n10674(n10674), .n10920(n10920), .n10923(n10923), 
            .n10977(n10977), .tx2_data({tx2_data}), .n5266(n5266), .n17412(n17412), 
            .n10976(n10976), .VCC_net(VCC_net), .n3(n3), .n8191(n8191), 
            .n11039(n11039), .n11038(n11038), .tx2_active(tx2_active), 
            .n11037(n11037), .tx2_o(tx2_o), .tx2_enable(tx2_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(404[10:77])
    uart_rx rx (.r_Bit_Index({r_Bit_Index_adj_27}), .n5244(n5244), .GND_net(GND_net), 
            .\r_SM_Main[1] (\r_SM_Main[1]_adj_21 ), .\r_SM_Main[2] (\r_SM_Main[2]_adj_22 ), 
            .n17361(n17361), .CLK_c(CLK_c), .n10983(n10983), .rx_data_ready(rx_data_ready), 
            .n11019(n11019), .n11031(n11031), .r_Rx_Data(r_Rx_Data), .rx_i(rx_i), 
            .n11139(n11139), .rx_data({rx_data}), .n13744(n13744), .n11136(n11136), 
            .n11135(n11135), .n1(n1_adj_23), .n13116(n13116), .n11112(n11112), 
            .n4(n4_adj_24), .n11090(n11090), .n11089(n11089), .n18008(n18008), 
            .n11034(n11034), .n11026(n11026), .VCC_net(VCC_net), .n10987(n10987), 
            .n13692(n13692), .n11018(n11018), .n4_adj_1(n4_adj_25), .n9999(n9999), 
            .n17708(n17708), .n17707(n17707), .n4_adj_2(n4_adj_26), .n10010(n10010)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(376[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n10969, n10966, n10963, n10960, n10957, GND_net, 
            n10954, n10951, n10994, VCC_net, \r_Bit_Index[2] , n16932, 
            r_Tx_Data, CLK_c, n16930, n16928, n16926, \r_Bit_Index[1] , 
            n10953, n10956, n10959, n10962, n10965, n10968, n10971, 
            n10974, n16924, n10996, \r_SM_Main_2__N_2034[0] , n16914, 
            n16902, n18199, n18073, tx_o, tx_active, n9257, n16912, 
            n5142, tx_active_prev, n65, n10972, tx_enable, n444) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output n10969;
    output n10966;
    output n10963;
    output n10960;
    output n10957;
    input GND_net;
    output n10954;
    output n10951;
    output n10994;
    input VCC_net;
    output \r_Bit_Index[2] ;
    input n16932;
    output [7:0]r_Tx_Data;
    input CLK_c;
    input n16930;
    input n16928;
    input n16926;
    output \r_Bit_Index[1] ;
    input n10953;
    input n10956;
    input n10959;
    input n10962;
    input n10965;
    input n10968;
    input n10971;
    input n10974;
    input n16924;
    input n10996;
    input \r_SM_Main_2__N_2034[0] ;
    input n16914;
    input n16902;
    input n18199;
    input n18073;
    output tx_o;
    output tx_active;
    output n9257;
    input n16912;
    output n5142;
    input tx_active_prev;
    output n65;
    output n10972;
    output tx_enable;
    output n444;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n16123, n16124, n16122, n16121, n16120, n16119, n10688;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n16830, n16118, n16117, n10, n77, n83, n55, n11285, 
        n11284, n6759, n11140, n11137, n31, n12, n10_adj_2133, 
        n13702, n10613, n11021, n17673, n12_adj_2134, n16910;
    
    SB_LUT4 add_59_9_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[7]), 
            .I2(r_SM_Main[2]), .I3(n16123), .O(n10969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_9 (.CI(n16123), .I0(r_Clock_Count[7]), .I1(r_SM_Main[2]), 
            .CO(n16124));
    SB_LUT4 add_59_8_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[6]), 
            .I2(r_SM_Main[2]), .I3(n16122), .O(n10966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_8 (.CI(n16122), .I0(r_Clock_Count[6]), .I1(r_SM_Main[2]), 
            .CO(n16123));
    SB_LUT4 add_59_7_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[5]), 
            .I2(r_SM_Main[2]), .I3(n16121), .O(n10963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_7 (.CI(n16121), .I0(r_Clock_Count[5]), .I1(r_SM_Main[2]), 
            .CO(n16122));
    SB_LUT4 add_59_6_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[4]), 
            .I2(r_SM_Main[2]), .I3(n16120), .O(n10960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_6 (.CI(n16120), .I0(r_Clock_Count[4]), .I1(r_SM_Main[2]), 
            .CO(n16121));
    SB_LUT4 add_59_5_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[3]), 
            .I2(r_SM_Main[2]), .I3(n16119), .O(n10957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i12_3_lut (.I0(n10688), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n16830));   // verilog/uart_tx.v(31[16:25])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_CARRY add_59_5 (.CI(n16119), .I0(r_Clock_Count[3]), .I1(r_SM_Main[2]), 
            .CO(n16120));
    SB_LUT4 add_59_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[2]), 
            .I2(r_SM_Main[2]), .I3(n16118), .O(n10954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_4 (.CI(n16118), .I0(r_Clock_Count[2]), .I1(r_SM_Main[2]), 
            .CO(n16119));
    SB_LUT4 add_59_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[1]), 
            .I2(r_SM_Main[2]), .I3(n16117), .O(n10951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_3 (.CI(n16117), .I0(r_Clock_Count[1]), .I1(r_SM_Main[2]), 
            .CO(n16118));
    SB_LUT4 add_59_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[0]), 
            .I2(r_SM_Main[2]), .I3(VCC_net), .O(n10994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(r_SM_Main[2]), 
            .CO(n16117));
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[3]), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[1]), .I1(n10), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n77));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i101_4_lut (.I0(r_Clock_Count[7]), .I1(n77), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[8]), .O(n83));   // verilog/uart_tx.v(32[16:29])
    defparam i101_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(n83), .O(n10688));
    defparam i1_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i12034_4_lut (.I0(n10688), .I1(n55), .I2(r_SM_Main[1]), .I3(\r_Bit_Index[2] ), 
            .O(n11285));   // verilog/uart_tx.v(31[16:25])
    defparam i12034_4_lut.LUT_INIT = 16'h35c0;
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .D(n16932));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .D(n16930));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .D(n16928));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .D(n16926));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(\r_Bit_Index[2] ), .C(CLK_c), .D(n11285));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(\r_Bit_Index[1] ), .C(CLK_c), .D(n11284));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .D(n10953));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .D(n10956));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .D(n10959));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .D(n10962));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .D(n10965));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .D(n10968));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .D(n10971));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .D(n10974));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .D(n16924));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n16830));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .D(n10996));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_2034[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n6759));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .D(n16914));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(VCC_net), .D(n16902));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n11140));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n11137));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i33_3_lut (.I0(n18199), .I1(n18073), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n31));   // verilog/uart_tx.v(33[16:27])
    defparam i33_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26_3_lut (.I0(n31), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n12));
    defparam i26_3_lut.LUT_INIT = 16'h1c1c;
    SB_LUT4 i25_3_lut (.I0(n12), .I1(tx_o), .I2(r_SM_Main[2]), .I3(GND_net), 
            .O(n10_adj_2133));
    defparam i25_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_4_lut_adj_399 (.I0(r_SM_Main[2]), .I1(n6759), .I2(n13702), 
            .I3(r_SM_Main[1]), .O(n10613));
    defparam i1_4_lut_adj_399.LUT_INIT = 16'h5044;
    SB_LUT4 i10020_3_lut (.I0(n10613), .I1(r_SM_Main[1]), .I2(tx_active), 
            .I3(GND_net), .O(n11021));   // verilog/uart_tx.v(31[16:25])
    defparam i10020_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i15099_4_lut (.I0(r_Bit_Index[0]), .I1(\r_Bit_Index[1] ), .I2(\r_Bit_Index[2] ), 
            .I3(n83), .O(n17673));   // verilog/uart_tx.v(31[16:25])
    defparam i15099_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i29_3_lut (.I0(\r_SM_Main_2__N_2034[0] ), .I1(n17673), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n12_adj_2134));   // verilog/uart_tx.v(31[16:25])
    defparam i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_400 (.I0(r_SM_Main[2]), .I1(n12_adj_2134), .I2(n83), 
            .I3(r_SM_Main[0]), .O(n16910));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut_adj_400.LUT_INIT = 16'h0544;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_SM_Main[1]), .I1(n83), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main[0]), .O(n11140));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i11999_4_lut_4_lut (.I0(n83), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n11137));   // verilog/uart_tx.v(31[16:25])
    defparam i11999_4_lut_4_lut.LUT_INIT = 16'h1320;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main_2__N_2034[0] ), .O(n9257));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .D(n16912));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(n83), .O(n5142));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h3301;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n16910));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n11021));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .D(n10_adj_2133));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i12039_4_lut_4_lut (.I0(r_Bit_Index[0]), .I1(n10688), .I2(\r_Bit_Index[1] ), 
            .I3(r_SM_Main[1]), .O(n11284));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12039_4_lut_4_lut.LUT_INIT = 16'h7830;
    SB_LUT4 i1_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(n10688), .I2(\r_Bit_Index[1] ), 
            .I3(GND_net), .O(n55));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_401 (.I0(tx_active), .I1(tx_active_prev), .I2(GND_net), 
            .I3(GND_net), .O(n65));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_401.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_402 (.I0(r_SM_Main[0]), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n13702));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_402.LUT_INIT = 16'h8888;
    SB_LUT4 add_59_10_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[8]), 
            .I2(r_SM_Main[2]), .I3(n16124), .O(n10972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_403 (.I0(tx_active), .I1(\r_SM_Main_2__N_2034[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n444));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_403.LUT_INIT = 16'heeee;
    
endmodule
//
// Verilog Description of module uart_tx_U0
//

module uart_tx_U0 (\r_SM_Main_2__N_2031[1] , r_SM_Main, \r_SM_Main_2__N_2034[0] , 
            n4, GND_net, r_Bit_Index, n18280, CLK_c, n10674, n10920, 
            n10923, n10977, tx2_data, n5266, n17412, n10976, VCC_net, 
            n3, n8191, n11039, n11038, tx2_active, n11037, tx2_o, 
            tx2_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output \r_SM_Main_2__N_2031[1] ;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_2034[0] ;
    output n4;
    input GND_net;
    output [2:0]r_Bit_Index;
    input n18280;
    input CLK_c;
    output n10674;
    input n10920;
    input n10923;
    input n10977;
    input [7:0]tx2_data;
    output n5266;
    output n17412;
    output n10976;
    input VCC_net;
    output n3;
    output n8191;
    input n11039;
    input n11038;
    output tx2_active;
    input n11037;
    output tx2_o;
    output tx2_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n17018, n10;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n18232, n18235;
    wire [8:0]n312;
    
    wire n10852, n18082, n18085, n9269, n16139, n16138, n13614, 
        n16137, n16136, n16135, n16134, n13748, n17322, n16133, 
        n16132, n11144, o_Tx_Serial_N_2062;
    
    SB_LUT4 i15179_4_lut_4_lut (.I0(\r_SM_Main_2__N_2031[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_2034[0] ), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i15179_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 i2_3_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n17018));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[4]), 
            .I3(r_Clock_Count[3]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n18232));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n18232_bdd_4_lut (.I0(n18232), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n18235));
    defparam n18232_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n18280));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n10674), 
            .D(n312[1]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n10674), 
            .D(n312[2]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n10674), 
            .D(n312[3]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n10674), 
            .D(n312[4]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n10674), 
            .D(n312[5]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n10674), 
            .D(n312[6]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n10674), 
            .D(n312[7]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n10674), 
            .D(n312[8]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .D(n10920));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_15415 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n18082));
    defparam r_Bit_Index_0__bdd_4_lut_15415.LUT_INIT = 16'he4aa;
    SB_LUT4 n18082_bdd_4_lut (.I0(n18082), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n18085));
    defparam n18082_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .D(n10923));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n10674), 
            .D(n312[0]), .R(n10852));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n10977));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n9269), .D(tx2_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n16139), .O(n312[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n16138), .O(n312[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_9 (.CI(n16138), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n16139));
    SB_LUT4 i2615_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5266));   // verilog/uart_tx.v(98[36:51])
    defparam i2615_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14643_3_lut (.I0(n17412), .I1(n13614), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n10976));
    defparam i14643_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n16137), .O(n312[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_8 (.CI(n16137), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n16138));
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n16136), .O(n312[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n16136), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n16137));
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n16135), .O(n312[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_6 (.CI(n16135), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n16136));
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n16134), .O(n312[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11067_2_lut_4_lut (.I0(r_Clock_Count[1]), .I1(n10), .I2(r_Clock_Count[5]), 
            .I3(r_SM_Main[2]), .O(n13748));
    defparam i11067_2_lut_4_lut.LUT_INIT = 16'hff80;
    SB_CARRY add_59_5 (.CI(n16134), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n16135));
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[0]), .I1(n17018), .I2(n13748), .I3(r_SM_Main[1]), 
            .O(n17322));
    defparam i1_4_lut.LUT_INIT = 16'h0302;
    SB_LUT4 i15218_2_lut (.I0(r_SM_Main[2]), .I1(n17322), .I2(GND_net), 
            .I3(GND_net), .O(n10852));
    defparam i15218_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n16133), .O(n312[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_Clock_Count[1]), .I1(n10), .I2(r_Clock_Count[5]), 
            .I3(n17018), .O(\r_SM_Main_2__N_2031[1] ));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff80;
    SB_CARRY add_59_4 (.CI(n16133), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n16134));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n16132), .O(n312[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n10674));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_59_3 (.CI(n16132), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n16133));
    SB_LUT4 add_59_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n312[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n16132));
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n11144));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i11130210_i1_3_lut (.I0(n18235), .I1(n18085), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_2062));
    defparam i11130210_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_2062), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i5661_4_lut (.I0(\r_SM_Main_2__N_2034[0] ), .I1(n13614), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_2031[1] ), .O(n8191));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5661_4_lut.LUT_INIT = 16'hca0a;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n9269), .D(tx2_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n9269), .D(tx2_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n9269), .D(tx2_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n9269), .D(tx2_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n9269), .D(tx2_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n9269), .D(tx2_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n9269), .D(tx2_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_2034[0] ), .O(n9269));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i14635_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_2031[1] ), .O(n17412));
    defparam i14635_3_lut_4_lut.LUT_INIT = 16'heefe;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n11039));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx2_active), .C(CLK_c), .D(n11038));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx2_o), .C(CLK_c), .D(n11037));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n13614));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx2_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx2_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8458_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_2031[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n11144));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i8458_3_lut_4_lut_4_lut.LUT_INIT = 16'h0078;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (r_Bit_Index, n5244, GND_net, \r_SM_Main[1] , \r_SM_Main[2] , 
            n17361, CLK_c, n10983, rx_data_ready, n11019, n11031, 
            r_Rx_Data, rx_i, n11139, rx_data, n13744, n11136, n11135, 
            n1, n13116, n11112, n4, n11090, n11089, n18008, n11034, 
            n11026, VCC_net, n10987, n13692, n11018, n4_adj_1, n9999, 
            n17708, n17707, n4_adj_2, n10010) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [2:0]r_Bit_Index;
    output n5244;
    input GND_net;
    output \r_SM_Main[1] ;
    output \r_SM_Main[2] ;
    output n17361;
    input CLK_c;
    input n10983;
    output rx_data_ready;
    input n11019;
    input n11031;
    output r_Rx_Data;
    input rx_i;
    input n11139;
    output [7:0]rx_data;
    input n13744;
    input n11136;
    input n11135;
    output n1;
    output n13116;
    input n11112;
    output n4;
    input n11090;
    input n11089;
    output n18008;
    input n11034;
    input n11026;
    input VCC_net;
    input n10987;
    output n13692;
    output n11018;
    output n4_adj_1;
    output n9999;
    output n17708;
    output n17707;
    output n4_adj_2;
    output n10010;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]r_SM_Main_2__N_2088;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    wire [31:0]n194;
    
    wire n10656;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n10845, n16802, r_Rx_Data_R, n6, n17022, n17080;
    wire [2:0]r_SM_Main_2__N_2094;
    
    wire n6_adj_2130, n17636, n17380, n17635, n16131, n16130, n17058, 
        n16129, n16128, n16127, n16126, n16125, n10158, n10620;
    
    SB_LUT4 i2593_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5244));   // verilog/uart_rx.v(102[36:51])
    defparam i2593_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14585_4_lut (.I0(r_SM_Main_2__N_2088[2]), .I1(r_SM_Main[0]), 
            .I2(\r_SM_Main[1] ), .I3(\r_SM_Main[2] ), .O(n17361));
    defparam i14585_4_lut.LUT_INIT = 16'hffdc;
    SB_DFFESR r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n10656), 
            .D(n194[1]), .R(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n10656), 
            .D(n194[2]), .R(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n10656), 
            .D(n194[3]), .R(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n10656), 
            .D(n194[4]), .R(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n10656), 
            .D(n194[5]), .R(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n10656), 
            .D(n194[6]), .R(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n10656), 
            .D(n194[7]), .R(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n10656), 
            .D(n194[0]), .R(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n10983));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n16802));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .D(n11019));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .D(n11031));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(rx_i));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(n6), 
            .I3(r_Clock_Count[3]), .O(n17022));
    defparam i1_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(GND_net), .O(n17080));   // verilog/uart_rx.v(68[17:52])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_395 (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_2094[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2130));
    defparam i2_2_lut_adj_395.LUT_INIT = 16'h2222;
    SB_LUT4 i15081_4_lut (.I0(r_Clock_Count[5]), .I1(n17080), .I2(\r_SM_Main[2] ), 
            .I3(n17022), .O(n17636));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15081_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i15000_4_lut (.I0(n17080), .I1(r_SM_Main[0]), .I2(n17022), 
            .I3(n17380), .O(n17635));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15000_4_lut.LUT_INIT = 16'h3373;
    SB_LUT4 i1_4_lut_adj_396 (.I0(\r_SM_Main[2] ), .I1(n17635), .I2(n17636), 
            .I3(\r_SM_Main[1] ), .O(n10845));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut_adj_396.LUT_INIT = 16'h5044;
    SB_LUT4 i15215_4_lut (.I0(\r_SM_Main[2] ), .I1(\r_SM_Main[1] ), .I2(n6_adj_2130), 
            .I3(r_SM_Main[0]), .O(n10656));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i15215_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 add_62_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n16131), .O(n194[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_62_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n16130), .O(n194[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n11139));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(CLK_c), .D(n13744));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n11136));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n11135));   // verilog/uart_rx.v(49[10] 144[8])
    SB_CARRY add_62_8 (.CI(n16130), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n16131));
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_2094[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFFSR r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(CLK_c), .D(r_SM_Main_2__N_2088[2]), 
            .R(n17058));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i10445_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n13116));
    defparam i10445_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n11112));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_52_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_52_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n11090));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n11089));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i15231_1_lut (.I0(rx_data_ready), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18008));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15231_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_62_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n16129), .O(n194[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_7 (.CI(n16129), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n16130));
    SB_LUT4 add_62_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n16128), .O(n194[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14604_2_lut_3_lut (.I0(r_Clock_Count[5]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_2094[0]), 
            .I3(GND_net), .O(n17380));
    defparam i14604_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_CARRY add_62_6 (.CI(n16128), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n16129));
    SB_LUT4 add_62_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n16127), .O(n194[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_5 (.CI(n16127), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n16128));
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n11034));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n16126), .O(n194[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(n17022), .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_2094[0]));   // verilog/uart_rx.v(68[17:52])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n11026));   // verilog/uart_rx.v(49[10] 144[8])
    SB_CARRY add_62_4 (.CI(n16126), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n16127));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n16125), .O(n194[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_3 (.CI(n16125), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n16126));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n194[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n16125));
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n10987));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut (.I0(r_Bit_Index[2]), 
            .I1(n5244), .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_2088[2]), 
            .O(n13692));
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut.LUT_INIT = 16'hf70f;
    SB_LUT4 i14631_3_lut_4_lut (.I0(r_Bit_Index[2]), .I1(n5244), .I2(\r_SM_Main[1] ), 
            .I3(n17361), .O(n11018));
    defparam i14631_3_lut_4_lut.LUT_INIT = 16'hff70;
    SB_LUT4 equal_55_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_55_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_397 (.I0(r_Bit_Index[0]), .I1(n10158), .I2(GND_net), 
            .I3(GND_net), .O(n9999));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_397.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[6]), 
            .I2(r_Clock_Count[7]), .I3(n17022), .O(r_SM_Main_2__N_2088[2]));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i15089_2_lut (.I0(r_SM_Main_2__N_2088[2]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17708));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i15089_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15113_3_lut (.I0(r_SM_Main_2__N_2094[0]), .I1(r_SM_Main[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n17707));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i15113_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(\r_SM_Main[1] ), 
            .I3(r_SM_Main_2__N_2088[2]), .O(n10158));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 equal_56_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_56_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_398 (.I0(r_Bit_Index[0]), .I1(n10158), .I2(GND_net), 
            .I3(GND_net), .O(n10010));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_398.LUT_INIT = 16'hdddd;
    SB_LUT4 i15224_2_lut_3_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n17058));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i15224_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), .I2(r_SM_Main_2__N_2088[2]), 
            .I3(r_SM_Main[0]), .O(n10620));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), .I2(n10620), 
            .I3(rx_data_ready), .O(n16802));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    
endmodule
