// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Aug 26 2019 00:03:50

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    inout PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    input PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    inout PIN_1;
    output LED;
    input CLK;

    wire N__23697;
    wire N__23696;
    wire N__23695;
    wire N__23688;
    wire N__23687;
    wire N__23686;
    wire N__23679;
    wire N__23678;
    wire N__23677;
    wire N__23670;
    wire N__23669;
    wire N__23668;
    wire N__23661;
    wire N__23660;
    wire N__23659;
    wire N__23652;
    wire N__23651;
    wire N__23650;
    wire N__23633;
    wire N__23632;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23605;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23575;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23548;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23521;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23494;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23486;
    wire N__23485;
    wire N__23484;
    wire N__23483;
    wire N__23482;
    wire N__23481;
    wire N__23480;
    wire N__23479;
    wire N__23478;
    wire N__23477;
    wire N__23476;
    wire N__23475;
    wire N__23474;
    wire N__23473;
    wire N__23472;
    wire N__23471;
    wire N__23470;
    wire N__23469;
    wire N__23468;
    wire N__23467;
    wire N__23466;
    wire N__23465;
    wire N__23464;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23408;
    wire N__23405;
    wire N__23396;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23369;
    wire N__23360;
    wire N__23349;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23317;
    wire N__23316;
    wire N__23315;
    wire N__23314;
    wire N__23313;
    wire N__23310;
    wire N__23309;
    wire N__23308;
    wire N__23307;
    wire N__23306;
    wire N__23299;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23264;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23249;
    wire N__23246;
    wire N__23245;
    wire N__23244;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23226;
    wire N__23221;
    wire N__23218;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23206;
    wire N__23205;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23193;
    wire N__23190;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23162;
    wire N__23161;
    wire N__23160;
    wire N__23155;
    wire N__23150;
    wire N__23145;
    wire N__23142;
    wire N__23137;
    wire N__23130;
    wire N__23125;
    wire N__23114;
    wire N__23113;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23101;
    wire N__23100;
    wire N__23099;
    wire N__23098;
    wire N__23097;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23080;
    wire N__23079;
    wire N__23078;
    wire N__23073;
    wire N__23072;
    wire N__23071;
    wire N__23070;
    wire N__23069;
    wire N__23062;
    wire N__23057;
    wire N__23054;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23038;
    wire N__23035;
    wire N__23018;
    wire N__23015;
    wire N__23014;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23003;
    wire N__23002;
    wire N__23001;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22993;
    wire N__22992;
    wire N__22991;
    wire N__22988;
    wire N__22979;
    wire N__22974;
    wire N__22967;
    wire N__22958;
    wire N__22957;
    wire N__22956;
    wire N__22955;
    wire N__22954;
    wire N__22953;
    wire N__22952;
    wire N__22951;
    wire N__22950;
    wire N__22949;
    wire N__22948;
    wire N__22947;
    wire N__22946;
    wire N__22945;
    wire N__22944;
    wire N__22943;
    wire N__22942;
    wire N__22941;
    wire N__22940;
    wire N__22939;
    wire N__22938;
    wire N__22937;
    wire N__22936;
    wire N__22935;
    wire N__22934;
    wire N__22933;
    wire N__22932;
    wire N__22931;
    wire N__22930;
    wire N__22929;
    wire N__22928;
    wire N__22927;
    wire N__22926;
    wire N__22925;
    wire N__22924;
    wire N__22923;
    wire N__22922;
    wire N__22921;
    wire N__22920;
    wire N__22919;
    wire N__22918;
    wire N__22917;
    wire N__22916;
    wire N__22915;
    wire N__22914;
    wire N__22913;
    wire N__22912;
    wire N__22911;
    wire N__22910;
    wire N__22909;
    wire N__22908;
    wire N__22907;
    wire N__22906;
    wire N__22905;
    wire N__22904;
    wire N__22903;
    wire N__22902;
    wire N__22901;
    wire N__22900;
    wire N__22899;
    wire N__22898;
    wire N__22897;
    wire N__22896;
    wire N__22895;
    wire N__22894;
    wire N__22893;
    wire N__22892;
    wire N__22891;
    wire N__22890;
    wire N__22889;
    wire N__22888;
    wire N__22887;
    wire N__22886;
    wire N__22885;
    wire N__22884;
    wire N__22883;
    wire N__22882;
    wire N__22881;
    wire N__22880;
    wire N__22879;
    wire N__22878;
    wire N__22877;
    wire N__22876;
    wire N__22875;
    wire N__22874;
    wire N__22873;
    wire N__22872;
    wire N__22871;
    wire N__22870;
    wire N__22869;
    wire N__22868;
    wire N__22867;
    wire N__22866;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22651;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22624;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22594;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22529;
    wire N__22526;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22477;
    wire N__22472;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22460;
    wire N__22459;
    wire N__22458;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22446;
    wire N__22439;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22431;
    wire N__22428;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22401;
    wire N__22398;
    wire N__22391;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22330;
    wire N__22329;
    wire N__22326;
    wire N__22325;
    wire N__22324;
    wire N__22319;
    wire N__22316;
    wire N__22311;
    wire N__22308;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22266;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22254;
    wire N__22253;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22239;
    wire N__22232;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22188;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22166;
    wire N__22163;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22151;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22143;
    wire N__22142;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22127;
    wire N__22120;
    wire N__22117;
    wire N__22116;
    wire N__22115;
    wire N__22114;
    wire N__22109;
    wire N__22106;
    wire N__22101;
    wire N__22098;
    wire N__22093;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22067;
    wire N__22064;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22043;
    wire N__22042;
    wire N__22039;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22031;
    wire N__22028;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__22000;
    wire N__21997;
    wire N__21996;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21987;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21959;
    wire N__21958;
    wire N__21957;
    wire N__21956;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21940;
    wire N__21935;
    wire N__21932;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21890;
    wire N__21889;
    wire N__21886;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21872;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21854;
    wire N__21853;
    wire N__21852;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21829;
    wire N__21824;
    wire N__21823;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21815;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21788;
    wire N__21779;
    wire N__21776;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21768;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21740;
    wire N__21737;
    wire N__21736;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21728;
    wire N__21725;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21676;
    wire N__21673;
    wire N__21672;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21651;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21603;
    wire N__21602;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21584;
    wire N__21583;
    wire N__21580;
    wire N__21579;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21565;
    wire N__21564;
    wire N__21563;
    wire N__21562;
    wire N__21561;
    wire N__21560;
    wire N__21559;
    wire N__21556;
    wire N__21555;
    wire N__21554;
    wire N__21551;
    wire N__21546;
    wire N__21545;
    wire N__21544;
    wire N__21543;
    wire N__21542;
    wire N__21541;
    wire N__21540;
    wire N__21539;
    wire N__21538;
    wire N__21537;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21526;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21501;
    wire N__21490;
    wire N__21487;
    wire N__21486;
    wire N__21485;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21466;
    wire N__21465;
    wire N__21464;
    wire N__21463;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21449;
    wire N__21448;
    wire N__21447;
    wire N__21446;
    wire N__21445;
    wire N__21444;
    wire N__21443;
    wire N__21442;
    wire N__21441;
    wire N__21440;
    wire N__21439;
    wire N__21438;
    wire N__21437;
    wire N__21436;
    wire N__21435;
    wire N__21434;
    wire N__21433;
    wire N__21430;
    wire N__21421;
    wire N__21414;
    wire N__21411;
    wire N__21406;
    wire N__21403;
    wire N__21398;
    wire N__21389;
    wire N__21384;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21338;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21307;
    wire N__21302;
    wire N__21289;
    wire N__21260;
    wire N__21259;
    wire N__21258;
    wire N__21257;
    wire N__21256;
    wire N__21255;
    wire N__21252;
    wire N__21251;
    wire N__21250;
    wire N__21249;
    wire N__21248;
    wire N__21247;
    wire N__21246;
    wire N__21243;
    wire N__21242;
    wire N__21239;
    wire N__21238;
    wire N__21235;
    wire N__21234;
    wire N__21229;
    wire N__21226;
    wire N__21221;
    wire N__21220;
    wire N__21219;
    wire N__21216;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21186;
    wire N__21185;
    wire N__21184;
    wire N__21183;
    wire N__21182;
    wire N__21181;
    wire N__21180;
    wire N__21179;
    wire N__21178;
    wire N__21177;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21162;
    wire N__21159;
    wire N__21154;
    wire N__21153;
    wire N__21152;
    wire N__21151;
    wire N__21150;
    wire N__21149;
    wire N__21148;
    wire N__21147;
    wire N__21146;
    wire N__21145;
    wire N__21144;
    wire N__21143;
    wire N__21142;
    wire N__21141;
    wire N__21140;
    wire N__21139;
    wire N__21138;
    wire N__21137;
    wire N__21136;
    wire N__21135;
    wire N__21134;
    wire N__21133;
    wire N__21132;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21114;
    wire N__21109;
    wire N__21098;
    wire N__21093;
    wire N__21084;
    wire N__21075;
    wire N__21070;
    wire N__21059;
    wire N__21048;
    wire N__21041;
    wire N__21032;
    wire N__21019;
    wire N__20990;
    wire N__20989;
    wire N__20986;
    wire N__20985;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20954;
    wire N__20951;
    wire N__20950;
    wire N__20947;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20923;
    wire N__20922;
    wire N__20917;
    wire N__20914;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20891;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20883;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20865;
    wire N__20858;
    wire N__20857;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20849;
    wire N__20846;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20825;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20807;
    wire N__20806;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20792;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20764;
    wire N__20761;
    wire N__20760;
    wire N__20759;
    wire N__20756;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20742;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20707;
    wire N__20706;
    wire N__20705;
    wire N__20702;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20694;
    wire N__20693;
    wire N__20690;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20682;
    wire N__20681;
    wire N__20680;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20660;
    wire N__20655;
    wire N__20650;
    wire N__20645;
    wire N__20644;
    wire N__20643;
    wire N__20640;
    wire N__20633;
    wire N__20628;
    wire N__20625;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20594;
    wire N__20591;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20583;
    wire N__20580;
    wire N__20579;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20564;
    wire N__20555;
    wire N__20554;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20550;
    wire N__20549;
    wire N__20548;
    wire N__20547;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20535;
    wire N__20532;
    wire N__20527;
    wire N__20520;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20513;
    wire N__20502;
    wire N__20497;
    wire N__20496;
    wire N__20495;
    wire N__20494;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20480;
    wire N__20479;
    wire N__20478;
    wire N__20477;
    wire N__20472;
    wire N__20467;
    wire N__20466;
    wire N__20465;
    wire N__20462;
    wire N__20457;
    wire N__20454;
    wire N__20453;
    wire N__20452;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20438;
    wire N__20433;
    wire N__20430;
    wire N__20425;
    wire N__20424;
    wire N__20423;
    wire N__20420;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20404;
    wire N__20401;
    wire N__20394;
    wire N__20389;
    wire N__20386;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20359;
    wire N__20358;
    wire N__20355;
    wire N__20350;
    wire N__20345;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20328;
    wire N__20327;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20288;
    wire N__20285;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20264;
    wire N__20263;
    wire N__20262;
    wire N__20259;
    wire N__20258;
    wire N__20257;
    wire N__20252;
    wire N__20247;
    wire N__20244;
    wire N__20237;
    wire N__20236;
    wire N__20235;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20198;
    wire N__20195;
    wire N__20194;
    wire N__20193;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20174;
    wire N__20171;
    wire N__20162;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20151;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20139;
    wire N__20136;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20096;
    wire N__20093;
    wire N__20092;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20074;
    wire N__20071;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20063;
    wire N__20062;
    wire N__20061;
    wire N__20060;
    wire N__20059;
    wire N__20058;
    wire N__20057;
    wire N__20056;
    wire N__20055;
    wire N__20054;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20030;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20014;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19984;
    wire N__19983;
    wire N__19982;
    wire N__19979;
    wire N__19972;
    wire N__19967;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19955;
    wire N__19954;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19946;
    wire N__19945;
    wire N__19940;
    wire N__19935;
    wire N__19932;
    wire N__19927;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19904;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19889;
    wire N__19886;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19878;
    wire N__19877;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19854;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19826;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19818;
    wire N__19817;
    wire N__19814;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19768;
    wire N__19767;
    wire N__19764;
    wire N__19759;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19685;
    wire N__19684;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19657;
    wire N__19656;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19644;
    wire N__19637;
    wire N__19634;
    wire N__19633;
    wire N__19632;
    wire N__19629;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19607;
    wire N__19604;
    wire N__19603;
    wire N__19602;
    wire N__19601;
    wire N__19598;
    wire N__19597;
    wire N__19596;
    wire N__19591;
    wire N__19590;
    wire N__19589;
    wire N__19586;
    wire N__19585;
    wire N__19582;
    wire N__19577;
    wire N__19574;
    wire N__19569;
    wire N__19568;
    wire N__19567;
    wire N__19566;
    wire N__19565;
    wire N__19562;
    wire N__19561;
    wire N__19558;
    wire N__19549;
    wire N__19546;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19522;
    wire N__19517;
    wire N__19512;
    wire N__19505;
    wire N__19502;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19286;
    wire N__19285;
    wire N__19282;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19270;
    wire N__19265;
    wire N__19262;
    wire N__19261;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19242;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19228;
    wire N__19227;
    wire N__19226;
    wire N__19223;
    wire N__19216;
    wire N__19211;
    wire N__19210;
    wire N__19209;
    wire N__19208;
    wire N__19207;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19199;
    wire N__19194;
    wire N__19189;
    wire N__19186;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19172;
    wire N__19169;
    wire N__19160;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19132;
    wire N__19127;
    wire N__19122;
    wire N__19119;
    wire N__19112;
    wire N__19111;
    wire N__19110;
    wire N__19107;
    wire N__19106;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19091;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18967;
    wire N__18966;
    wire N__18965;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18905;
    wire N__18902;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18894;
    wire N__18889;
    wire N__18888;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18764;
    wire N__18761;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18749;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18734;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18722;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18710;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18698;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18683;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18585;
    wire N__18584;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18563;
    wire N__18562;
    wire N__18559;
    wire N__18558;
    wire N__18557;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18533;
    wire N__18530;
    wire N__18523;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18511;
    wire N__18510;
    wire N__18509;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18486;
    wire N__18479;
    wire N__18476;
    wire N__18475;
    wire N__18472;
    wire N__18471;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18459;
    wire N__18452;
    wire N__18451;
    wire N__18450;
    wire N__18447;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18432;
    wire N__18427;
    wire N__18424;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18365;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18357;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18337;
    wire N__18332;
    wire N__18329;
    wire N__18328;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18315;
    wire N__18314;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18266;
    wire N__18265;
    wire N__18262;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18215;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18173;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18088;
    wire N__18085;
    wire N__18082;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18067;
    wire N__18064;
    wire N__18061;
    wire N__18056;
    wire N__18055;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17981;
    wire N__17978;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17932;
    wire N__17931;
    wire N__17930;
    wire N__17929;
    wire N__17926;
    wire N__17925;
    wire N__17924;
    wire N__17921;
    wire N__17914;
    wire N__17907;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17890;
    wire N__17889;
    wire N__17888;
    wire N__17887;
    wire N__17886;
    wire N__17883;
    wire N__17880;
    wire N__17875;
    wire N__17870;
    wire N__17861;
    wire N__17858;
    wire N__17857;
    wire N__17856;
    wire N__17855;
    wire N__17852;
    wire N__17847;
    wire N__17846;
    wire N__17843;
    wire N__17838;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17809;
    wire N__17808;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17796;
    wire N__17789;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17781;
    wire N__17780;
    wire N__17779;
    wire N__17778;
    wire N__17773;
    wire N__17768;
    wire N__17767;
    wire N__17766;
    wire N__17763;
    wire N__17762;
    wire N__17761;
    wire N__17760;
    wire N__17757;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17745;
    wire N__17736;
    wire N__17733;
    wire N__17730;
    wire N__17727;
    wire N__17720;
    wire N__17711;
    wire N__17710;
    wire N__17709;
    wire N__17708;
    wire N__17707;
    wire N__17706;
    wire N__17705;
    wire N__17702;
    wire N__17697;
    wire N__17688;
    wire N__17687;
    wire N__17686;
    wire N__17685;
    wire N__17684;
    wire N__17683;
    wire N__17680;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17655;
    wire N__17646;
    wire N__17639;
    wire N__17638;
    wire N__17637;
    wire N__17634;
    wire N__17633;
    wire N__17632;
    wire N__17631;
    wire N__17630;
    wire N__17629;
    wire N__17628;
    wire N__17627;
    wire N__17622;
    wire N__17621;
    wire N__17620;
    wire N__17619;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17607;
    wire N__17598;
    wire N__17595;
    wire N__17588;
    wire N__17585;
    wire N__17576;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17557;
    wire N__17556;
    wire N__17555;
    wire N__17554;
    wire N__17553;
    wire N__17552;
    wire N__17551;
    wire N__17550;
    wire N__17545;
    wire N__17544;
    wire N__17543;
    wire N__17542;
    wire N__17537;
    wire N__17528;
    wire N__17525;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17517;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17499;
    wire N__17496;
    wire N__17489;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17451;
    wire N__17446;
    wire N__17443;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17419;
    wire N__17418;
    wire N__17417;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17396;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17374;
    wire N__17373;
    wire N__17372;
    wire N__17369;
    wire N__17368;
    wire N__17367;
    wire N__17364;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17276;
    wire N__17273;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17265;
    wire N__17262;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17242;
    wire N__17237;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17222;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17207;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17192;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17129;
    wire N__17128;
    wire N__17127;
    wire N__17126;
    wire N__17121;
    wire N__17120;
    wire N__17117;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17103;
    wire N__17102;
    wire N__17101;
    wire N__17100;
    wire N__17099;
    wire N__17098;
    wire N__17097;
    wire N__17096;
    wire N__17095;
    wire N__17094;
    wire N__17093;
    wire N__17092;
    wire N__17091;
    wire N__17090;
    wire N__17089;
    wire N__17088;
    wire N__17087;
    wire N__17080;
    wire N__17075;
    wire N__17070;
    wire N__17069;
    wire N__17066;
    wire N__17065;
    wire N__17064;
    wire N__17063;
    wire N__17062;
    wire N__17061;
    wire N__17060;
    wire N__17059;
    wire N__17058;
    wire N__17057;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17049;
    wire N__17046;
    wire N__17041;
    wire N__17038;
    wire N__17033;
    wire N__17028;
    wire N__17025;
    wire N__17024;
    wire N__17023;
    wire N__17022;
    wire N__17021;
    wire N__17020;
    wire N__17019;
    wire N__17012;
    wire N__17003;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16999;
    wire N__16998;
    wire N__16997;
    wire N__16996;
    wire N__16989;
    wire N__16988;
    wire N__16987;
    wire N__16986;
    wire N__16985;
    wire N__16974;
    wire N__16973;
    wire N__16972;
    wire N__16971;
    wire N__16970;
    wire N__16965;
    wire N__16962;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16932;
    wire N__16929;
    wire N__16924;
    wire N__16923;
    wire N__16922;
    wire N__16921;
    wire N__16920;
    wire N__16919;
    wire N__16918;
    wire N__16917;
    wire N__16908;
    wire N__16907;
    wire N__16906;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16893;
    wire N__16884;
    wire N__16881;
    wire N__16874;
    wire N__16871;
    wire N__16866;
    wire N__16863;
    wire N__16856;
    wire N__16843;
    wire N__16832;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16816;
    wire N__16811;
    wire N__16806;
    wire N__16801;
    wire N__16790;
    wire N__16787;
    wire N__16780;
    wire N__16763;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16752;
    wire N__16751;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16676;
    wire N__16675;
    wire N__16672;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16657;
    wire N__16654;
    wire N__16651;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16639;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16591;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16579;
    wire N__16578;
    wire N__16577;
    wire N__16572;
    wire N__16567;
    wire N__16562;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16474;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16464;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16429;
    wire N__16428;
    wire N__16425;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16396;
    wire N__16395;
    wire N__16394;
    wire N__16393;
    wire N__16392;
    wire N__16391;
    wire N__16388;
    wire N__16383;
    wire N__16378;
    wire N__16373;
    wire N__16364;
    wire N__16363;
    wire N__16362;
    wire N__16361;
    wire N__16360;
    wire N__16359;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16344;
    wire N__16339;
    wire N__16328;
    wire N__16327;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16306;
    wire N__16305;
    wire N__16304;
    wire N__16301;
    wire N__16298;
    wire N__16293;
    wire N__16290;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16273;
    wire N__16272;
    wire N__16271;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16256;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16225;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16180;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16170;
    wire N__16163;
    wire N__16162;
    wire N__16159;
    wire N__16158;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16144;
    wire N__16143;
    wire N__16136;
    wire N__16133;
    wire N__16132;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16088;
    wire N__16087;
    wire N__16086;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16033;
    wire N__16032;
    wire N__16031;
    wire N__16028;
    wire N__16027;
    wire N__16026;
    wire N__16021;
    wire N__16016;
    wire N__16011;
    wire N__16004;
    wire N__16001;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15902;
    wire N__15899;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15887;
    wire N__15884;
    wire N__15883;
    wire N__15882;
    wire N__15879;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15854;
    wire N__15853;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15825;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15787;
    wire N__15786;
    wire N__15785;
    wire N__15784;
    wire N__15783;
    wire N__15782;
    wire N__15779;
    wire N__15778;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15767;
    wire N__15766;
    wire N__15765;
    wire N__15762;
    wire N__15761;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15747;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15735;
    wire N__15732;
    wire N__15731;
    wire N__15728;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15714;
    wire N__15711;
    wire N__15706;
    wire N__15705;
    wire N__15698;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15672;
    wire N__15669;
    wire N__15664;
    wire N__15661;
    wire N__15656;
    wire N__15647;
    wire N__15646;
    wire N__15641;
    wire N__15640;
    wire N__15639;
    wire N__15638;
    wire N__15637;
    wire N__15636;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15609;
    wire N__15608;
    wire N__15605;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15571;
    wire N__15560;
    wire N__15559;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15548;
    wire N__15547;
    wire N__15546;
    wire N__15545;
    wire N__15544;
    wire N__15537;
    wire N__15532;
    wire N__15529;
    wire N__15528;
    wire N__15527;
    wire N__15526;
    wire N__15525;
    wire N__15522;
    wire N__15521;
    wire N__15520;
    wire N__15519;
    wire N__15518;
    wire N__15517;
    wire N__15516;
    wire N__15515;
    wire N__15514;
    wire N__15513;
    wire N__15512;
    wire N__15511;
    wire N__15510;
    wire N__15507;
    wire N__15502;
    wire N__15499;
    wire N__15496;
    wire N__15495;
    wire N__15492;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15471;
    wire N__15470;
    wire N__15469;
    wire N__15468;
    wire N__15467;
    wire N__15466;
    wire N__15461;
    wire N__15454;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15436;
    wire N__15433;
    wire N__15432;
    wire N__15431;
    wire N__15430;
    wire N__15427;
    wire N__15418;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15402;
    wire N__15397;
    wire N__15390;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15364;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15332;
    wire N__15329;
    wire N__15328;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15310;
    wire N__15305;
    wire N__15302;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15229;
    wire N__15228;
    wire N__15227;
    wire N__15226;
    wire N__15225;
    wire N__15224;
    wire N__15223;
    wire N__15222;
    wire N__15219;
    wire N__15208;
    wire N__15201;
    wire N__15194;
    wire N__15193;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15183;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15143;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15131;
    wire N__15128;
    wire N__15127;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15106;
    wire N__15105;
    wire N__15102;
    wire N__15097;
    wire N__15092;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15079;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15047;
    wire N__15046;
    wire N__15045;
    wire N__15044;
    wire N__15043;
    wire N__15042;
    wire N__15039;
    wire N__15038;
    wire N__15037;
    wire N__15036;
    wire N__15035;
    wire N__15034;
    wire N__15033;
    wire N__15032;
    wire N__15031;
    wire N__15030;
    wire N__15029;
    wire N__15028;
    wire N__15027;
    wire N__15026;
    wire N__15025;
    wire N__15024;
    wire N__15023;
    wire N__15022;
    wire N__15021;
    wire N__15020;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15016;
    wire N__15015;
    wire N__15014;
    wire N__15013;
    wire N__15012;
    wire N__15011;
    wire N__15010;
    wire N__15009;
    wire N__15006;
    wire N__15001;
    wire N__14998;
    wire N__14997;
    wire N__14994;
    wire N__14989;
    wire N__14984;
    wire N__14979;
    wire N__14978;
    wire N__14977;
    wire N__14974;
    wire N__14965;
    wire N__14964;
    wire N__14963;
    wire N__14962;
    wire N__14961;
    wire N__14960;
    wire N__14959;
    wire N__14958;
    wire N__14957;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14946;
    wire N__14945;
    wire N__14944;
    wire N__14941;
    wire N__14940;
    wire N__14939;
    wire N__14938;
    wire N__14937;
    wire N__14936;
    wire N__14935;
    wire N__14934;
    wire N__14933;
    wire N__14932;
    wire N__14931;
    wire N__14930;
    wire N__14929;
    wire N__14928;
    wire N__14919;
    wire N__14914;
    wire N__14901;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14881;
    wire N__14872;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14839;
    wire N__14836;
    wire N__14831;
    wire N__14826;
    wire N__14823;
    wire N__14818;
    wire N__14811;
    wire N__14804;
    wire N__14791;
    wire N__14786;
    wire N__14777;
    wire N__14772;
    wire N__14765;
    wire N__14762;
    wire N__14751;
    wire N__14726;
    wire N__14725;
    wire N__14724;
    wire N__14723;
    wire N__14722;
    wire N__14721;
    wire N__14720;
    wire N__14717;
    wire N__14716;
    wire N__14715;
    wire N__14714;
    wire N__14713;
    wire N__14712;
    wire N__14711;
    wire N__14708;
    wire N__14707;
    wire N__14706;
    wire N__14705;
    wire N__14704;
    wire N__14703;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14695;
    wire N__14694;
    wire N__14693;
    wire N__14690;
    wire N__14689;
    wire N__14688;
    wire N__14687;
    wire N__14686;
    wire N__14685;
    wire N__14684;
    wire N__14681;
    wire N__14674;
    wire N__14671;
    wire N__14670;
    wire N__14669;
    wire N__14666;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14655;
    wire N__14654;
    wire N__14653;
    wire N__14652;
    wire N__14647;
    wire N__14646;
    wire N__14645;
    wire N__14644;
    wire N__14643;
    wire N__14642;
    wire N__14641;
    wire N__14640;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14629;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14621;
    wire N__14612;
    wire N__14607;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14591;
    wire N__14590;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14579;
    wire N__14578;
    wire N__14575;
    wire N__14574;
    wire N__14571;
    wire N__14570;
    wire N__14567;
    wire N__14562;
    wire N__14555;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14531;
    wire N__14518;
    wire N__14509;
    wire N__14502;
    wire N__14501;
    wire N__14496;
    wire N__14495;
    wire N__14494;
    wire N__14493;
    wire N__14490;
    wire N__14487;
    wire N__14486;
    wire N__14485;
    wire N__14484;
    wire N__14481;
    wire N__14474;
    wire N__14473;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14465;
    wire N__14464;
    wire N__14459;
    wire N__14454;
    wire N__14451;
    wire N__14432;
    wire N__14429;
    wire N__14428;
    wire N__14425;
    wire N__14420;
    wire N__14407;
    wire N__14406;
    wire N__14405;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14389;
    wire N__14384;
    wire N__14381;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14367;
    wire N__14362;
    wire N__14359;
    wire N__14354;
    wire N__14351;
    wire N__14346;
    wire N__14337;
    wire N__14334;
    wire N__14315;
    wire N__14312;
    wire N__14311;
    wire N__14310;
    wire N__14307;
    wire N__14304;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14288;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14276;
    wire N__14273;
    wire N__14272;
    wire N__14271;
    wire N__14268;
    wire N__14265;
    wire N__14262;
    wire N__14255;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14247;
    wire N__14242;
    wire N__14239;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14227;
    wire N__14226;
    wire N__14223;
    wire N__14220;
    wire N__14217;
    wire N__14210;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14202;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14182;
    wire N__14177;
    wire N__14174;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14162;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14150;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14142;
    wire N__14139;
    wire N__14134;
    wire N__14129;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14118;
    wire N__14115;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14090;
    wire N__14087;
    wire N__14086;
    wire N__14085;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14060;
    wire N__14057;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14014;
    wire N__14013;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13976;
    wire N__13973;
    wire N__13972;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13964;
    wire N__13963;
    wire N__13960;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13940;
    wire N__13939;
    wire N__13936;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13914;
    wire N__13907;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13897;
    wire N__13896;
    wire N__13895;
    wire N__13890;
    wire N__13887;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13835;
    wire N__13832;
    wire N__13831;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13821;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13796;
    wire N__13793;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13785;
    wire N__13784;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13763;
    wire N__13760;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13752;
    wire N__13751;
    wire N__13746;
    wire N__13743;
    wire N__13742;
    wire N__13739;
    wire N__13734;
    wire N__13731;
    wire N__13724;
    wire N__13723;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13692;
    wire N__13685;
    wire N__13682;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13674;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13645;
    wire N__13644;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13636;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13613;
    wire N__13612;
    wire N__13609;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13598;
    wire N__13597;
    wire N__13594;
    wire N__13591;
    wire N__13588;
    wire N__13585;
    wire N__13582;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13558;
    wire N__13555;
    wire N__13554;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13542;
    wire N__13535;
    wire N__13532;
    wire N__13531;
    wire N__13530;
    wire N__13527;
    wire N__13526;
    wire N__13525;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13499;
    wire N__13496;
    wire N__13495;
    wire N__13492;
    wire N__13489;
    wire N__13486;
    wire N__13485;
    wire N__13482;
    wire N__13481;
    wire N__13480;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13466;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13447;
    wire N__13444;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13433;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13417;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13369;
    wire N__13368;
    wire N__13367;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13357;
    wire N__13352;
    wire N__13343;
    wire N__13342;
    wire N__13341;
    wire N__13338;
    wire N__13335;
    wire N__13332;
    wire N__13329;
    wire N__13328;
    wire N__13327;
    wire N__13324;
    wire N__13321;
    wire N__13318;
    wire N__13313;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13297;
    wire N__13294;
    wire N__13293;
    wire N__13290;
    wire N__13285;
    wire N__13284;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13272;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13260;
    wire N__13257;
    wire N__13254;
    wire N__13251;
    wire N__13250;
    wire N__13249;
    wire N__13242;
    wire N__13237;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13222;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13193;
    wire N__13190;
    wire N__13189;
    wire N__13186;
    wire N__13185;
    wire N__13184;
    wire N__13183;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13151;
    wire N__13148;
    wire N__13147;
    wire N__13146;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13121;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13099;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13091;
    wire N__13086;
    wire N__13081;
    wire N__13076;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13046;
    wire N__13045;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13031;
    wire N__13028;
    wire N__13023;
    wire N__13022;
    wire N__13019;
    wire N__13014;
    wire N__13011;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12965;
    wire N__12962;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12895;
    wire N__12892;
    wire N__12889;
    wire N__12886;
    wire N__12883;
    wire N__12878;
    wire N__12877;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12835;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12814;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12794;
    wire N__12791;
    wire N__12790;
    wire N__12787;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12724;
    wire N__12723;
    wire N__12720;
    wire N__12715;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12694;
    wire N__12693;
    wire N__12692;
    wire N__12689;
    wire N__12688;
    wire N__12685;
    wire N__12680;
    wire N__12677;
    wire N__12672;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12649;
    wire N__12648;
    wire N__12645;
    wire N__12644;
    wire N__12641;
    wire N__12640;
    wire N__12639;
    wire N__12638;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12624;
    wire N__12623;
    wire N__12620;
    wire N__12619;
    wire N__12616;
    wire N__12609;
    wire N__12604;
    wire N__12601;
    wire N__12600;
    wire N__12595;
    wire N__12592;
    wire N__12587;
    wire N__12584;
    wire N__12579;
    wire N__12572;
    wire N__12571;
    wire N__12570;
    wire N__12569;
    wire N__12566;
    wire N__12565;
    wire N__12562;
    wire N__12561;
    wire N__12560;
    wire N__12559;
    wire N__12558;
    wire N__12555;
    wire N__12554;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12534;
    wire N__12529;
    wire N__12528;
    wire N__12525;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12504;
    wire N__12501;
    wire N__12494;
    wire N__12489;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12463;
    wire N__12462;
    wire N__12461;
    wire N__12460;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12450;
    wire N__12449;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12414;
    wire N__12413;
    wire N__12412;
    wire N__12411;
    wire N__12410;
    wire N__12409;
    wire N__12408;
    wire N__12407;
    wire N__12398;
    wire N__12389;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12371;
    wire N__12368;
    wire N__12361;
    wire N__12356;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12323;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12310;
    wire N__12309;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12291;
    wire N__12284;
    wire N__12283;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12273;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12202;
    wire N__12199;
    wire N__12196;
    wire N__12191;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12164;
    wire N__12163;
    wire N__12160;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12143;
    wire N__12140;
    wire N__12139;
    wire N__12138;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12113;
    wire N__12112;
    wire N__12109;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12084;
    wire N__12077;
    wire N__12074;
    wire N__12073;
    wire N__12068;
    wire N__12065;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12047;
    wire N__12046;
    wire N__12043;
    wire N__12042;
    wire N__12039;
    wire N__12038;
    wire N__12037;
    wire N__12034;
    wire N__12031;
    wire N__12028;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12008;
    wire N__12007;
    wire N__12004;
    wire N__12003;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11991;
    wire N__11984;
    wire N__11983;
    wire N__11980;
    wire N__11979;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11948;
    wire N__11945;
    wire N__11944;
    wire N__11943;
    wire N__11940;
    wire N__11935;
    wire N__11932;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11917;
    wire N__11914;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11902;
    wire N__11897;
    wire N__11896;
    wire N__11893;
    wire N__11892;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11870;
    wire N__11867;
    wire N__11866;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11839;
    wire N__11838;
    wire N__11835;
    wire N__11834;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11806;
    wire N__11805;
    wire N__11802;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11761;
    wire N__11758;
    wire N__11757;
    wire N__11756;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11716;
    wire N__11715;
    wire N__11712;
    wire N__11707;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11685;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11673;
    wire N__11666;
    wire N__11663;
    wire N__11662;
    wire N__11661;
    wire N__11658;
    wire N__11655;
    wire N__11654;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11636;
    wire N__11635;
    wire N__11632;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11603;
    wire N__11602;
    wire N__11597;
    wire N__11596;
    wire N__11593;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11498;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11487;
    wire N__11482;
    wire N__11479;
    wire N__11474;
    wire N__11471;
    wire N__11470;
    wire N__11469;
    wire N__11466;
    wire N__11461;
    wire N__11458;
    wire N__11453;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11440;
    wire N__11439;
    wire N__11436;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11421;
    wire N__11414;
    wire N__11413;
    wire N__11412;
    wire N__11411;
    wire N__11404;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11387;
    wire N__11384;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11357;
    wire N__11356;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11339;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11248;
    wire N__11247;
    wire N__11246;
    wire N__11243;
    wire N__11236;
    wire N__11231;
    wire N__11230;
    wire N__11229;
    wire N__11228;
    wire N__11227;
    wire N__11224;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11204;
    wire N__11201;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11134;
    wire N__11129;
    wire N__11126;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11114;
    wire N__11113;
    wire N__11108;
    wire N__11105;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11093;
    wire N__11090;
    wire N__11089;
    wire N__11084;
    wire N__11081;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11069;
    wire N__11068;
    wire N__11065;
    wire N__11060;
    wire N__11057;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11000;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10989;
    wire N__10988;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10976;
    wire N__10973;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10934;
    wire N__10933;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10916;
    wire N__10915;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10898;
    wire N__10897;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10887;
    wire N__10884;
    wire N__10877;
    wire N__10876;
    wire N__10875;
    wire N__10872;
    wire N__10869;
    wire N__10866;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10849;
    wire N__10848;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10822;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10805;
    wire N__10802;
    wire N__10801;
    wire N__10800;
    wire N__10799;
    wire N__10798;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10788;
    wire N__10785;
    wire N__10780;
    wire N__10769;
    wire N__10768;
    wire N__10767;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10755;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10699;
    wire N__10696;
    wire N__10693;
    wire N__10690;
    wire N__10685;
    wire N__10684;
    wire N__10681;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10654;
    wire N__10653;
    wire N__10650;
    wire N__10645;
    wire N__10640;
    wire N__10637;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10625;
    wire N__10622;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10603;
    wire N__10602;
    wire N__10599;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10556;
    wire N__10553;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10500;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10478;
    wire N__10475;
    wire N__10474;
    wire N__10471;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10454;
    wire N__10451;
    wire N__10450;
    wire N__10447;
    wire N__10446;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10424;
    wire N__10423;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10375;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10358;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10346;
    wire N__10343;
    wire N__10342;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10331;
    wire N__10330;
    wire N__10323;
    wire N__10318;
    wire N__10313;
    wire N__10310;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10302;
    wire N__10301;
    wire N__10296;
    wire N__10295;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10272;
    wire N__10267;
    wire N__10266;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10198;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10174;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10163;
    wire N__10160;
    wire N__10155;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10133;
    wire N__10132;
    wire N__10131;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10120;
    wire N__10119;
    wire N__10116;
    wire N__10113;
    wire N__10108;
    wire N__10105;
    wire N__10100;
    wire N__10091;
    wire N__10088;
    wire N__10087;
    wire N__10086;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10066;
    wire N__10061;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10053;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10041;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10021;
    wire N__10020;
    wire N__10019;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9943;
    wire N__9942;
    wire N__9939;
    wire N__9934;
    wire N__9929;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9921;
    wire N__9920;
    wire N__9919;
    wire N__9914;
    wire N__9909;
    wire N__9906;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9866;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9854;
    wire N__9851;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9829;
    wire N__9828;
    wire N__9827;
    wire N__9824;
    wire N__9819;
    wire N__9816;
    wire N__9809;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9801;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9776;
    wire N__9773;
    wire N__9772;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9764;
    wire N__9761;
    wire N__9756;
    wire N__9751;
    wire N__9746;
    wire N__9743;
    wire N__9742;
    wire N__9741;
    wire N__9738;
    wire N__9733;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9697;
    wire N__9696;
    wire N__9693;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9637;
    wire N__9634;
    wire N__9633;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9613;
    wire N__9612;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9580;
    wire N__9579;
    wire N__9576;
    wire N__9575;
    wire N__9574;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9551;
    wire N__9550;
    wire N__9549;
    wire N__9548;
    wire N__9545;
    wire N__9544;
    wire N__9543;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9528;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9506;
    wire N__9505;
    wire N__9502;
    wire N__9501;
    wire N__9500;
    wire N__9499;
    wire N__9498;
    wire N__9495;
    wire N__9492;
    wire N__9491;
    wire N__9490;
    wire N__9485;
    wire N__9480;
    wire N__9475;
    wire N__9470;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9409;
    wire N__9408;
    wire N__9405;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9367;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9345;
    wire N__9338;
    wire N__9337;
    wire N__9336;
    wire N__9333;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9310;
    wire N__9305;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9290;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9273;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9261;
    wire N__9254;
    wire N__9251;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9219;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9181;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9131;
    wire N__9130;
    wire N__9129;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9107;
    wire N__9104;
    wire N__9103;
    wire N__9100;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9083;
    wire N__9082;
    wire N__9079;
    wire N__9078;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9066;
    wire N__9063;
    wire N__9056;
    wire N__9055;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8977;
    wire N__8974;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8957;
    wire N__8956;
    wire N__8953;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8945;
    wire N__8942;
    wire N__8937;
    wire N__8934;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8920;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8899;
    wire N__8894;
    wire N__8891;
    wire N__8890;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8857;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8843;
    wire N__8840;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8825;
    wire N__8822;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8797;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8767;
    wire N__8762;
    wire N__8759;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8714;
    wire N__8713;
    wire N__8712;
    wire N__8709;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8671;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8653;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire n26;
    wire bfn_1_22_0_;
    wire n25;
    wire n3851;
    wire n24;
    wire n3852;
    wire n23;
    wire n3853;
    wire n22;
    wire n3854;
    wire n21;
    wire n3855;
    wire n20;
    wire n3856;
    wire n19;
    wire n3857;
    wire n3858;
    wire n18;
    wire bfn_1_23_0_;
    wire n17;
    wire n3859;
    wire n16;
    wire n3860;
    wire n15;
    wire n3861;
    wire n14;
    wire n3862;
    wire n13;
    wire n3863;
    wire n12;
    wire n3864;
    wire n11;
    wire n3865;
    wire n3866;
    wire n10;
    wire bfn_1_24_0_;
    wire n9;
    wire n3867;
    wire n8;
    wire n3868;
    wire n7;
    wire n3869;
    wire n6;
    wire n3870;
    wire n3871;
    wire n3872;
    wire n3873;
    wire n3874;
    wire bfn_1_25_0_;
    wire n3875;
    wire \c0.n4849_cascade_ ;
    wire \c0.n4568 ;
    wire \c0.n4582 ;
    wire \c0.n4591_cascade_ ;
    wire \c0.n28_cascade_ ;
    wire \c0.n22 ;
    wire \c0.data_in_frame_6_6 ;
    wire \c0.n4592 ;
    wire \c0.n25_cascade_ ;
    wire data_in_1_5;
    wire \c0.n28_adj_868 ;
    wire \c0.n26 ;
    wire \c0.data_in_frame_7_3 ;
    wire \c0.n4601 ;
    wire \c0.data_in_frame_6_3 ;
    wire \c0.data_in_frame_7_6 ;
    wire \c0.n4831 ;
    wire tx2_data_6_keep_cascade_;
    wire r_Tx_Data_6_adj_958;
    wire \c0.data_in_frame_6_4 ;
    wire \c0.data_in_frame_7_2 ;
    wire \c0.n4604_cascade_ ;
    wire \c0.data_in_frame_6_7 ;
    wire \c0.n4583 ;
    wire \c0.data_in_frame_7_7 ;
    wire \c0.data_in_frame_7_4 ;
    wire \c0.n4555 ;
    wire tx2_data_7_keep;
    wire r_Tx_Data_5_adj_959;
    wire n4624;
    wire \c0.n4801_cascade_ ;
    wire tx2_data_1_keep_cascade_;
    wire r_Tx_Data_1_adj_963;
    wire r_Tx_Data_7_adj_957;
    wire n4625;
    wire \c0.n4540 ;
    wire \c0.n4606 ;
    wire \c0.n4552 ;
    wire \c0.n4553_cascade_ ;
    wire tx2_data_5_keep;
    wire data_in_0_5;
    wire data_in_1_0;
    wire data_in_5_6;
    wire \c0.n4594 ;
    wire \c0.n4825 ;
    wire \c0.n4813 ;
    wire tx2_data_3_keep_cascade_;
    wire r_Tx_Data_3_adj_961;
    wire \c0.n4600 ;
    wire data_in_0_6;
    wire data_in_1_3;
    wire data_in_0_0;
    wire \c0.n30 ;
    wire \c0.n25_adj_870_cascade_ ;
    wire \c0.n3933 ;
    wire \c0.n1197_cascade_ ;
    wire \c0.data_in_frame_6_0 ;
    wire data_in_3_5;
    wire \c0.data_in_frame_7_0 ;
    wire data_in_2_6;
    wire rx_data_2;
    wire PIN_2_c;
    wire data_in_1_6;
    wire \c0.n26_adj_869 ;
    wire data_in_2_0;
    wire \c0.n27 ;
    wire \c0.rx.r_Rx_Data_R ;
    wire data_in_1_4;
    wire data_in_1_7;
    wire n11_adj_941;
    wire n4638_cascade_;
    wire tx2_done;
    wire \c0.n4598 ;
    wire \c0.n4807 ;
    wire tx2_data_2_keep_cascade_;
    wire r_Tx_Data_2_adj_962;
    wire n9_adj_939;
    wire n4512_cascade_;
    wire \c0.n4546 ;
    wire \c0.n4603 ;
    wire n1611;
    wire n2326_cascade_;
    wire n4514;
    wire n4512;
    wire n4523;
    wire n4522_cascade_;
    wire n4777;
    wire r_Bit_Index_1;
    wire r_Bit_Index_0_adj_956;
    wire r_Bit_Index_2_adj_955;
    wire \c0.data_in_field_22 ;
    wire \c0.n4556 ;
    wire \c0.n10_adj_874_cascade_ ;
    wire \c0.n4567 ;
    wire data_in_0_7;
    wire \c0.n4541 ;
    wire \c0.n4544 ;
    wire \c0.data_in_field_6 ;
    wire \c0.n1284 ;
    wire \c0.n4408_cascade_ ;
    wire \c0.n4468 ;
    wire data_in_2_3;
    wire data_in_3_2;
    wire data_in_2_5;
    wire \c0.n1271_cascade_ ;
    wire \c0.n4429_cascade_ ;
    wire \c0.n4429 ;
    wire \c0.data_in_field_46 ;
    wire \c0.n6_adj_877 ;
    wire \c0.data_in_field_5 ;
    wire \c0.n4450 ;
    wire data_in_0_4;
    wire \c0.data_in_field_31 ;
    wire \c0.n1261_cascade_ ;
    wire \c0.n4411 ;
    wire \c0.n4411_cascade_ ;
    wire \c0.data_in_frame_6_5 ;
    wire \c0.n4595 ;
    wire \c0.n1340_cascade_ ;
    wire \c0.data_in_field_16 ;
    wire \c0.data_in_field_33 ;
    wire data_in_2_2;
    wire \c0.data_in_field_18 ;
    wire data_in_2_1;
    wire \c0.data_in_field_17 ;
    wire \c0.data_in_field_15 ;
    wire \c0.data_in_field_27 ;
    wire \c0.n4547 ;
    wire data_in_0_3;
    wire \c0.data_in_frame_7_5 ;
    wire \c0.data_in_field_34 ;
    wire \c0.data_in_field_3 ;
    wire \c0.data_in_field_19 ;
    wire \c0.n10 ;
    wire \c0.data_in_field_29 ;
    wire rx_data_3;
    wire data_in_0_1;
    wire data_in_5_5;
    wire data_in_4_5;
    wire \c0.rx.n4873_cascade_ ;
    wire data_in_3_7;
    wire data_in_4_1;
    wire data_in_3_1;
    wire bfn_4_21_0_;
    wire n1710;
    wire \c0.tx2.n3891 ;
    wire \c0.tx2.n3892 ;
    wire \c0.tx2.n3893 ;
    wire \c0.tx2.n3894 ;
    wire n1698;
    wire \c0.tx2.n3895 ;
    wire \c0.tx2.n3896 ;
    wire \c0.tx2.n3897 ;
    wire \c0.tx2.n3898 ;
    wire bfn_4_22_0_;
    wire n1689;
    wire n1704;
    wire n1707;
    wire n1768;
    wire \c0.tx2.r_Clock_Count_0 ;
    wire \c0.tx2.r_Clock_Count_2 ;
    wire \c0.tx2.r_Clock_Count_5 ;
    wire \c0.tx2.r_Clock_Count_1 ;
    wire \c0.tx2.r_Clock_Count_3 ;
    wire \c0.tx2.n5_cascade_ ;
    wire n1701;
    wire \c0.tx2.r_Clock_Count_4 ;
    wire n1692;
    wire \c0.tx2.r_Clock_Count_7 ;
    wire r_SM_Main_2_N_759_1_cascade_;
    wire \c0.tx2.r_Clock_Count_8 ;
    wire \c0.tx2.n2902 ;
    wire n4_adj_965;
    wire \c0.n4543 ;
    wire blink_counter_22;
    wire blink_counter_24;
    wire blink_counter_21;
    wire blink_counter_23;
    wire \c0.n4580 ;
    wire \c0.n4571 ;
    wire \c0.n4855_cascade_ ;
    wire tx2_data_0_keep_cascade_;
    wire r_Tx_Data_0_adj_964;
    wire \c0.data_in_field_32 ;
    wire \c0.n4579 ;
    wire \c0.n4819 ;
    wire \c0.n4549_cascade_ ;
    wire n1030;
    wire tx2_data_4_keep_cascade_;
    wire r_Tx_Data_4_adj_960;
    wire \c0.n4597 ;
    wire \c0.data_in_field_20 ;
    wire \c0.n4550 ;
    wire \c0.tx2.n23 ;
    wire n865_cascade_;
    wire r_SM_Main_2_N_759_1;
    wire n4366_cascade_;
    wire data_in_4_2;
    wire \c0.data_in_field_11 ;
    wire \c0.n8_adj_879_cascade_ ;
    wire \c0.n4451_cascade_ ;
    wire \c0.n8_adj_880 ;
    wire \c0.n10_adj_876 ;
    wire \c0.n4469 ;
    wire \c0.n1357_cascade_ ;
    wire \c0.n4399 ;
    wire \c0.n17 ;
    wire \c0.n4430 ;
    wire \c0.n15_adj_885 ;
    wire \c0.n16_adj_884 ;
    wire \c0.n17_adj_889_cascade_ ;
    wire \c0.n4387_cascade_ ;
    wire data_in_4_7;
    wire data_in_5_7;
    wire \c0.n1296 ;
    wire \c0.n11_adj_888 ;
    wire data_in_2_7;
    wire data_in_1_1;
    wire \c0.n8_adj_871_cascade_ ;
    wire \c0.n12 ;
    wire \c0.n1418 ;
    wire \c0.data_in_field_4 ;
    wire \c0.n1418_cascade_ ;
    wire \c0.n4474_cascade_ ;
    wire data_in_4_6;
    wire \c0.n4396 ;
    wire \c0.data_in_field_21 ;
    wire \c0.n4396_cascade_ ;
    wire \c0.data_in_field_7 ;
    wire \c0.data_in_field_0 ;
    wire \c0.data_in_field_8 ;
    wire \c0.n4570 ;
    wire \c0.data_in_field_39 ;
    wire \c0.data_in_field_38 ;
    wire data_in_6_4;
    wire data_in_4_4;
    wire \c0.n8_adj_872 ;
    wire data_in_0_2;
    wire \c0.data_in_field_2 ;
    wire \c0.data_in_frame_7_1 ;
    wire \c0.n4607 ;
    wire data_in_3_6;
    wire \c0.data_in_frame_6_1 ;
    wire data_in_5_4;
    wire \c0.data_in_field_44 ;
    wire data_in_3_4;
    wire data_in_2_4;
    wire rx_data_5;
    wire rx_data_7;
    wire r_SM_Main_0_adj_954;
    wire r_SM_Main_1_adj_953;
    wire n4780;
    wire r_SM_Main_2_adj_952;
    wire n3_cascade_;
    wire rx_data_6;
    wire \c0.rx.n4876 ;
    wire tx_enable;
    wire data_in_7_5;
    wire data_in_6_5;
    wire n4519;
    wire n4520;
    wire blink_counter_25;
    wire LED_c;
    wire bfn_5_24_0_;
    wire \c0.n3921 ;
    wire \c0.n3922 ;
    wire \c0.n1675 ;
    wire \c0.n688 ;
    wire tx2_active;
    wire \c0.n2643 ;
    wire \c0.n2643_cascade_ ;
    wire \c0.tx2_transmit ;
    wire \c0.n21 ;
    wire \c0.n22_adj_881 ;
    wire \c0.n30_adj_892_cascade_ ;
    wire \c0.n25_adj_893 ;
    wire \c0.n2637 ;
    wire \c0.n1261 ;
    wire \c0.data_in_field_45 ;
    wire \c0.n14 ;
    wire \c0.n12_adj_873 ;
    wire \c0.n16_cascade_ ;
    wire \c0.n15 ;
    wire \c0.n24 ;
    wire \c0.n4388 ;
    wire \c0.n4445 ;
    wire \c0.n26_adj_890 ;
    wire \c0.data_in_frame_6_2 ;
    wire \c0.n1280 ;
    wire \c0.n4390 ;
    wire \c0.data_in_field_47 ;
    wire \c0.n4391 ;
    wire \c0.data_in_field_1 ;
    wire \c0.data_in_field_14 ;
    wire \c0.n4474 ;
    wire \c0.n12_adj_887 ;
    wire data_in_7_7;
    wire data_in_6_7;
    wire \c0.data_in_field_35 ;
    wire \c0.data_in_field_36 ;
    wire \c0.n11 ;
    wire \c0.data_in_field_43 ;
    wire \c0.data_in_field_26 ;
    wire \c0.n4415_cascade_ ;
    wire \c0.data_in_field_9 ;
    wire \c0.n23 ;
    wire \c0.data_in_field_30 ;
    wire \c0.n4927 ;
    wire \c0.n1267 ;
    wire \c0.n4421 ;
    wire \c0.data_in_field_23 ;
    wire \c0.data_in_field_37 ;
    wire \c0.n8_adj_883 ;
    wire \c0.data_in_field_25 ;
    wire \c0.n1290 ;
    wire \c0.n4441 ;
    wire \c0.data_in_field_28 ;
    wire \c0.data_in_field_42 ;
    wire \c0.data_in_field_13 ;
    wire \c0.n4414 ;
    wire data_in_7_3;
    wire data_in_7_6;
    wire tx2_o_adj_949;
    wire tx2_enable;
    wire \c0.data_in_field_12 ;
    wire \c0.data_in_field_40 ;
    wire data_in_6_6;
    wire \c0.data_in_field_41 ;
    wire \c0.n12_adj_878 ;
    wire rx_data_4;
    wire data_in_7_4;
    wire data_in_3_0;
    wire \c0.data_in_field_24 ;
    wire data_in_1_2;
    wire \c0.n1197 ;
    wire \c0.FRAME_MATCHER_wait_for_transmission ;
    wire \c0.data_in_field_10 ;
    wire n2651;
    wire data_in_5_0;
    wire data_in_4_0;
    wire data_in_4_3;
    wire data_in_3_3;
    wire data_in_5_2;
    wire n1222;
    wire n1222_cascade_;
    wire rx_data_0;
    wire n4_adj_950;
    wire n4;
    wire \c0.rx.n2269 ;
    wire \c0.rx.n2269_cascade_ ;
    wire n1227;
    wire n1227_cascade_;
    wire bfn_5_32_0_;
    wire \c0.rx.n3884 ;
    wire \c0.rx.n3885 ;
    wire \c0.rx.n3886 ;
    wire \c0.rx.n3887 ;
    wire \c0.rx.n3888 ;
    wire \c0.rx.n3889 ;
    wire \c0.rx.n3890 ;
    wire n1695;
    wire n6_adj_940;
    wire \c0.tx2.r_Clock_Count_6 ;
    wire bfn_6_25_0_;
    wire \c0.n3906 ;
    wire \c0.n3907 ;
    wire \c0.n3908 ;
    wire \c0.n3909 ;
    wire \c0.n3910 ;
    wire \c0.n3911 ;
    wire \c0.n3912 ;
    wire \c0.n3913 ;
    wire bfn_6_26_0_;
    wire \c0.n3914 ;
    wire \c0.n3915 ;
    wire \c0.n3916 ;
    wire \c0.n3917 ;
    wire \c0.n3918 ;
    wire \c0.n3919 ;
    wire \c0.n3920 ;
    wire \c0.byte_transmit_counter2_2 ;
    wire \c0.byte_transmit_counter2_1 ;
    wire \c0.byte_transmit_counter2_0 ;
    wire \c0.FRAME_MATCHER_wait_for_transmission_N_423 ;
    wire \c0.data_9 ;
    wire \c0.n4619_cascade_ ;
    wire \c0.data_1 ;
    wire data_in_7_2;
    wire data_in_6_2;
    wire \c0.n4517_cascade_ ;
    wire \c0.n4867_cascade_ ;
    wire tx_data_2_keep_cascade_;
    wire \c0.n4564 ;
    wire \c0.n4408 ;
    wire \c0.n1271 ;
    wire \c0.n4409 ;
    wire \c0.rx.n232_cascade_ ;
    wire \c0.n4516 ;
    wire \c0.rx.n1464_cascade_ ;
    wire n1527;
    wire n1527_cascade_;
    wire n2142;
    wire data_in_7_0;
    wire data_in_6_0;
    wire \c0.rx.n232 ;
    wire \c0.rx.r_SM_Main_2_N_816_2_cascade_ ;
    wire \c0.rx.n4678 ;
    wire r_Bit_Index_0;
    wire n4_adj_943;
    wire n223;
    wire \c0.rx.n214 ;
    wire r_Clock_Count_3;
    wire \c0.rx.n214_cascade_ ;
    wire \c0.rx.n4_cascade_ ;
    wire r_Bit_Index_2;
    wire \c0.rx.r_Bit_Index_1 ;
    wire n4_adj_951;
    wire \c0.rx.n4679 ;
    wire \c0.rx.r_Clock_Count_1 ;
    wire n219;
    wire r_Clock_Count_7;
    wire \c0.rx.n4677 ;
    wire n226;
    wire n573_cascade_;
    wire r_Clock_Count_0;
    wire n222;
    wire r_Clock_Count_4;
    wire \c0.rx.n4641_cascade_ ;
    wire \c0.rx.n8 ;
    wire \c0.rx.n4 ;
    wire \c0.rx.n7 ;
    wire \c0.rx.n4093_cascade_ ;
    wire \c0.rx.n2246 ;
    wire n221;
    wire r_Clock_Count_5;
    wire \c0.n4783_cascade_ ;
    wire \c0.n4526 ;
    wire tx_data_3_keep_cascade_;
    wire \c0.n4622 ;
    wire \c0.n4621 ;
    wire \c0.n4525 ;
    wire data_in_6_3;
    wire data_in_5_3;
    wire \c0.n4768_cascade_ ;
    wire tx_data_7_keep_cascade_;
    wire \c0.n4843_cascade_ ;
    wire tx_data_1_keep_cascade_;
    wire r_Tx_Data_7;
    wire \c0.n4585 ;
    wire r_Tx_Data_6;
    wire \c0.n4861_cascade_ ;
    wire tx_data_0_keep_cascade_;
    wire \c0.n4586 ;
    wire \c0.n4573 ;
    wire \c0.n4789 ;
    wire tx_data_4_keep_cascade_;
    wire r_Tx_Data_4;
    wire \c0.n4576 ;
    wire \c0.tx.n4589 ;
    wire \c0.tx.n4588 ;
    wire tx_data_5_keep_cascade_;
    wire r_Tx_Data_5;
    wire \c0.tx.n1588 ;
    wire \c0.tx.n4715_cascade_ ;
    wire rx_data_1;
    wire data_in_7_1;
    wire r_Tx_Data_1;
    wire r_Tx_Data_0;
    wire r_Tx_Data_3;
    wire r_Tx_Data_2;
    wire \c0.tx.n4558 ;
    wire \c0.tx.n4559_cascade_ ;
    wire \c0.tx.n4837 ;
    wire tx_o;
    wire rx_data_ready_keep;
    wire data_in_6_1;
    wire data_in_5_1;
    wire n224;
    wire r_Clock_Count_2;
    wire \c0.n4528 ;
    wire \c0.rx.r_SM_Main_2_N_816_2 ;
    wire \c0.rx.n1024 ;
    wire \c0.tx.o_Tx_Serial_N_790 ;
    wire \c0.tx.n12 ;
    wire \c0.rx.n6_cascade_ ;
    wire \c0.rx.n357 ;
    wire \c0.rx.n4093 ;
    wire \c0.rx.n4378 ;
    wire \c0.rx.n13_cascade_ ;
    wire \c0.rx.n6 ;
    wire n1554;
    wire n220;
    wire n573;
    wire n1554_cascade_;
    wire r_Clock_Count_6;
    wire \c0.rx.n2179 ;
    wire \c0.rx.r_SM_Main_0 ;
    wire r_Rx_Data;
    wire \c0.rx.r_SM_Main_2 ;
    wire \c0.rx.n4666_cascade_ ;
    wire \c0.rx.n4667 ;
    wire \c0.rx.r_SM_Main_1 ;
    wire bfn_9_25_0_;
    wire \c0.n3899 ;
    wire \c0.n3900 ;
    wire \c0.n3901 ;
    wire \c0.n3902 ;
    wire \c0.n3903 ;
    wire \c0.n3904 ;
    wire \c0.n3905 ;
    wire data_out_6_1;
    wire \c0.data_15 ;
    wire \c0.n4888 ;
    wire \c0.n2429 ;
    wire \c0.data_6 ;
    wire \c0.data_7 ;
    wire \c0.data_14 ;
    wire data_out_7_3;
    wire \c0.data_8 ;
    wire n8_adj_932_cascade_;
    wire data_out_7_2;
    wire data_out_7_1;
    wire \c0.n4574 ;
    wire \c0.data_10 ;
    wire data_out_field_19;
    wire n8_adj_936;
    wire data_out_6_2;
    wire \c0.n4565 ;
    wire n11_adj_967_cascade_;
    wire data_out_7_4;
    wire data_out_field_11;
    wire \c0.n6_cascade_ ;
    wire data_out_field_24;
    wire \c0.n4456_cascade_ ;
    wire \c0.data_0 ;
    wire data_out_field_17;
    wire \c0.n4562 ;
    wire \c0.data_out_field_47_N_682_41 ;
    wire \c0.data_out_field_47_N_682_34 ;
    wire \c0.n1384_cascade_ ;
    wire \c0.data_out_field_47_N_682_32 ;
    wire data_out_field_3;
    wire data_out_field_4;
    wire \c0.n4529 ;
    wire n7_adj_937;
    wire \c0.delay_counter_6 ;
    wire \c0.delay_counter_0 ;
    wire \c0.delay_counter_2 ;
    wire \c0.delay_counter_4 ;
    wire \c0.delay_counter_5 ;
    wire \c0.delay_counter_1 ;
    wire \c0.delay_counter_7 ;
    wire \c0.delay_counter_3 ;
    wire \c0.n13 ;
    wire \c0.n14_adj_902_cascade_ ;
    wire \c0.data_4 ;
    wire n3580_cascade_;
    wire \c0.data_11 ;
    wire \c0.data_3 ;
    wire n7_adj_933;
    wire \c0.n4885 ;
    wire \c0.data_5 ;
    wire \c0.n6_adj_904_cascade_ ;
    wire n7_adj_938_cascade_;
    wire data_out_6_3;
    wire \c0.n4380 ;
    wire \c0.data_out_field_47_N_682_33 ;
    wire \c0.n4393 ;
    wire n12_adj_966;
    wire n1677_cascade_;
    wire data_out_6_7;
    wire n7_adj_935;
    wire n8_adj_934_cascade_;
    wire data_out_7_7;
    wire \c0.n1333 ;
    wire \c0.n4447_cascade_ ;
    wire n9_adj_972;
    wire \c0.n4795 ;
    wire n11_adj_945;
    wire n4_adj_970;
    wire data_out_field_16;
    wire \c0.n4447 ;
    wire n7_adj_969_cascade_;
    wire \c0.tx.r_Bit_Index_2 ;
    wire \c0.tx.r_Bit_Index_1 ;
    wire \c0.tx.r_Bit_Index_0 ;
    wire data_out_6_5;
    wire \c0.n4616 ;
    wire data_out_field_25;
    wire \c0.data_out_field_47_N_682_40 ;
    wire \c0.n4561 ;
    wire \c0.data_2 ;
    wire \c0.n4771_cascade_ ;
    wire \c0.n4774_cascade_ ;
    wire tx_data_6_keep;
    wire n10_adj_971;
    wire \c0.data_12 ;
    wire data_out_field_7;
    wire data_out_field_6;
    wire n1246_cascade_;
    wire data_out_field_22;
    wire bfn_11_27_0_;
    wire \c0.n3844 ;
    wire \c0.byte_transmit_counter_2 ;
    wire \c0.n3845 ;
    wire \c0.byte_transmit_counter_3 ;
    wire \c0.tx_transmit_N_274_3 ;
    wire \c0.n3846 ;
    wire \c0.byte_transmit_counter_4 ;
    wire \c0.tx_transmit_N_274_4 ;
    wire \c0.n3847 ;
    wire \c0.byte_transmit_counter_5 ;
    wire \c0.tx_transmit_N_274_5 ;
    wire \c0.n3848 ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.tx_transmit_N_274_6 ;
    wire \c0.n3849 ;
    wire \c0.byte_transmit_counter_7 ;
    wire \c0.n3850 ;
    wire \c0.tx_transmit_N_274_7 ;
    wire \c0.data_out_field_47_N_682_35 ;
    wire n10_adj_947;
    wire n9_adj_948_cascade_;
    wire data_out_field_27;
    wire n4_adj_942;
    wire \c0.n4531 ;
    wire n8_adj_968;
    wire data_out_7_0;
    wire data_out_6_0;
    wire \c0.n4577 ;
    wire n1255;
    wire data_out_6_4;
    wire data_out_field_5;
    wire data_out_field_18;
    wire data_out_field_20;
    wire data_out_field_12;
    wire \c0.n4432_cascade_ ;
    wire \c0.n4417 ;
    wire \c0.n4483 ;
    wire \c0.n10_adj_900_cascade_ ;
    wire n4438;
    wire \c0.n4489 ;
    wire \c0.n4532 ;
    wire n1677;
    wire \c0.n4465 ;
    wire \c0.data_out_7_5 ;
    wire \c0.data_out_field_47_N_682_45 ;
    wire \c0.n4615 ;
    wire data_out_6_6;
    wire data_out_7_6;
    wire \c0.n4879_cascade_ ;
    wire \c0.data_out_field_47_N_682_46 ;
    wire \c0.n4882 ;
    wire data_out_field_13;
    wire data_out_field_28;
    wire \c0.data_out_field_47_N_682_44 ;
    wire \c0.data_out_field_47_N_682_36 ;
    wire \c0.n4618 ;
    wire data_out_field_21;
    wire n1246;
    wire n4663;
    wire \c0.byte_transmit_counter_1 ;
    wire data_out_field_31;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.n4765 ;
    wire data_out_field_14;
    wire \c0.data_out_field_47_N_682_42 ;
    wire n4423;
    wire n4462;
    wire data_out_field_26;
    wire n4655;
    wire data_out_field_2;
    wire data_out_field_43;
    wire data_out_field_15;
    wire data_out_field_30;
    wire \c0.tx.n1514 ;
    wire data_out_field_38;
    wire data_out_field_9;
    wire \c0.data_out_field_47_N_682_39 ;
    wire n4426;
    wire n4426_cascade_;
    wire data_out_field_10;
    wire n4659;
    wire \c0.data_13 ;
    wire \c0.data_out_field_47_N_682_37 ;
    wire n3580;
    wire n7_adj_938;
    wire data_out_field_1;
    wire data_out_field_29;
    wire \c0.n4453 ;
    wire \c0.n1312 ;
    wire \c0.n1306_cascade_ ;
    wire \c0.data_out_field_47_N_682_47 ;
    wire n4454;
    wire \c0.tx_active_prev ;
    wire \c0.n50 ;
    wire \c0.tx.n2908_cascade_ ;
    wire \c0.tx.n1457_cascade_ ;
    wire \c0.tx_active ;
    wire data_out_field_8;
    wire data_out_field_23;
    wire n1325;
    wire n1025;
    wire \c0.tx.n752 ;
    wire \c0.tx_transmit ;
    wire data_out_field_0;
    wire \c0.n1421 ;
    wire \c0.n1306 ;
    wire \c0.tx.n6 ;
    wire \c0.tx.n5_cascade_ ;
    wire \c0.tx.n17_cascade_ ;
    wire \c0.n1378 ;
    wire \c0.n4477 ;
    wire n4480;
    wire \c0.n4456 ;
    wire n12_adj_944;
    wire n4_adj_946_cascade_;
    wire n88;
    wire tx_done;
    wire \c0.tx.n84 ;
    wire \c0.tx.n3643 ;
    wire r_SM_Main_1;
    wire n4375;
    wire \c0.tx.n25_cascade_ ;
    wire \c0.tx.n17 ;
    wire r_SM_Main_0;
    wire CLK_c;
    wire \c0.tx.r_Clock_Count_0 ;
    wire \c0.tx.n1979 ;
    wire bfn_14_27_0_;
    wire \c0.tx.r_Clock_Count_1 ;
    wire \c0.tx.n1754 ;
    wire \c0.tx.n3876 ;
    wire \c0.tx.r_Clock_Count_2 ;
    wire \c0.tx.n1751 ;
    wire \c0.tx.n3877 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire \c0.tx.n1748 ;
    wire \c0.tx.n3878 ;
    wire \c0.tx.r_Clock_Count_4 ;
    wire \c0.tx.n1745 ;
    wire \c0.tx.n3879 ;
    wire \c0.tx.r_Clock_Count_5 ;
    wire \c0.tx.n1742 ;
    wire \c0.tx.n3880 ;
    wire \c0.tx.r_Clock_Count_6 ;
    wire \c0.tx.n1739 ;
    wire \c0.tx.n3881 ;
    wire \c0.tx.r_Clock_Count_7 ;
    wire \c0.tx.n1736 ;
    wire \c0.tx.n3882 ;
    wire \c0.tx.n3883 ;
    wire \c0.tx.r_Clock_Count_8 ;
    wire r_SM_Main_2;
    wire bfn_14_28_0_;
    wire \c0.tx.n1733 ;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__23697),
            .DIN(N__23696),
            .DOUT(N__23695),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__23697),
            .PADOUT(N__23696),
            .PADIN(N__23695),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12218),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_2_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_2_pad_iopad (
            .OE(N__23688),
            .DIN(N__23687),
            .DOUT(N__23686),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_2_pad_preio (
            .PADOEN(N__23688),
            .PADOUT(N__23687),
            .PADIN(N__23686),
            .CLOCKENABLE(),
            .DIN0(PIN_2_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__23679),
            .DIN(N__23678),
            .DOUT(N__23677),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__23679),
            .PADOUT(N__23678),
            .PADIN(N__23677),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx2_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx2_output_iopad.PULLUP=1'b1;
    IO_PAD tx2_output_iopad (
            .OE(N__23670),
            .DIN(N__23669),
            .DOUT(N__23668),
            .PACKAGEPIN(PIN_3));
    defparam tx2_output_preio.PIN_TYPE=6'b101001;
    defparam tx2_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx2_output_preio (
            .PADOEN(N__23670),
            .PADOUT(N__23669),
            .PADIN(N__23668),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14060),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__14033));
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__23661),
            .DIN(N__23660),
            .DOUT(N__23659),
            .PACKAGEPIN(PIN_1));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__23661),
            .PADOUT(N__23660),
            .PADIN(N__23659),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__17162),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__12317));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__23652),
            .DIN(N__23651),
            .DOUT(N__23650),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__23652),
            .PADOUT(N__23651),
            .PADIN(N__23650),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__5783 (
            .O(N__23633),
            .I(N__23628));
    InMux I__5782 (
            .O(N__23632),
            .I(N__23625));
    InMux I__5781 (
            .O(N__23631),
            .I(N__23622));
    LocalMux I__5780 (
            .O(N__23628),
            .I(\c0.tx.r_Clock_Count_4 ));
    LocalMux I__5779 (
            .O(N__23625),
            .I(\c0.tx.r_Clock_Count_4 ));
    LocalMux I__5778 (
            .O(N__23622),
            .I(\c0.tx.r_Clock_Count_4 ));
    InMux I__5777 (
            .O(N__23615),
            .I(N__23612));
    LocalMux I__5776 (
            .O(N__23612),
            .I(\c0.tx.n1745 ));
    InMux I__5775 (
            .O(N__23609),
            .I(\c0.tx.n3879 ));
    InMux I__5774 (
            .O(N__23606),
            .I(N__23601));
    InMux I__5773 (
            .O(N__23605),
            .I(N__23598));
    InMux I__5772 (
            .O(N__23604),
            .I(N__23595));
    LocalMux I__5771 (
            .O(N__23601),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__5770 (
            .O(N__23598),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__5769 (
            .O(N__23595),
            .I(\c0.tx.r_Clock_Count_5 ));
    CascadeMux I__5768 (
            .O(N__23588),
            .I(N__23585));
    InMux I__5767 (
            .O(N__23585),
            .I(N__23582));
    LocalMux I__5766 (
            .O(N__23582),
            .I(\c0.tx.n1742 ));
    InMux I__5765 (
            .O(N__23579),
            .I(\c0.tx.n3880 ));
    InMux I__5764 (
            .O(N__23576),
            .I(N__23571));
    InMux I__5763 (
            .O(N__23575),
            .I(N__23568));
    InMux I__5762 (
            .O(N__23574),
            .I(N__23565));
    LocalMux I__5761 (
            .O(N__23571),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__5760 (
            .O(N__23568),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__5759 (
            .O(N__23565),
            .I(\c0.tx.r_Clock_Count_6 ));
    InMux I__5758 (
            .O(N__23558),
            .I(N__23555));
    LocalMux I__5757 (
            .O(N__23555),
            .I(\c0.tx.n1739 ));
    InMux I__5756 (
            .O(N__23552),
            .I(\c0.tx.n3881 ));
    InMux I__5755 (
            .O(N__23549),
            .I(N__23544));
    InMux I__5754 (
            .O(N__23548),
            .I(N__23541));
    InMux I__5753 (
            .O(N__23547),
            .I(N__23538));
    LocalMux I__5752 (
            .O(N__23544),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__5751 (
            .O(N__23541),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__5750 (
            .O(N__23538),
            .I(\c0.tx.r_Clock_Count_7 ));
    InMux I__5749 (
            .O(N__23531),
            .I(N__23528));
    LocalMux I__5748 (
            .O(N__23528),
            .I(\c0.tx.n1736 ));
    InMux I__5747 (
            .O(N__23525),
            .I(\c0.tx.n3882 ));
    InMux I__5746 (
            .O(N__23522),
            .I(N__23517));
    InMux I__5745 (
            .O(N__23521),
            .I(N__23514));
    InMux I__5744 (
            .O(N__23520),
            .I(N__23511));
    LocalMux I__5743 (
            .O(N__23517),
            .I(N__23508));
    LocalMux I__5742 (
            .O(N__23514),
            .I(\c0.tx.r_Clock_Count_8 ));
    LocalMux I__5741 (
            .O(N__23511),
            .I(\c0.tx.r_Clock_Count_8 ));
    Odrv4 I__5740 (
            .O(N__23508),
            .I(\c0.tx.r_Clock_Count_8 ));
    InMux I__5739 (
            .O(N__23501),
            .I(N__23498));
    LocalMux I__5738 (
            .O(N__23498),
            .I(N__23495));
    Span4Mux_s2_v I__5737 (
            .O(N__23495),
            .I(N__23490));
    CascadeMux I__5736 (
            .O(N__23494),
            .I(N__23487));
    CascadeMux I__5735 (
            .O(N__23493),
            .I(N__23460));
    Span4Mux_h I__5734 (
            .O(N__23490),
            .I(N__23457));
    InMux I__5733 (
            .O(N__23487),
            .I(N__23454));
    CascadeMux I__5732 (
            .O(N__23486),
            .I(N__23450));
    CascadeMux I__5731 (
            .O(N__23485),
            .I(N__23447));
    CascadeMux I__5730 (
            .O(N__23484),
            .I(N__23444));
    CascadeMux I__5729 (
            .O(N__23483),
            .I(N__23441));
    CascadeMux I__5728 (
            .O(N__23482),
            .I(N__23438));
    CascadeMux I__5727 (
            .O(N__23481),
            .I(N__23435));
    CascadeMux I__5726 (
            .O(N__23480),
            .I(N__23432));
    CascadeMux I__5725 (
            .O(N__23479),
            .I(N__23429));
    InMux I__5724 (
            .O(N__23478),
            .I(N__23422));
    InMux I__5723 (
            .O(N__23477),
            .I(N__23422));
    InMux I__5722 (
            .O(N__23476),
            .I(N__23422));
    InMux I__5721 (
            .O(N__23475),
            .I(N__23419));
    InMux I__5720 (
            .O(N__23474),
            .I(N__23416));
    InMux I__5719 (
            .O(N__23473),
            .I(N__23413));
    InMux I__5718 (
            .O(N__23472),
            .I(N__23408));
    InMux I__5717 (
            .O(N__23471),
            .I(N__23408));
    InMux I__5716 (
            .O(N__23470),
            .I(N__23405));
    InMux I__5715 (
            .O(N__23469),
            .I(N__23396));
    InMux I__5714 (
            .O(N__23468),
            .I(N__23396));
    InMux I__5713 (
            .O(N__23467),
            .I(N__23396));
    InMux I__5712 (
            .O(N__23466),
            .I(N__23396));
    InMux I__5711 (
            .O(N__23465),
            .I(N__23387));
    InMux I__5710 (
            .O(N__23464),
            .I(N__23387));
    InMux I__5709 (
            .O(N__23463),
            .I(N__23387));
    InMux I__5708 (
            .O(N__23460),
            .I(N__23387));
    Span4Mux_v I__5707 (
            .O(N__23457),
            .I(N__23384));
    LocalMux I__5706 (
            .O(N__23454),
            .I(N__23381));
    InMux I__5705 (
            .O(N__23453),
            .I(N__23378));
    InMux I__5704 (
            .O(N__23450),
            .I(N__23369));
    InMux I__5703 (
            .O(N__23447),
            .I(N__23369));
    InMux I__5702 (
            .O(N__23444),
            .I(N__23369));
    InMux I__5701 (
            .O(N__23441),
            .I(N__23369));
    InMux I__5700 (
            .O(N__23438),
            .I(N__23360));
    InMux I__5699 (
            .O(N__23435),
            .I(N__23360));
    InMux I__5698 (
            .O(N__23432),
            .I(N__23360));
    InMux I__5697 (
            .O(N__23429),
            .I(N__23360));
    LocalMux I__5696 (
            .O(N__23422),
            .I(N__23349));
    LocalMux I__5695 (
            .O(N__23419),
            .I(N__23349));
    LocalMux I__5694 (
            .O(N__23416),
            .I(N__23349));
    LocalMux I__5693 (
            .O(N__23413),
            .I(N__23349));
    LocalMux I__5692 (
            .O(N__23408),
            .I(N__23349));
    LocalMux I__5691 (
            .O(N__23405),
            .I(r_SM_Main_2));
    LocalMux I__5690 (
            .O(N__23396),
            .I(r_SM_Main_2));
    LocalMux I__5689 (
            .O(N__23387),
            .I(r_SM_Main_2));
    Odrv4 I__5688 (
            .O(N__23384),
            .I(r_SM_Main_2));
    Odrv4 I__5687 (
            .O(N__23381),
            .I(r_SM_Main_2));
    LocalMux I__5686 (
            .O(N__23378),
            .I(r_SM_Main_2));
    LocalMux I__5685 (
            .O(N__23369),
            .I(r_SM_Main_2));
    LocalMux I__5684 (
            .O(N__23360),
            .I(r_SM_Main_2));
    Odrv4 I__5683 (
            .O(N__23349),
            .I(r_SM_Main_2));
    InMux I__5682 (
            .O(N__23330),
            .I(bfn_14_28_0_));
    InMux I__5681 (
            .O(N__23327),
            .I(N__23324));
    LocalMux I__5680 (
            .O(N__23324),
            .I(\c0.tx.n1733 ));
    CascadeMux I__5679 (
            .O(N__23321),
            .I(n4_adj_946_cascade_));
    CascadeMux I__5678 (
            .O(N__23318),
            .I(N__23310));
    InMux I__5677 (
            .O(N__23317),
            .I(N__23299));
    InMux I__5676 (
            .O(N__23316),
            .I(N__23299));
    InMux I__5675 (
            .O(N__23315),
            .I(N__23299));
    InMux I__5674 (
            .O(N__23314),
            .I(N__23288));
    InMux I__5673 (
            .O(N__23313),
            .I(N__23288));
    InMux I__5672 (
            .O(N__23310),
            .I(N__23288));
    InMux I__5671 (
            .O(N__23309),
            .I(N__23288));
    InMux I__5670 (
            .O(N__23308),
            .I(N__23288));
    CascadeMux I__5669 (
            .O(N__23307),
            .I(N__23285));
    InMux I__5668 (
            .O(N__23306),
            .I(N__23282));
    LocalMux I__5667 (
            .O(N__23299),
            .I(N__23279));
    LocalMux I__5666 (
            .O(N__23288),
            .I(N__23276));
    InMux I__5665 (
            .O(N__23285),
            .I(N__23273));
    LocalMux I__5664 (
            .O(N__23282),
            .I(n88));
    Odrv4 I__5663 (
            .O(N__23279),
            .I(n88));
    Odrv4 I__5662 (
            .O(N__23276),
            .I(n88));
    LocalMux I__5661 (
            .O(N__23273),
            .I(n88));
    CascadeMux I__5660 (
            .O(N__23264),
            .I(N__23260));
    InMux I__5659 (
            .O(N__23263),
            .I(N__23257));
    InMux I__5658 (
            .O(N__23260),
            .I(N__23254));
    LocalMux I__5657 (
            .O(N__23257),
            .I(tx_done));
    LocalMux I__5656 (
            .O(N__23254),
            .I(tx_done));
    InMux I__5655 (
            .O(N__23249),
            .I(N__23246));
    LocalMux I__5654 (
            .O(N__23246),
            .I(N__23241));
    InMux I__5653 (
            .O(N__23245),
            .I(N__23238));
    InMux I__5652 (
            .O(N__23244),
            .I(N__23235));
    Span4Mux_v I__5651 (
            .O(N__23241),
            .I(N__23232));
    LocalMux I__5650 (
            .O(N__23238),
            .I(N__23229));
    LocalMux I__5649 (
            .O(N__23235),
            .I(N__23226));
    Span4Mux_h I__5648 (
            .O(N__23232),
            .I(N__23221));
    Span4Mux_h I__5647 (
            .O(N__23229),
            .I(N__23221));
    Span4Mux_h I__5646 (
            .O(N__23226),
            .I(N__23218));
    Odrv4 I__5645 (
            .O(N__23221),
            .I(\c0.tx.n84 ));
    Odrv4 I__5644 (
            .O(N__23218),
            .I(\c0.tx.n84 ));
    InMux I__5643 (
            .O(N__23213),
            .I(N__23210));
    LocalMux I__5642 (
            .O(N__23210),
            .I(\c0.tx.n3643 ));
    InMux I__5641 (
            .O(N__23207),
            .I(N__23202));
    InMux I__5640 (
            .O(N__23206),
            .I(N__23197));
    InMux I__5639 (
            .O(N__23205),
            .I(N__23194));
    LocalMux I__5638 (
            .O(N__23202),
            .I(N__23190));
    CascadeMux I__5637 (
            .O(N__23201),
            .I(N__23186));
    CascadeMux I__5636 (
            .O(N__23200),
            .I(N__23183));
    LocalMux I__5635 (
            .O(N__23197),
            .I(N__23179));
    LocalMux I__5634 (
            .O(N__23194),
            .I(N__23176));
    CascadeMux I__5633 (
            .O(N__23193),
            .I(N__23173));
    Span4Mux_v I__5632 (
            .O(N__23190),
            .I(N__23169));
    InMux I__5631 (
            .O(N__23189),
            .I(N__23166));
    InMux I__5630 (
            .O(N__23186),
            .I(N__23163));
    InMux I__5629 (
            .O(N__23183),
            .I(N__23155));
    InMux I__5628 (
            .O(N__23182),
            .I(N__23155));
    Span4Mux_s3_v I__5627 (
            .O(N__23179),
            .I(N__23150));
    Span4Mux_v I__5626 (
            .O(N__23176),
            .I(N__23150));
    InMux I__5625 (
            .O(N__23173),
            .I(N__23145));
    InMux I__5624 (
            .O(N__23172),
            .I(N__23145));
    Span4Mux_h I__5623 (
            .O(N__23169),
            .I(N__23142));
    LocalMux I__5622 (
            .O(N__23166),
            .I(N__23137));
    LocalMux I__5621 (
            .O(N__23163),
            .I(N__23137));
    InMux I__5620 (
            .O(N__23162),
            .I(N__23130));
    InMux I__5619 (
            .O(N__23161),
            .I(N__23130));
    InMux I__5618 (
            .O(N__23160),
            .I(N__23130));
    LocalMux I__5617 (
            .O(N__23155),
            .I(N__23125));
    Span4Mux_h I__5616 (
            .O(N__23150),
            .I(N__23125));
    LocalMux I__5615 (
            .O(N__23145),
            .I(r_SM_Main_1));
    Odrv4 I__5614 (
            .O(N__23142),
            .I(r_SM_Main_1));
    Odrv4 I__5613 (
            .O(N__23137),
            .I(r_SM_Main_1));
    LocalMux I__5612 (
            .O(N__23130),
            .I(r_SM_Main_1));
    Odrv4 I__5611 (
            .O(N__23125),
            .I(r_SM_Main_1));
    InMux I__5610 (
            .O(N__23114),
            .I(N__23108));
    InMux I__5609 (
            .O(N__23113),
            .I(N__23108));
    LocalMux I__5608 (
            .O(N__23108),
            .I(n4375));
    CascadeMux I__5607 (
            .O(N__23105),
            .I(\c0.tx.n25_cascade_ ));
    CascadeMux I__5606 (
            .O(N__23102),
            .I(N__23093));
    CascadeMux I__5605 (
            .O(N__23101),
            .I(N__23090));
    CascadeMux I__5604 (
            .O(N__23100),
            .I(N__23087));
    CascadeMux I__5603 (
            .O(N__23099),
            .I(N__23084));
    CascadeMux I__5602 (
            .O(N__23098),
            .I(N__23081));
    InMux I__5601 (
            .O(N__23097),
            .I(N__23073));
    InMux I__5600 (
            .O(N__23096),
            .I(N__23073));
    InMux I__5599 (
            .O(N__23093),
            .I(N__23062));
    InMux I__5598 (
            .O(N__23090),
            .I(N__23062));
    InMux I__5597 (
            .O(N__23087),
            .I(N__23062));
    InMux I__5596 (
            .O(N__23084),
            .I(N__23057));
    InMux I__5595 (
            .O(N__23081),
            .I(N__23057));
    InMux I__5594 (
            .O(N__23080),
            .I(N__23054));
    InMux I__5593 (
            .O(N__23079),
            .I(N__23049));
    InMux I__5592 (
            .O(N__23078),
            .I(N__23049));
    LocalMux I__5591 (
            .O(N__23073),
            .I(N__23046));
    InMux I__5590 (
            .O(N__23072),
            .I(N__23043));
    InMux I__5589 (
            .O(N__23071),
            .I(N__23038));
    InMux I__5588 (
            .O(N__23070),
            .I(N__23038));
    InMux I__5587 (
            .O(N__23069),
            .I(N__23035));
    LocalMux I__5586 (
            .O(N__23062),
            .I(\c0.tx.n17 ));
    LocalMux I__5585 (
            .O(N__23057),
            .I(\c0.tx.n17 ));
    LocalMux I__5584 (
            .O(N__23054),
            .I(\c0.tx.n17 ));
    LocalMux I__5583 (
            .O(N__23049),
            .I(\c0.tx.n17 ));
    Odrv4 I__5582 (
            .O(N__23046),
            .I(\c0.tx.n17 ));
    LocalMux I__5581 (
            .O(N__23043),
            .I(\c0.tx.n17 ));
    LocalMux I__5580 (
            .O(N__23038),
            .I(\c0.tx.n17 ));
    LocalMux I__5579 (
            .O(N__23035),
            .I(\c0.tx.n17 ));
    InMux I__5578 (
            .O(N__23018),
            .I(N__23015));
    LocalMux I__5577 (
            .O(N__23015),
            .I(N__23010));
    InMux I__5576 (
            .O(N__23014),
            .I(N__23007));
    InMux I__5575 (
            .O(N__23013),
            .I(N__23004));
    Span4Mux_h I__5574 (
            .O(N__23010),
            .I(N__22997));
    LocalMux I__5573 (
            .O(N__23007),
            .I(N__22994));
    LocalMux I__5572 (
            .O(N__23004),
            .I(N__22988));
    InMux I__5571 (
            .O(N__23003),
            .I(N__22979));
    InMux I__5570 (
            .O(N__23002),
            .I(N__22979));
    InMux I__5569 (
            .O(N__23001),
            .I(N__22979));
    InMux I__5568 (
            .O(N__23000),
            .I(N__22979));
    Span4Mux_h I__5567 (
            .O(N__22997),
            .I(N__22974));
    Span4Mux_h I__5566 (
            .O(N__22994),
            .I(N__22974));
    InMux I__5565 (
            .O(N__22993),
            .I(N__22967));
    InMux I__5564 (
            .O(N__22992),
            .I(N__22967));
    InMux I__5563 (
            .O(N__22991),
            .I(N__22967));
    Odrv12 I__5562 (
            .O(N__22988),
            .I(r_SM_Main_0));
    LocalMux I__5561 (
            .O(N__22979),
            .I(r_SM_Main_0));
    Odrv4 I__5560 (
            .O(N__22974),
            .I(r_SM_Main_0));
    LocalMux I__5559 (
            .O(N__22967),
            .I(r_SM_Main_0));
    ClkMux I__5558 (
            .O(N__22958),
            .I(N__22679));
    ClkMux I__5557 (
            .O(N__22957),
            .I(N__22679));
    ClkMux I__5556 (
            .O(N__22956),
            .I(N__22679));
    ClkMux I__5555 (
            .O(N__22955),
            .I(N__22679));
    ClkMux I__5554 (
            .O(N__22954),
            .I(N__22679));
    ClkMux I__5553 (
            .O(N__22953),
            .I(N__22679));
    ClkMux I__5552 (
            .O(N__22952),
            .I(N__22679));
    ClkMux I__5551 (
            .O(N__22951),
            .I(N__22679));
    ClkMux I__5550 (
            .O(N__22950),
            .I(N__22679));
    ClkMux I__5549 (
            .O(N__22949),
            .I(N__22679));
    ClkMux I__5548 (
            .O(N__22948),
            .I(N__22679));
    ClkMux I__5547 (
            .O(N__22947),
            .I(N__22679));
    ClkMux I__5546 (
            .O(N__22946),
            .I(N__22679));
    ClkMux I__5545 (
            .O(N__22945),
            .I(N__22679));
    ClkMux I__5544 (
            .O(N__22944),
            .I(N__22679));
    ClkMux I__5543 (
            .O(N__22943),
            .I(N__22679));
    ClkMux I__5542 (
            .O(N__22942),
            .I(N__22679));
    ClkMux I__5541 (
            .O(N__22941),
            .I(N__22679));
    ClkMux I__5540 (
            .O(N__22940),
            .I(N__22679));
    ClkMux I__5539 (
            .O(N__22939),
            .I(N__22679));
    ClkMux I__5538 (
            .O(N__22938),
            .I(N__22679));
    ClkMux I__5537 (
            .O(N__22937),
            .I(N__22679));
    ClkMux I__5536 (
            .O(N__22936),
            .I(N__22679));
    ClkMux I__5535 (
            .O(N__22935),
            .I(N__22679));
    ClkMux I__5534 (
            .O(N__22934),
            .I(N__22679));
    ClkMux I__5533 (
            .O(N__22933),
            .I(N__22679));
    ClkMux I__5532 (
            .O(N__22932),
            .I(N__22679));
    ClkMux I__5531 (
            .O(N__22931),
            .I(N__22679));
    ClkMux I__5530 (
            .O(N__22930),
            .I(N__22679));
    ClkMux I__5529 (
            .O(N__22929),
            .I(N__22679));
    ClkMux I__5528 (
            .O(N__22928),
            .I(N__22679));
    ClkMux I__5527 (
            .O(N__22927),
            .I(N__22679));
    ClkMux I__5526 (
            .O(N__22926),
            .I(N__22679));
    ClkMux I__5525 (
            .O(N__22925),
            .I(N__22679));
    ClkMux I__5524 (
            .O(N__22924),
            .I(N__22679));
    ClkMux I__5523 (
            .O(N__22923),
            .I(N__22679));
    ClkMux I__5522 (
            .O(N__22922),
            .I(N__22679));
    ClkMux I__5521 (
            .O(N__22921),
            .I(N__22679));
    ClkMux I__5520 (
            .O(N__22920),
            .I(N__22679));
    ClkMux I__5519 (
            .O(N__22919),
            .I(N__22679));
    ClkMux I__5518 (
            .O(N__22918),
            .I(N__22679));
    ClkMux I__5517 (
            .O(N__22917),
            .I(N__22679));
    ClkMux I__5516 (
            .O(N__22916),
            .I(N__22679));
    ClkMux I__5515 (
            .O(N__22915),
            .I(N__22679));
    ClkMux I__5514 (
            .O(N__22914),
            .I(N__22679));
    ClkMux I__5513 (
            .O(N__22913),
            .I(N__22679));
    ClkMux I__5512 (
            .O(N__22912),
            .I(N__22679));
    ClkMux I__5511 (
            .O(N__22911),
            .I(N__22679));
    ClkMux I__5510 (
            .O(N__22910),
            .I(N__22679));
    ClkMux I__5509 (
            .O(N__22909),
            .I(N__22679));
    ClkMux I__5508 (
            .O(N__22908),
            .I(N__22679));
    ClkMux I__5507 (
            .O(N__22907),
            .I(N__22679));
    ClkMux I__5506 (
            .O(N__22906),
            .I(N__22679));
    ClkMux I__5505 (
            .O(N__22905),
            .I(N__22679));
    ClkMux I__5504 (
            .O(N__22904),
            .I(N__22679));
    ClkMux I__5503 (
            .O(N__22903),
            .I(N__22679));
    ClkMux I__5502 (
            .O(N__22902),
            .I(N__22679));
    ClkMux I__5501 (
            .O(N__22901),
            .I(N__22679));
    ClkMux I__5500 (
            .O(N__22900),
            .I(N__22679));
    ClkMux I__5499 (
            .O(N__22899),
            .I(N__22679));
    ClkMux I__5498 (
            .O(N__22898),
            .I(N__22679));
    ClkMux I__5497 (
            .O(N__22897),
            .I(N__22679));
    ClkMux I__5496 (
            .O(N__22896),
            .I(N__22679));
    ClkMux I__5495 (
            .O(N__22895),
            .I(N__22679));
    ClkMux I__5494 (
            .O(N__22894),
            .I(N__22679));
    ClkMux I__5493 (
            .O(N__22893),
            .I(N__22679));
    ClkMux I__5492 (
            .O(N__22892),
            .I(N__22679));
    ClkMux I__5491 (
            .O(N__22891),
            .I(N__22679));
    ClkMux I__5490 (
            .O(N__22890),
            .I(N__22679));
    ClkMux I__5489 (
            .O(N__22889),
            .I(N__22679));
    ClkMux I__5488 (
            .O(N__22888),
            .I(N__22679));
    ClkMux I__5487 (
            .O(N__22887),
            .I(N__22679));
    ClkMux I__5486 (
            .O(N__22886),
            .I(N__22679));
    ClkMux I__5485 (
            .O(N__22885),
            .I(N__22679));
    ClkMux I__5484 (
            .O(N__22884),
            .I(N__22679));
    ClkMux I__5483 (
            .O(N__22883),
            .I(N__22679));
    ClkMux I__5482 (
            .O(N__22882),
            .I(N__22679));
    ClkMux I__5481 (
            .O(N__22881),
            .I(N__22679));
    ClkMux I__5480 (
            .O(N__22880),
            .I(N__22679));
    ClkMux I__5479 (
            .O(N__22879),
            .I(N__22679));
    ClkMux I__5478 (
            .O(N__22878),
            .I(N__22679));
    ClkMux I__5477 (
            .O(N__22877),
            .I(N__22679));
    ClkMux I__5476 (
            .O(N__22876),
            .I(N__22679));
    ClkMux I__5475 (
            .O(N__22875),
            .I(N__22679));
    ClkMux I__5474 (
            .O(N__22874),
            .I(N__22679));
    ClkMux I__5473 (
            .O(N__22873),
            .I(N__22679));
    ClkMux I__5472 (
            .O(N__22872),
            .I(N__22679));
    ClkMux I__5471 (
            .O(N__22871),
            .I(N__22679));
    ClkMux I__5470 (
            .O(N__22870),
            .I(N__22679));
    ClkMux I__5469 (
            .O(N__22869),
            .I(N__22679));
    ClkMux I__5468 (
            .O(N__22868),
            .I(N__22679));
    ClkMux I__5467 (
            .O(N__22867),
            .I(N__22679));
    ClkMux I__5466 (
            .O(N__22866),
            .I(N__22679));
    GlobalMux I__5465 (
            .O(N__22679),
            .I(N__22676));
    gio2CtrlBuf I__5464 (
            .O(N__22676),
            .I(CLK_c));
    InMux I__5463 (
            .O(N__22673),
            .I(N__22669));
    InMux I__5462 (
            .O(N__22672),
            .I(N__22666));
    LocalMux I__5461 (
            .O(N__22669),
            .I(\c0.tx.r_Clock_Count_0 ));
    LocalMux I__5460 (
            .O(N__22666),
            .I(\c0.tx.r_Clock_Count_0 ));
    InMux I__5459 (
            .O(N__22661),
            .I(N__22658));
    LocalMux I__5458 (
            .O(N__22658),
            .I(\c0.tx.n1979 ));
    InMux I__5457 (
            .O(N__22655),
            .I(bfn_14_27_0_));
    InMux I__5456 (
            .O(N__22652),
            .I(N__22647));
    InMux I__5455 (
            .O(N__22651),
            .I(N__22644));
    InMux I__5454 (
            .O(N__22650),
            .I(N__22641));
    LocalMux I__5453 (
            .O(N__22647),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__5452 (
            .O(N__22644),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__5451 (
            .O(N__22641),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__5450 (
            .O(N__22634),
            .I(N__22631));
    LocalMux I__5449 (
            .O(N__22631),
            .I(\c0.tx.n1754 ));
    InMux I__5448 (
            .O(N__22628),
            .I(\c0.tx.n3876 ));
    CascadeMux I__5447 (
            .O(N__22625),
            .I(N__22620));
    InMux I__5446 (
            .O(N__22624),
            .I(N__22617));
    InMux I__5445 (
            .O(N__22623),
            .I(N__22614));
    InMux I__5444 (
            .O(N__22620),
            .I(N__22611));
    LocalMux I__5443 (
            .O(N__22617),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__5442 (
            .O(N__22614),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__5441 (
            .O(N__22611),
            .I(\c0.tx.r_Clock_Count_2 ));
    InMux I__5440 (
            .O(N__22604),
            .I(N__22601));
    LocalMux I__5439 (
            .O(N__22601),
            .I(\c0.tx.n1751 ));
    InMux I__5438 (
            .O(N__22598),
            .I(\c0.tx.n3877 ));
    InMux I__5437 (
            .O(N__22595),
            .I(N__22590));
    InMux I__5436 (
            .O(N__22594),
            .I(N__22587));
    InMux I__5435 (
            .O(N__22593),
            .I(N__22584));
    LocalMux I__5434 (
            .O(N__22590),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__5433 (
            .O(N__22587),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__5432 (
            .O(N__22584),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__5431 (
            .O(N__22577),
            .I(N__22574));
    LocalMux I__5430 (
            .O(N__22574),
            .I(\c0.tx.n1748 ));
    InMux I__5429 (
            .O(N__22571),
            .I(\c0.tx.n3878 ));
    InMux I__5428 (
            .O(N__22568),
            .I(N__22565));
    LocalMux I__5427 (
            .O(N__22565),
            .I(\c0.tx.n6 ));
    CascadeMux I__5426 (
            .O(N__22562),
            .I(\c0.tx.n5_cascade_ ));
    CascadeMux I__5425 (
            .O(N__22559),
            .I(\c0.tx.n17_cascade_ ));
    InMux I__5424 (
            .O(N__22556),
            .I(N__22553));
    LocalMux I__5423 (
            .O(N__22553),
            .I(N__22550));
    Odrv4 I__5422 (
            .O(N__22550),
            .I(\c0.n1378 ));
    InMux I__5421 (
            .O(N__22547),
            .I(N__22544));
    LocalMux I__5420 (
            .O(N__22544),
            .I(N__22541));
    Span4Mux_h I__5419 (
            .O(N__22541),
            .I(N__22537));
    InMux I__5418 (
            .O(N__22540),
            .I(N__22534));
    Odrv4 I__5417 (
            .O(N__22537),
            .I(\c0.n4477 ));
    LocalMux I__5416 (
            .O(N__22534),
            .I(\c0.n4477 ));
    CascadeMux I__5415 (
            .O(N__22529),
            .I(N__22526));
    InMux I__5414 (
            .O(N__22526),
            .I(N__22522));
    InMux I__5413 (
            .O(N__22525),
            .I(N__22519));
    LocalMux I__5412 (
            .O(N__22522),
            .I(N__22516));
    LocalMux I__5411 (
            .O(N__22519),
            .I(N__22513));
    Span4Mux_h I__5410 (
            .O(N__22516),
            .I(N__22510));
    Span4Mux_h I__5409 (
            .O(N__22513),
            .I(N__22507));
    Odrv4 I__5408 (
            .O(N__22510),
            .I(n4480));
    Odrv4 I__5407 (
            .O(N__22507),
            .I(n4480));
    InMux I__5406 (
            .O(N__22502),
            .I(N__22499));
    LocalMux I__5405 (
            .O(N__22499),
            .I(N__22496));
    Span4Mux_h I__5404 (
            .O(N__22496),
            .I(N__22493));
    Odrv4 I__5403 (
            .O(N__22493),
            .I(\c0.n4456 ));
    InMux I__5402 (
            .O(N__22490),
            .I(N__22487));
    LocalMux I__5401 (
            .O(N__22487),
            .I(N__22484));
    Odrv12 I__5400 (
            .O(N__22484),
            .I(n12_adj_944));
    CascadeMux I__5399 (
            .O(N__22481),
            .I(N__22478));
    InMux I__5398 (
            .O(N__22478),
            .I(N__22472));
    InMux I__5397 (
            .O(N__22477),
            .I(N__22472));
    LocalMux I__5396 (
            .O(N__22472),
            .I(N__22468));
    InMux I__5395 (
            .O(N__22471),
            .I(N__22465));
    Span4Mux_v I__5394 (
            .O(N__22468),
            .I(N__22460));
    LocalMux I__5393 (
            .O(N__22465),
            .I(N__22460));
    Span4Mux_h I__5392 (
            .O(N__22460),
            .I(N__22454));
    InMux I__5391 (
            .O(N__22459),
            .I(N__22451));
    InMux I__5390 (
            .O(N__22458),
            .I(N__22446));
    InMux I__5389 (
            .O(N__22457),
            .I(N__22446));
    Odrv4 I__5388 (
            .O(N__22454),
            .I(\c0.tx_transmit ));
    LocalMux I__5387 (
            .O(N__22451),
            .I(\c0.tx_transmit ));
    LocalMux I__5386 (
            .O(N__22446),
            .I(\c0.tx_transmit ));
    InMux I__5385 (
            .O(N__22439),
            .I(N__22435));
    InMux I__5384 (
            .O(N__22438),
            .I(N__22432));
    LocalMux I__5383 (
            .O(N__22435),
            .I(N__22428));
    LocalMux I__5382 (
            .O(N__22432),
            .I(N__22424));
    InMux I__5381 (
            .O(N__22431),
            .I(N__22421));
    Span4Mux_v I__5380 (
            .O(N__22428),
            .I(N__22418));
    InMux I__5379 (
            .O(N__22427),
            .I(N__22415));
    Span4Mux_v I__5378 (
            .O(N__22424),
            .I(N__22412));
    LocalMux I__5377 (
            .O(N__22421),
            .I(N__22409));
    Span4Mux_h I__5376 (
            .O(N__22418),
            .I(N__22406));
    LocalMux I__5375 (
            .O(N__22415),
            .I(N__22401));
    Span4Mux_h I__5374 (
            .O(N__22412),
            .I(N__22401));
    Span4Mux_v I__5373 (
            .O(N__22409),
            .I(N__22398));
    Odrv4 I__5372 (
            .O(N__22406),
            .I(data_out_field_0));
    Odrv4 I__5371 (
            .O(N__22401),
            .I(data_out_field_0));
    Odrv4 I__5370 (
            .O(N__22398),
            .I(data_out_field_0));
    InMux I__5369 (
            .O(N__22391),
            .I(N__22387));
    InMux I__5368 (
            .O(N__22390),
            .I(N__22384));
    LocalMux I__5367 (
            .O(N__22387),
            .I(\c0.n1421 ));
    LocalMux I__5366 (
            .O(N__22384),
            .I(\c0.n1421 ));
    InMux I__5365 (
            .O(N__22379),
            .I(N__22376));
    LocalMux I__5364 (
            .O(N__22376),
            .I(\c0.n1306 ));
    InMux I__5363 (
            .O(N__22373),
            .I(N__22370));
    LocalMux I__5362 (
            .O(N__22370),
            .I(N__22366));
    InMux I__5361 (
            .O(N__22369),
            .I(N__22363));
    Span4Mux_h I__5360 (
            .O(N__22366),
            .I(N__22360));
    LocalMux I__5359 (
            .O(N__22363),
            .I(\c0.n4453 ));
    Odrv4 I__5358 (
            .O(N__22360),
            .I(\c0.n4453 ));
    InMux I__5357 (
            .O(N__22355),
            .I(N__22352));
    LocalMux I__5356 (
            .O(N__22352),
            .I(N__22349));
    Span4Mux_h I__5355 (
            .O(N__22349),
            .I(N__22345));
    InMux I__5354 (
            .O(N__22348),
            .I(N__22342));
    Odrv4 I__5353 (
            .O(N__22345),
            .I(\c0.n1312 ));
    LocalMux I__5352 (
            .O(N__22342),
            .I(\c0.n1312 ));
    CascadeMux I__5351 (
            .O(N__22337),
            .I(\c0.n1306_cascade_ ));
    InMux I__5350 (
            .O(N__22334),
            .I(N__22331));
    LocalMux I__5349 (
            .O(N__22331),
            .I(N__22326));
    InMux I__5348 (
            .O(N__22330),
            .I(N__22319));
    InMux I__5347 (
            .O(N__22329),
            .I(N__22319));
    Span4Mux_v I__5346 (
            .O(N__22326),
            .I(N__22316));
    InMux I__5345 (
            .O(N__22325),
            .I(N__22311));
    InMux I__5344 (
            .O(N__22324),
            .I(N__22311));
    LocalMux I__5343 (
            .O(N__22319),
            .I(N__22308));
    Odrv4 I__5342 (
            .O(N__22316),
            .I(\c0.data_out_field_47_N_682_47 ));
    LocalMux I__5341 (
            .O(N__22311),
            .I(\c0.data_out_field_47_N_682_47 ));
    Odrv4 I__5340 (
            .O(N__22308),
            .I(\c0.data_out_field_47_N_682_47 ));
    CascadeMux I__5339 (
            .O(N__22301),
            .I(N__22298));
    InMux I__5338 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__5337 (
            .O(N__22295),
            .I(N__22292));
    Odrv12 I__5336 (
            .O(N__22292),
            .I(n4454));
    InMux I__5335 (
            .O(N__22289),
            .I(N__22286));
    LocalMux I__5334 (
            .O(N__22286),
            .I(\c0.tx_active_prev ));
    InMux I__5333 (
            .O(N__22283),
            .I(N__22280));
    LocalMux I__5332 (
            .O(N__22280),
            .I(\c0.n50 ));
    CascadeMux I__5331 (
            .O(N__22277),
            .I(\c0.tx.n2908_cascade_ ));
    CascadeMux I__5330 (
            .O(N__22274),
            .I(\c0.tx.n1457_cascade_ ));
    InMux I__5329 (
            .O(N__22271),
            .I(N__22266));
    InMux I__5328 (
            .O(N__22270),
            .I(N__22261));
    InMux I__5327 (
            .O(N__22269),
            .I(N__22261));
    LocalMux I__5326 (
            .O(N__22266),
            .I(N__22258));
    LocalMux I__5325 (
            .O(N__22261),
            .I(N__22255));
    Span4Mux_v I__5324 (
            .O(N__22258),
            .I(N__22249));
    Span4Mux_h I__5323 (
            .O(N__22255),
            .I(N__22246));
    InMux I__5322 (
            .O(N__22254),
            .I(N__22239));
    InMux I__5321 (
            .O(N__22253),
            .I(N__22239));
    InMux I__5320 (
            .O(N__22252),
            .I(N__22239));
    Odrv4 I__5319 (
            .O(N__22249),
            .I(\c0.tx_active ));
    Odrv4 I__5318 (
            .O(N__22246),
            .I(\c0.tx_active ));
    LocalMux I__5317 (
            .O(N__22239),
            .I(\c0.tx_active ));
    InMux I__5316 (
            .O(N__22232),
            .I(N__22228));
    InMux I__5315 (
            .O(N__22231),
            .I(N__22225));
    LocalMux I__5314 (
            .O(N__22228),
            .I(N__22222));
    LocalMux I__5313 (
            .O(N__22225),
            .I(N__22218));
    Span4Mux_v I__5312 (
            .O(N__22222),
            .I(N__22215));
    InMux I__5311 (
            .O(N__22221),
            .I(N__22211));
    Span4Mux_h I__5310 (
            .O(N__22218),
            .I(N__22208));
    Span4Mux_h I__5309 (
            .O(N__22215),
            .I(N__22205));
    InMux I__5308 (
            .O(N__22214),
            .I(N__22202));
    LocalMux I__5307 (
            .O(N__22211),
            .I(data_out_field_8));
    Odrv4 I__5306 (
            .O(N__22208),
            .I(data_out_field_8));
    Odrv4 I__5305 (
            .O(N__22205),
            .I(data_out_field_8));
    LocalMux I__5304 (
            .O(N__22202),
            .I(data_out_field_8));
    InMux I__5303 (
            .O(N__22193),
            .I(N__22188));
    InMux I__5302 (
            .O(N__22192),
            .I(N__22184));
    InMux I__5301 (
            .O(N__22191),
            .I(N__22181));
    LocalMux I__5300 (
            .O(N__22188),
            .I(N__22178));
    InMux I__5299 (
            .O(N__22187),
            .I(N__22175));
    LocalMux I__5298 (
            .O(N__22184),
            .I(data_out_field_23));
    LocalMux I__5297 (
            .O(N__22181),
            .I(data_out_field_23));
    Odrv4 I__5296 (
            .O(N__22178),
            .I(data_out_field_23));
    LocalMux I__5295 (
            .O(N__22175),
            .I(data_out_field_23));
    InMux I__5294 (
            .O(N__22166),
            .I(N__22163));
    LocalMux I__5293 (
            .O(N__22163),
            .I(N__22159));
    InMux I__5292 (
            .O(N__22162),
            .I(N__22156));
    Odrv4 I__5291 (
            .O(N__22159),
            .I(n1325));
    LocalMux I__5290 (
            .O(N__22156),
            .I(n1325));
    InMux I__5289 (
            .O(N__22151),
            .I(N__22147));
    InMux I__5288 (
            .O(N__22150),
            .I(N__22144));
    LocalMux I__5287 (
            .O(N__22147),
            .I(N__22138));
    LocalMux I__5286 (
            .O(N__22144),
            .I(N__22135));
    InMux I__5285 (
            .O(N__22143),
            .I(N__22132));
    InMux I__5284 (
            .O(N__22142),
            .I(N__22127));
    InMux I__5283 (
            .O(N__22141),
            .I(N__22127));
    Span4Mux_v I__5282 (
            .O(N__22138),
            .I(N__22120));
    Span4Mux_h I__5281 (
            .O(N__22135),
            .I(N__22120));
    LocalMux I__5280 (
            .O(N__22132),
            .I(N__22120));
    LocalMux I__5279 (
            .O(N__22127),
            .I(N__22117));
    Span4Mux_v I__5278 (
            .O(N__22120),
            .I(N__22109));
    Span4Mux_v I__5277 (
            .O(N__22117),
            .I(N__22109));
    InMux I__5276 (
            .O(N__22116),
            .I(N__22106));
    InMux I__5275 (
            .O(N__22115),
            .I(N__22101));
    InMux I__5274 (
            .O(N__22114),
            .I(N__22101));
    Span4Mux_h I__5273 (
            .O(N__22109),
            .I(N__22098));
    LocalMux I__5272 (
            .O(N__22106),
            .I(N__22093));
    LocalMux I__5271 (
            .O(N__22101),
            .I(N__22093));
    Odrv4 I__5270 (
            .O(N__22098),
            .I(n1025));
    Odrv12 I__5269 (
            .O(N__22093),
            .I(n1025));
    InMux I__5268 (
            .O(N__22088),
            .I(N__22085));
    LocalMux I__5267 (
            .O(N__22085),
            .I(\c0.tx.n752 ));
    InMux I__5266 (
            .O(N__22082),
            .I(N__22078));
    InMux I__5265 (
            .O(N__22081),
            .I(N__22075));
    LocalMux I__5264 (
            .O(N__22078),
            .I(N__22072));
    LocalMux I__5263 (
            .O(N__22075),
            .I(n4423));
    Odrv4 I__5262 (
            .O(N__22072),
            .I(n4423));
    CascadeMux I__5261 (
            .O(N__22067),
            .I(N__22064));
    InMux I__5260 (
            .O(N__22064),
            .I(N__22060));
    InMux I__5259 (
            .O(N__22063),
            .I(N__22057));
    LocalMux I__5258 (
            .O(N__22060),
            .I(N__22054));
    LocalMux I__5257 (
            .O(N__22057),
            .I(N__22051));
    Span4Mux_h I__5256 (
            .O(N__22054),
            .I(N__22048));
    Odrv4 I__5255 (
            .O(N__22051),
            .I(n4462));
    Odrv4 I__5254 (
            .O(N__22048),
            .I(n4462));
    InMux I__5253 (
            .O(N__22043),
            .I(N__22039));
    InMux I__5252 (
            .O(N__22042),
            .I(N__22035));
    LocalMux I__5251 (
            .O(N__22039),
            .I(N__22032));
    InMux I__5250 (
            .O(N__22038),
            .I(N__22028));
    LocalMux I__5249 (
            .O(N__22035),
            .I(N__22023));
    Span4Mux_v I__5248 (
            .O(N__22032),
            .I(N__22023));
    InMux I__5247 (
            .O(N__22031),
            .I(N__22020));
    LocalMux I__5246 (
            .O(N__22028),
            .I(N__22017));
    Odrv4 I__5245 (
            .O(N__22023),
            .I(data_out_field_26));
    LocalMux I__5244 (
            .O(N__22020),
            .I(data_out_field_26));
    Odrv12 I__5243 (
            .O(N__22017),
            .I(data_out_field_26));
    CascadeMux I__5242 (
            .O(N__22010),
            .I(N__22007));
    InMux I__5241 (
            .O(N__22007),
            .I(N__22004));
    LocalMux I__5240 (
            .O(N__22004),
            .I(n4655));
    InMux I__5239 (
            .O(N__22001),
            .I(N__21997));
    CascadeMux I__5238 (
            .O(N__22000),
            .I(N__21993));
    LocalMux I__5237 (
            .O(N__21997),
            .I(N__21987));
    InMux I__5236 (
            .O(N__21996),
            .I(N__21982));
    InMux I__5235 (
            .O(N__21993),
            .I(N__21982));
    InMux I__5234 (
            .O(N__21992),
            .I(N__21979));
    InMux I__5233 (
            .O(N__21991),
            .I(N__21976));
    InMux I__5232 (
            .O(N__21990),
            .I(N__21973));
    Span12Mux_s10_h I__5231 (
            .O(N__21987),
            .I(N__21970));
    LocalMux I__5230 (
            .O(N__21982),
            .I(data_out_field_2));
    LocalMux I__5229 (
            .O(N__21979),
            .I(data_out_field_2));
    LocalMux I__5228 (
            .O(N__21976),
            .I(data_out_field_2));
    LocalMux I__5227 (
            .O(N__21973),
            .I(data_out_field_2));
    Odrv12 I__5226 (
            .O(N__21970),
            .I(data_out_field_2));
    InMux I__5225 (
            .O(N__21959),
            .I(N__21951));
    InMux I__5224 (
            .O(N__21958),
            .I(N__21951));
    InMux I__5223 (
            .O(N__21957),
            .I(N__21948));
    InMux I__5222 (
            .O(N__21956),
            .I(N__21945));
    LocalMux I__5221 (
            .O(N__21951),
            .I(N__21940));
    LocalMux I__5220 (
            .O(N__21948),
            .I(N__21940));
    LocalMux I__5219 (
            .O(N__21945),
            .I(data_out_field_43));
    Odrv12 I__5218 (
            .O(N__21940),
            .I(data_out_field_43));
    CascadeMux I__5217 (
            .O(N__21935),
            .I(N__21932));
    InMux I__5216 (
            .O(N__21932),
            .I(N__21928));
    CascadeMux I__5215 (
            .O(N__21931),
            .I(N__21925));
    LocalMux I__5214 (
            .O(N__21928),
            .I(N__21922));
    InMux I__5213 (
            .O(N__21925),
            .I(N__21919));
    Span4Mux_h I__5212 (
            .O(N__21922),
            .I(N__21912));
    LocalMux I__5211 (
            .O(N__21919),
            .I(N__21912));
    InMux I__5210 (
            .O(N__21918),
            .I(N__21909));
    InMux I__5209 (
            .O(N__21917),
            .I(N__21906));
    Span4Mux_h I__5208 (
            .O(N__21912),
            .I(N__21903));
    LocalMux I__5207 (
            .O(N__21909),
            .I(N__21900));
    LocalMux I__5206 (
            .O(N__21906),
            .I(data_out_field_15));
    Odrv4 I__5205 (
            .O(N__21903),
            .I(data_out_field_15));
    Odrv4 I__5204 (
            .O(N__21900),
            .I(data_out_field_15));
    InMux I__5203 (
            .O(N__21893),
            .I(N__21886));
    InMux I__5202 (
            .O(N__21892),
            .I(N__21879));
    InMux I__5201 (
            .O(N__21891),
            .I(N__21879));
    InMux I__5200 (
            .O(N__21890),
            .I(N__21879));
    InMux I__5199 (
            .O(N__21889),
            .I(N__21876));
    LocalMux I__5198 (
            .O(N__21886),
            .I(N__21873));
    LocalMux I__5197 (
            .O(N__21879),
            .I(N__21867));
    LocalMux I__5196 (
            .O(N__21876),
            .I(N__21867));
    Span4Mux_h I__5195 (
            .O(N__21873),
            .I(N__21864));
    InMux I__5194 (
            .O(N__21872),
            .I(N__21861));
    Odrv4 I__5193 (
            .O(N__21867),
            .I(data_out_field_30));
    Odrv4 I__5192 (
            .O(N__21864),
            .I(data_out_field_30));
    LocalMux I__5191 (
            .O(N__21861),
            .I(data_out_field_30));
    InMux I__5190 (
            .O(N__21854),
            .I(N__21847));
    InMux I__5189 (
            .O(N__21853),
            .I(N__21847));
    InMux I__5188 (
            .O(N__21852),
            .I(N__21844));
    LocalMux I__5187 (
            .O(N__21847),
            .I(N__21841));
    LocalMux I__5186 (
            .O(N__21844),
            .I(N__21838));
    Span4Mux_h I__5185 (
            .O(N__21841),
            .I(N__21835));
    Span4Mux_h I__5184 (
            .O(N__21838),
            .I(N__21832));
    Span4Mux_h I__5183 (
            .O(N__21835),
            .I(N__21829));
    Odrv4 I__5182 (
            .O(N__21832),
            .I(\c0.tx.n1514 ));
    Odrv4 I__5181 (
            .O(N__21829),
            .I(\c0.tx.n1514 ));
    InMux I__5180 (
            .O(N__21824),
            .I(N__21819));
    InMux I__5179 (
            .O(N__21823),
            .I(N__21816));
    InMux I__5178 (
            .O(N__21822),
            .I(N__21811));
    LocalMux I__5177 (
            .O(N__21819),
            .I(N__21808));
    LocalMux I__5176 (
            .O(N__21816),
            .I(N__21805));
    InMux I__5175 (
            .O(N__21815),
            .I(N__21802));
    InMux I__5174 (
            .O(N__21814),
            .I(N__21799));
    LocalMux I__5173 (
            .O(N__21811),
            .I(N__21796));
    Span4Mux_h I__5172 (
            .O(N__21808),
            .I(N__21793));
    Span4Mux_h I__5171 (
            .O(N__21805),
            .I(N__21788));
    LocalMux I__5170 (
            .O(N__21802),
            .I(N__21788));
    LocalMux I__5169 (
            .O(N__21799),
            .I(data_out_field_38));
    Odrv12 I__5168 (
            .O(N__21796),
            .I(data_out_field_38));
    Odrv4 I__5167 (
            .O(N__21793),
            .I(data_out_field_38));
    Odrv4 I__5166 (
            .O(N__21788),
            .I(data_out_field_38));
    CascadeMux I__5165 (
            .O(N__21779),
            .I(N__21776));
    InMux I__5164 (
            .O(N__21776),
            .I(N__21772));
    InMux I__5163 (
            .O(N__21775),
            .I(N__21769));
    LocalMux I__5162 (
            .O(N__21772),
            .I(N__21764));
    LocalMux I__5161 (
            .O(N__21769),
            .I(N__21761));
    InMux I__5160 (
            .O(N__21768),
            .I(N__21758));
    InMux I__5159 (
            .O(N__21767),
            .I(N__21755));
    Span4Mux_h I__5158 (
            .O(N__21764),
            .I(N__21752));
    Span4Mux_v I__5157 (
            .O(N__21761),
            .I(N__21749));
    LocalMux I__5156 (
            .O(N__21758),
            .I(data_out_field_9));
    LocalMux I__5155 (
            .O(N__21755),
            .I(data_out_field_9));
    Odrv4 I__5154 (
            .O(N__21752),
            .I(data_out_field_9));
    Odrv4 I__5153 (
            .O(N__21749),
            .I(data_out_field_9));
    CascadeMux I__5152 (
            .O(N__21740),
            .I(N__21737));
    InMux I__5151 (
            .O(N__21737),
            .I(N__21732));
    InMux I__5150 (
            .O(N__21736),
            .I(N__21729));
    CascadeMux I__5149 (
            .O(N__21735),
            .I(N__21725));
    LocalMux I__5148 (
            .O(N__21732),
            .I(N__21721));
    LocalMux I__5147 (
            .O(N__21729),
            .I(N__21718));
    InMux I__5146 (
            .O(N__21728),
            .I(N__21715));
    InMux I__5145 (
            .O(N__21725),
            .I(N__21710));
    InMux I__5144 (
            .O(N__21724),
            .I(N__21710));
    Span4Mux_v I__5143 (
            .O(N__21721),
            .I(N__21707));
    Span4Mux_h I__5142 (
            .O(N__21718),
            .I(N__21704));
    LocalMux I__5141 (
            .O(N__21715),
            .I(N__21701));
    LocalMux I__5140 (
            .O(N__21710),
            .I(\c0.data_out_field_47_N_682_39 ));
    Odrv4 I__5139 (
            .O(N__21707),
            .I(\c0.data_out_field_47_N_682_39 ));
    Odrv4 I__5138 (
            .O(N__21704),
            .I(\c0.data_out_field_47_N_682_39 ));
    Odrv12 I__5137 (
            .O(N__21701),
            .I(\c0.data_out_field_47_N_682_39 ));
    InMux I__5136 (
            .O(N__21692),
            .I(N__21689));
    LocalMux I__5135 (
            .O(N__21689),
            .I(N__21686));
    Odrv12 I__5134 (
            .O(N__21686),
            .I(n4426));
    CascadeMux I__5133 (
            .O(N__21683),
            .I(n4426_cascade_));
    InMux I__5132 (
            .O(N__21680),
            .I(N__21677));
    LocalMux I__5131 (
            .O(N__21677),
            .I(N__21673));
    InMux I__5130 (
            .O(N__21676),
            .I(N__21668));
    Span4Mux_v I__5129 (
            .O(N__21673),
            .I(N__21665));
    InMux I__5128 (
            .O(N__21672),
            .I(N__21662));
    InMux I__5127 (
            .O(N__21671),
            .I(N__21659));
    LocalMux I__5126 (
            .O(N__21668),
            .I(N__21656));
    Span4Mux_h I__5125 (
            .O(N__21665),
            .I(N__21651));
    LocalMux I__5124 (
            .O(N__21662),
            .I(N__21651));
    LocalMux I__5123 (
            .O(N__21659),
            .I(data_out_field_10));
    Odrv4 I__5122 (
            .O(N__21656),
            .I(data_out_field_10));
    Odrv4 I__5121 (
            .O(N__21651),
            .I(data_out_field_10));
    InMux I__5120 (
            .O(N__21644),
            .I(N__21641));
    LocalMux I__5119 (
            .O(N__21641),
            .I(N__21638));
    Span4Mux_h I__5118 (
            .O(N__21638),
            .I(N__21635));
    Odrv4 I__5117 (
            .O(N__21635),
            .I(n4659));
    CascadeMux I__5116 (
            .O(N__21632),
            .I(N__21629));
    InMux I__5115 (
            .O(N__21629),
            .I(N__21626));
    LocalMux I__5114 (
            .O(N__21626),
            .I(N__21623));
    Span4Mux_v I__5113 (
            .O(N__21623),
            .I(N__21620));
    Span4Mux_h I__5112 (
            .O(N__21620),
            .I(N__21616));
    InMux I__5111 (
            .O(N__21619),
            .I(N__21613));
    Odrv4 I__5110 (
            .O(N__21616),
            .I(\c0.data_13 ));
    LocalMux I__5109 (
            .O(N__21613),
            .I(\c0.data_13 ));
    InMux I__5108 (
            .O(N__21608),
            .I(N__21603));
    InMux I__5107 (
            .O(N__21607),
            .I(N__21597));
    InMux I__5106 (
            .O(N__21606),
            .I(N__21597));
    LocalMux I__5105 (
            .O(N__21603),
            .I(N__21594));
    InMux I__5104 (
            .O(N__21602),
            .I(N__21591));
    LocalMux I__5103 (
            .O(N__21597),
            .I(\c0.data_out_field_47_N_682_37 ));
    Odrv4 I__5102 (
            .O(N__21594),
            .I(\c0.data_out_field_47_N_682_37 ));
    LocalMux I__5101 (
            .O(N__21591),
            .I(\c0.data_out_field_47_N_682_37 ));
    CascadeMux I__5100 (
            .O(N__21584),
            .I(N__21580));
    InMux I__5099 (
            .O(N__21583),
            .I(N__21565));
    InMux I__5098 (
            .O(N__21580),
            .I(N__21565));
    InMux I__5097 (
            .O(N__21579),
            .I(N__21565));
    InMux I__5096 (
            .O(N__21578),
            .I(N__21565));
    InMux I__5095 (
            .O(N__21577),
            .I(N__21565));
    InMux I__5094 (
            .O(N__21576),
            .I(N__21556));
    LocalMux I__5093 (
            .O(N__21565),
            .I(N__21551));
    InMux I__5092 (
            .O(N__21564),
            .I(N__21546));
    InMux I__5091 (
            .O(N__21563),
            .I(N__21546));
    InMux I__5090 (
            .O(N__21562),
            .I(N__21533));
    InMux I__5089 (
            .O(N__21561),
            .I(N__21530));
    InMux I__5088 (
            .O(N__21560),
            .I(N__21527));
    InMux I__5087 (
            .O(N__21559),
            .I(N__21515));
    LocalMux I__5086 (
            .O(N__21556),
            .I(N__21512));
    InMux I__5085 (
            .O(N__21555),
            .I(N__21509));
    InMux I__5084 (
            .O(N__21554),
            .I(N__21506));
    Span4Mux_v I__5083 (
            .O(N__21551),
            .I(N__21501));
    LocalMux I__5082 (
            .O(N__21546),
            .I(N__21501));
    InMux I__5081 (
            .O(N__21545),
            .I(N__21490));
    InMux I__5080 (
            .O(N__21544),
            .I(N__21490));
    InMux I__5079 (
            .O(N__21543),
            .I(N__21490));
    InMux I__5078 (
            .O(N__21542),
            .I(N__21490));
    InMux I__5077 (
            .O(N__21541),
            .I(N__21490));
    InMux I__5076 (
            .O(N__21540),
            .I(N__21487));
    InMux I__5075 (
            .O(N__21539),
            .I(N__21476));
    InMux I__5074 (
            .O(N__21538),
            .I(N__21476));
    InMux I__5073 (
            .O(N__21537),
            .I(N__21476));
    InMux I__5072 (
            .O(N__21536),
            .I(N__21476));
    LocalMux I__5071 (
            .O(N__21533),
            .I(N__21473));
    LocalMux I__5070 (
            .O(N__21530),
            .I(N__21470));
    LocalMux I__5069 (
            .O(N__21527),
            .I(N__21467));
    CascadeMux I__5068 (
            .O(N__21526),
            .I(N__21459));
    InMux I__5067 (
            .O(N__21525),
            .I(N__21456));
    InMux I__5066 (
            .O(N__21524),
            .I(N__21453));
    InMux I__5065 (
            .O(N__21523),
            .I(N__21450));
    InMux I__5064 (
            .O(N__21522),
            .I(N__21430));
    InMux I__5063 (
            .O(N__21521),
            .I(N__21421));
    InMux I__5062 (
            .O(N__21520),
            .I(N__21421));
    InMux I__5061 (
            .O(N__21519),
            .I(N__21421));
    InMux I__5060 (
            .O(N__21518),
            .I(N__21421));
    LocalMux I__5059 (
            .O(N__21515),
            .I(N__21414));
    Span4Mux_h I__5058 (
            .O(N__21512),
            .I(N__21414));
    LocalMux I__5057 (
            .O(N__21509),
            .I(N__21414));
    LocalMux I__5056 (
            .O(N__21506),
            .I(N__21411));
    Span4Mux_h I__5055 (
            .O(N__21501),
            .I(N__21406));
    LocalMux I__5054 (
            .O(N__21490),
            .I(N__21406));
    LocalMux I__5053 (
            .O(N__21487),
            .I(N__21403));
    InMux I__5052 (
            .O(N__21486),
            .I(N__21398));
    InMux I__5051 (
            .O(N__21485),
            .I(N__21398));
    LocalMux I__5050 (
            .O(N__21476),
            .I(N__21389));
    Span4Mux_v I__5049 (
            .O(N__21473),
            .I(N__21389));
    Span4Mux_v I__5048 (
            .O(N__21470),
            .I(N__21389));
    Span4Mux_v I__5047 (
            .O(N__21467),
            .I(N__21389));
    InMux I__5046 (
            .O(N__21466),
            .I(N__21384));
    InMux I__5045 (
            .O(N__21465),
            .I(N__21384));
    InMux I__5044 (
            .O(N__21464),
            .I(N__21375));
    InMux I__5043 (
            .O(N__21463),
            .I(N__21375));
    InMux I__5042 (
            .O(N__21462),
            .I(N__21375));
    InMux I__5041 (
            .O(N__21459),
            .I(N__21375));
    LocalMux I__5040 (
            .O(N__21456),
            .I(N__21372));
    LocalMux I__5039 (
            .O(N__21453),
            .I(N__21369));
    LocalMux I__5038 (
            .O(N__21450),
            .I(N__21366));
    InMux I__5037 (
            .O(N__21449),
            .I(N__21361));
    InMux I__5036 (
            .O(N__21448),
            .I(N__21361));
    InMux I__5035 (
            .O(N__21447),
            .I(N__21358));
    InMux I__5034 (
            .O(N__21446),
            .I(N__21355));
    InMux I__5033 (
            .O(N__21445),
            .I(N__21352));
    InMux I__5032 (
            .O(N__21444),
            .I(N__21349));
    InMux I__5031 (
            .O(N__21443),
            .I(N__21338));
    InMux I__5030 (
            .O(N__21442),
            .I(N__21338));
    InMux I__5029 (
            .O(N__21441),
            .I(N__21338));
    InMux I__5028 (
            .O(N__21440),
            .I(N__21338));
    InMux I__5027 (
            .O(N__21439),
            .I(N__21338));
    InMux I__5026 (
            .O(N__21438),
            .I(N__21327));
    InMux I__5025 (
            .O(N__21437),
            .I(N__21327));
    InMux I__5024 (
            .O(N__21436),
            .I(N__21327));
    InMux I__5023 (
            .O(N__21435),
            .I(N__21327));
    InMux I__5022 (
            .O(N__21434),
            .I(N__21327));
    InMux I__5021 (
            .O(N__21433),
            .I(N__21324));
    LocalMux I__5020 (
            .O(N__21430),
            .I(N__21321));
    LocalMux I__5019 (
            .O(N__21421),
            .I(N__21318));
    Span4Mux_v I__5018 (
            .O(N__21414),
            .I(N__21315));
    Span4Mux_v I__5017 (
            .O(N__21411),
            .I(N__21312));
    Span4Mux_h I__5016 (
            .O(N__21406),
            .I(N__21307));
    Span4Mux_h I__5015 (
            .O(N__21403),
            .I(N__21307));
    LocalMux I__5014 (
            .O(N__21398),
            .I(N__21302));
    Span4Mux_h I__5013 (
            .O(N__21389),
            .I(N__21302));
    LocalMux I__5012 (
            .O(N__21384),
            .I(N__21289));
    LocalMux I__5011 (
            .O(N__21375),
            .I(N__21289));
    Span4Mux_h I__5010 (
            .O(N__21372),
            .I(N__21289));
    Span4Mux_v I__5009 (
            .O(N__21369),
            .I(N__21289));
    Span4Mux_v I__5008 (
            .O(N__21366),
            .I(N__21289));
    LocalMux I__5007 (
            .O(N__21361),
            .I(N__21289));
    LocalMux I__5006 (
            .O(N__21358),
            .I(n3580));
    LocalMux I__5005 (
            .O(N__21355),
            .I(n3580));
    LocalMux I__5004 (
            .O(N__21352),
            .I(n3580));
    LocalMux I__5003 (
            .O(N__21349),
            .I(n3580));
    LocalMux I__5002 (
            .O(N__21338),
            .I(n3580));
    LocalMux I__5001 (
            .O(N__21327),
            .I(n3580));
    LocalMux I__5000 (
            .O(N__21324),
            .I(n3580));
    Odrv4 I__4999 (
            .O(N__21321),
            .I(n3580));
    Odrv12 I__4998 (
            .O(N__21318),
            .I(n3580));
    Odrv4 I__4997 (
            .O(N__21315),
            .I(n3580));
    Odrv4 I__4996 (
            .O(N__21312),
            .I(n3580));
    Odrv4 I__4995 (
            .O(N__21307),
            .I(n3580));
    Odrv4 I__4994 (
            .O(N__21302),
            .I(n3580));
    Odrv4 I__4993 (
            .O(N__21289),
            .I(n3580));
    InMux I__4992 (
            .O(N__21260),
            .I(N__21252));
    InMux I__4991 (
            .O(N__21259),
            .I(N__21243));
    InMux I__4990 (
            .O(N__21258),
            .I(N__21239));
    InMux I__4989 (
            .O(N__21257),
            .I(N__21235));
    InMux I__4988 (
            .O(N__21256),
            .I(N__21229));
    InMux I__4987 (
            .O(N__21255),
            .I(N__21229));
    LocalMux I__4986 (
            .O(N__21252),
            .I(N__21226));
    InMux I__4985 (
            .O(N__21251),
            .I(N__21221));
    InMux I__4984 (
            .O(N__21250),
            .I(N__21221));
    InMux I__4983 (
            .O(N__21249),
            .I(N__21216));
    InMux I__4982 (
            .O(N__21248),
            .I(N__21208));
    InMux I__4981 (
            .O(N__21247),
            .I(N__21208));
    InMux I__4980 (
            .O(N__21246),
            .I(N__21205));
    LocalMux I__4979 (
            .O(N__21243),
            .I(N__21202));
    InMux I__4978 (
            .O(N__21242),
            .I(N__21199));
    LocalMux I__4977 (
            .O(N__21239),
            .I(N__21196));
    InMux I__4976 (
            .O(N__21238),
            .I(N__21193));
    LocalMux I__4975 (
            .O(N__21235),
            .I(N__21190));
    InMux I__4974 (
            .O(N__21234),
            .I(N__21187));
    LocalMux I__4973 (
            .O(N__21229),
            .I(N__21173));
    Span4Mux_h I__4972 (
            .O(N__21226),
            .I(N__21170));
    LocalMux I__4971 (
            .O(N__21221),
            .I(N__21167));
    InMux I__4970 (
            .O(N__21220),
            .I(N__21162));
    InMux I__4969 (
            .O(N__21219),
            .I(N__21162));
    LocalMux I__4968 (
            .O(N__21216),
            .I(N__21159));
    InMux I__4967 (
            .O(N__21215),
            .I(N__21154));
    InMux I__4966 (
            .O(N__21214),
            .I(N__21154));
    InMux I__4965 (
            .O(N__21213),
            .I(N__21128));
    LocalMux I__4964 (
            .O(N__21208),
            .I(N__21125));
    LocalMux I__4963 (
            .O(N__21205),
            .I(N__21114));
    Span4Mux_h I__4962 (
            .O(N__21202),
            .I(N__21114));
    LocalMux I__4961 (
            .O(N__21199),
            .I(N__21114));
    Span4Mux_v I__4960 (
            .O(N__21196),
            .I(N__21114));
    LocalMux I__4959 (
            .O(N__21193),
            .I(N__21114));
    Span4Mux_h I__4958 (
            .O(N__21190),
            .I(N__21109));
    LocalMux I__4957 (
            .O(N__21187),
            .I(N__21109));
    InMux I__4956 (
            .O(N__21186),
            .I(N__21098));
    InMux I__4955 (
            .O(N__21185),
            .I(N__21098));
    InMux I__4954 (
            .O(N__21184),
            .I(N__21098));
    InMux I__4953 (
            .O(N__21183),
            .I(N__21098));
    InMux I__4952 (
            .O(N__21182),
            .I(N__21098));
    InMux I__4951 (
            .O(N__21181),
            .I(N__21093));
    InMux I__4950 (
            .O(N__21180),
            .I(N__21093));
    InMux I__4949 (
            .O(N__21179),
            .I(N__21084));
    InMux I__4948 (
            .O(N__21178),
            .I(N__21084));
    InMux I__4947 (
            .O(N__21177),
            .I(N__21084));
    InMux I__4946 (
            .O(N__21176),
            .I(N__21084));
    Span4Mux_h I__4945 (
            .O(N__21173),
            .I(N__21075));
    Span4Mux_v I__4944 (
            .O(N__21170),
            .I(N__21075));
    Span4Mux_v I__4943 (
            .O(N__21167),
            .I(N__21075));
    LocalMux I__4942 (
            .O(N__21162),
            .I(N__21075));
    Span4Mux_h I__4941 (
            .O(N__21159),
            .I(N__21070));
    LocalMux I__4940 (
            .O(N__21154),
            .I(N__21070));
    InMux I__4939 (
            .O(N__21153),
            .I(N__21059));
    InMux I__4938 (
            .O(N__21152),
            .I(N__21059));
    InMux I__4937 (
            .O(N__21151),
            .I(N__21059));
    InMux I__4936 (
            .O(N__21150),
            .I(N__21059));
    InMux I__4935 (
            .O(N__21149),
            .I(N__21059));
    InMux I__4934 (
            .O(N__21148),
            .I(N__21048));
    InMux I__4933 (
            .O(N__21147),
            .I(N__21048));
    InMux I__4932 (
            .O(N__21146),
            .I(N__21048));
    InMux I__4931 (
            .O(N__21145),
            .I(N__21048));
    InMux I__4930 (
            .O(N__21144),
            .I(N__21048));
    InMux I__4929 (
            .O(N__21143),
            .I(N__21041));
    InMux I__4928 (
            .O(N__21142),
            .I(N__21041));
    InMux I__4927 (
            .O(N__21141),
            .I(N__21041));
    InMux I__4926 (
            .O(N__21140),
            .I(N__21032));
    InMux I__4925 (
            .O(N__21139),
            .I(N__21032));
    InMux I__4924 (
            .O(N__21138),
            .I(N__21032));
    InMux I__4923 (
            .O(N__21137),
            .I(N__21032));
    InMux I__4922 (
            .O(N__21136),
            .I(N__21019));
    InMux I__4921 (
            .O(N__21135),
            .I(N__21019));
    InMux I__4920 (
            .O(N__21134),
            .I(N__21019));
    InMux I__4919 (
            .O(N__21133),
            .I(N__21019));
    InMux I__4918 (
            .O(N__21132),
            .I(N__21019));
    InMux I__4917 (
            .O(N__21131),
            .I(N__21019));
    LocalMux I__4916 (
            .O(N__21128),
            .I(n7_adj_938));
    Odrv4 I__4915 (
            .O(N__21125),
            .I(n7_adj_938));
    Odrv4 I__4914 (
            .O(N__21114),
            .I(n7_adj_938));
    Odrv4 I__4913 (
            .O(N__21109),
            .I(n7_adj_938));
    LocalMux I__4912 (
            .O(N__21098),
            .I(n7_adj_938));
    LocalMux I__4911 (
            .O(N__21093),
            .I(n7_adj_938));
    LocalMux I__4910 (
            .O(N__21084),
            .I(n7_adj_938));
    Odrv4 I__4909 (
            .O(N__21075),
            .I(n7_adj_938));
    Odrv4 I__4908 (
            .O(N__21070),
            .I(n7_adj_938));
    LocalMux I__4907 (
            .O(N__21059),
            .I(n7_adj_938));
    LocalMux I__4906 (
            .O(N__21048),
            .I(n7_adj_938));
    LocalMux I__4905 (
            .O(N__21041),
            .I(n7_adj_938));
    LocalMux I__4904 (
            .O(N__21032),
            .I(n7_adj_938));
    LocalMux I__4903 (
            .O(N__21019),
            .I(n7_adj_938));
    CascadeMux I__4902 (
            .O(N__20990),
            .I(N__20986));
    InMux I__4901 (
            .O(N__20989),
            .I(N__20981));
    InMux I__4900 (
            .O(N__20986),
            .I(N__20978));
    InMux I__4899 (
            .O(N__20985),
            .I(N__20975));
    InMux I__4898 (
            .O(N__20984),
            .I(N__20972));
    LocalMux I__4897 (
            .O(N__20981),
            .I(N__20969));
    LocalMux I__4896 (
            .O(N__20978),
            .I(N__20966));
    LocalMux I__4895 (
            .O(N__20975),
            .I(N__20963));
    LocalMux I__4894 (
            .O(N__20972),
            .I(data_out_field_1));
    Odrv4 I__4893 (
            .O(N__20969),
            .I(data_out_field_1));
    Odrv4 I__4892 (
            .O(N__20966),
            .I(data_out_field_1));
    Odrv4 I__4891 (
            .O(N__20963),
            .I(data_out_field_1));
    InMux I__4890 (
            .O(N__20954),
            .I(N__20951));
    LocalMux I__4889 (
            .O(N__20951),
            .I(N__20947));
    InMux I__4888 (
            .O(N__20950),
            .I(N__20943));
    Span4Mux_v I__4887 (
            .O(N__20947),
            .I(N__20940));
    InMux I__4886 (
            .O(N__20946),
            .I(N__20937));
    LocalMux I__4885 (
            .O(N__20943),
            .I(data_out_field_29));
    Odrv4 I__4884 (
            .O(N__20940),
            .I(data_out_field_29));
    LocalMux I__4883 (
            .O(N__20937),
            .I(data_out_field_29));
    InMux I__4882 (
            .O(N__20930),
            .I(N__20927));
    LocalMux I__4881 (
            .O(N__20927),
            .I(\c0.n4882 ));
    InMux I__4880 (
            .O(N__20924),
            .I(N__20917));
    InMux I__4879 (
            .O(N__20923),
            .I(N__20917));
    InMux I__4878 (
            .O(N__20922),
            .I(N__20914));
    LocalMux I__4877 (
            .O(N__20917),
            .I(N__20910));
    LocalMux I__4876 (
            .O(N__20914),
            .I(N__20907));
    InMux I__4875 (
            .O(N__20913),
            .I(N__20904));
    Span4Mux_v I__4874 (
            .O(N__20910),
            .I(N__20901));
    Span4Mux_h I__4873 (
            .O(N__20907),
            .I(N__20898));
    LocalMux I__4872 (
            .O(N__20904),
            .I(data_out_field_13));
    Odrv4 I__4871 (
            .O(N__20901),
            .I(data_out_field_13));
    Odrv4 I__4870 (
            .O(N__20898),
            .I(data_out_field_13));
    InMux I__4869 (
            .O(N__20891),
            .I(N__20887));
    InMux I__4868 (
            .O(N__20890),
            .I(N__20884));
    LocalMux I__4867 (
            .O(N__20887),
            .I(N__20879));
    LocalMux I__4866 (
            .O(N__20884),
            .I(N__20876));
    InMux I__4865 (
            .O(N__20883),
            .I(N__20873));
    InMux I__4864 (
            .O(N__20882),
            .I(N__20870));
    Span4Mux_s3_v I__4863 (
            .O(N__20879),
            .I(N__20865));
    Span4Mux_h I__4862 (
            .O(N__20876),
            .I(N__20865));
    LocalMux I__4861 (
            .O(N__20873),
            .I(data_out_field_28));
    LocalMux I__4860 (
            .O(N__20870),
            .I(data_out_field_28));
    Odrv4 I__4859 (
            .O(N__20865),
            .I(data_out_field_28));
    InMux I__4858 (
            .O(N__20858),
            .I(N__20853));
    InMux I__4857 (
            .O(N__20857),
            .I(N__20850));
    InMux I__4856 (
            .O(N__20856),
            .I(N__20846));
    LocalMux I__4855 (
            .O(N__20853),
            .I(N__20842));
    LocalMux I__4854 (
            .O(N__20850),
            .I(N__20839));
    InMux I__4853 (
            .O(N__20849),
            .I(N__20836));
    LocalMux I__4852 (
            .O(N__20846),
            .I(N__20833));
    InMux I__4851 (
            .O(N__20845),
            .I(N__20830));
    Span4Mux_v I__4850 (
            .O(N__20842),
            .I(N__20825));
    Span4Mux_h I__4849 (
            .O(N__20839),
            .I(N__20825));
    LocalMux I__4848 (
            .O(N__20836),
            .I(\c0.data_out_field_47_N_682_44 ));
    Odrv4 I__4847 (
            .O(N__20833),
            .I(\c0.data_out_field_47_N_682_44 ));
    LocalMux I__4846 (
            .O(N__20830),
            .I(\c0.data_out_field_47_N_682_44 ));
    Odrv4 I__4845 (
            .O(N__20825),
            .I(\c0.data_out_field_47_N_682_44 ));
    InMux I__4844 (
            .O(N__20816),
            .I(N__20813));
    LocalMux I__4843 (
            .O(N__20813),
            .I(N__20810));
    Span4Mux_h I__4842 (
            .O(N__20810),
            .I(N__20803));
    InMux I__4841 (
            .O(N__20809),
            .I(N__20800));
    InMux I__4840 (
            .O(N__20808),
            .I(N__20797));
    InMux I__4839 (
            .O(N__20807),
            .I(N__20792));
    InMux I__4838 (
            .O(N__20806),
            .I(N__20792));
    Odrv4 I__4837 (
            .O(N__20803),
            .I(\c0.data_out_field_47_N_682_36 ));
    LocalMux I__4836 (
            .O(N__20800),
            .I(\c0.data_out_field_47_N_682_36 ));
    LocalMux I__4835 (
            .O(N__20797),
            .I(\c0.data_out_field_47_N_682_36 ));
    LocalMux I__4834 (
            .O(N__20792),
            .I(\c0.data_out_field_47_N_682_36 ));
    InMux I__4833 (
            .O(N__20783),
            .I(N__20780));
    LocalMux I__4832 (
            .O(N__20780),
            .I(N__20777));
    Span4Mux_h I__4831 (
            .O(N__20777),
            .I(N__20774));
    Span4Mux_h I__4830 (
            .O(N__20774),
            .I(N__20771));
    Odrv4 I__4829 (
            .O(N__20771),
            .I(\c0.n4618 ));
    InMux I__4828 (
            .O(N__20768),
            .I(N__20765));
    LocalMux I__4827 (
            .O(N__20765),
            .I(N__20761));
    CascadeMux I__4826 (
            .O(N__20764),
            .I(N__20756));
    Span4Mux_v I__4825 (
            .O(N__20761),
            .I(N__20752));
    InMux I__4824 (
            .O(N__20760),
            .I(N__20749));
    InMux I__4823 (
            .O(N__20759),
            .I(N__20742));
    InMux I__4822 (
            .O(N__20756),
            .I(N__20742));
    InMux I__4821 (
            .O(N__20755),
            .I(N__20742));
    Odrv4 I__4820 (
            .O(N__20752),
            .I(data_out_field_21));
    LocalMux I__4819 (
            .O(N__20749),
            .I(data_out_field_21));
    LocalMux I__4818 (
            .O(N__20742),
            .I(data_out_field_21));
    CascadeMux I__4817 (
            .O(N__20735),
            .I(N__20732));
    InMux I__4816 (
            .O(N__20732),
            .I(N__20729));
    LocalMux I__4815 (
            .O(N__20729),
            .I(N__20726));
    Odrv4 I__4814 (
            .O(N__20726),
            .I(n1246));
    CascadeMux I__4813 (
            .O(N__20723),
            .I(N__20720));
    InMux I__4812 (
            .O(N__20720),
            .I(N__20717));
    LocalMux I__4811 (
            .O(N__20717),
            .I(N__20714));
    Span4Mux_h I__4810 (
            .O(N__20714),
            .I(N__20711));
    Odrv4 I__4809 (
            .O(N__20711),
            .I(n4663));
    InMux I__4808 (
            .O(N__20708),
            .I(N__20702));
    InMux I__4807 (
            .O(N__20707),
            .I(N__20698));
    InMux I__4806 (
            .O(N__20706),
            .I(N__20695));
    InMux I__4805 (
            .O(N__20705),
            .I(N__20690));
    LocalMux I__4804 (
            .O(N__20702),
            .I(N__20686));
    InMux I__4803 (
            .O(N__20701),
            .I(N__20683));
    LocalMux I__4802 (
            .O(N__20698),
            .I(N__20676));
    LocalMux I__4801 (
            .O(N__20695),
            .I(N__20673));
    InMux I__4800 (
            .O(N__20694),
            .I(N__20670));
    InMux I__4799 (
            .O(N__20693),
            .I(N__20667));
    LocalMux I__4798 (
            .O(N__20690),
            .I(N__20664));
    InMux I__4797 (
            .O(N__20689),
            .I(N__20661));
    Span4Mux_v I__4796 (
            .O(N__20686),
            .I(N__20655));
    LocalMux I__4795 (
            .O(N__20683),
            .I(N__20655));
    InMux I__4794 (
            .O(N__20682),
            .I(N__20650));
    InMux I__4793 (
            .O(N__20681),
            .I(N__20650));
    InMux I__4792 (
            .O(N__20680),
            .I(N__20645));
    InMux I__4791 (
            .O(N__20679),
            .I(N__20645));
    Span4Mux_v I__4790 (
            .O(N__20676),
            .I(N__20640));
    Span12Mux_s5_v I__4789 (
            .O(N__20673),
            .I(N__20633));
    LocalMux I__4788 (
            .O(N__20670),
            .I(N__20633));
    LocalMux I__4787 (
            .O(N__20667),
            .I(N__20633));
    Span4Mux_h I__4786 (
            .O(N__20664),
            .I(N__20628));
    LocalMux I__4785 (
            .O(N__20661),
            .I(N__20628));
    InMux I__4784 (
            .O(N__20660),
            .I(N__20625));
    Span4Mux_h I__4783 (
            .O(N__20655),
            .I(N__20620));
    LocalMux I__4782 (
            .O(N__20650),
            .I(N__20620));
    LocalMux I__4781 (
            .O(N__20645),
            .I(N__20617));
    InMux I__4780 (
            .O(N__20644),
            .I(N__20614));
    InMux I__4779 (
            .O(N__20643),
            .I(N__20611));
    Odrv4 I__4778 (
            .O(N__20640),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv12 I__4777 (
            .O(N__20633),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__4776 (
            .O(N__20628),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__4775 (
            .O(N__20625),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__4774 (
            .O(N__20620),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__4773 (
            .O(N__20617),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__4772 (
            .O(N__20614),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__4771 (
            .O(N__20611),
            .I(\c0.byte_transmit_counter_1 ));
    CascadeMux I__4770 (
            .O(N__20594),
            .I(N__20591));
    InMux I__4769 (
            .O(N__20591),
            .I(N__20587));
    CascadeMux I__4768 (
            .O(N__20590),
            .I(N__20584));
    LocalMux I__4767 (
            .O(N__20587),
            .I(N__20580));
    InMux I__4766 (
            .O(N__20584),
            .I(N__20575));
    InMux I__4765 (
            .O(N__20583),
            .I(N__20572));
    Span4Mux_h I__4764 (
            .O(N__20580),
            .I(N__20569));
    InMux I__4763 (
            .O(N__20579),
            .I(N__20564));
    InMux I__4762 (
            .O(N__20578),
            .I(N__20564));
    LocalMux I__4761 (
            .O(N__20575),
            .I(data_out_field_31));
    LocalMux I__4760 (
            .O(N__20572),
            .I(data_out_field_31));
    Odrv4 I__4759 (
            .O(N__20569),
            .I(data_out_field_31));
    LocalMux I__4758 (
            .O(N__20564),
            .I(data_out_field_31));
    InMux I__4757 (
            .O(N__20555),
            .I(N__20543));
    InMux I__4756 (
            .O(N__20554),
            .I(N__20540));
    InMux I__4755 (
            .O(N__20553),
            .I(N__20535));
    InMux I__4754 (
            .O(N__20552),
            .I(N__20535));
    InMux I__4753 (
            .O(N__20551),
            .I(N__20532));
    InMux I__4752 (
            .O(N__20550),
            .I(N__20527));
    InMux I__4751 (
            .O(N__20549),
            .I(N__20527));
    InMux I__4750 (
            .O(N__20548),
            .I(N__20520));
    InMux I__4749 (
            .O(N__20547),
            .I(N__20520));
    InMux I__4748 (
            .O(N__20546),
            .I(N__20520));
    LocalMux I__4747 (
            .O(N__20543),
            .I(N__20513));
    LocalMux I__4746 (
            .O(N__20540),
            .I(N__20502));
    LocalMux I__4745 (
            .O(N__20535),
            .I(N__20502));
    LocalMux I__4744 (
            .O(N__20532),
            .I(N__20502));
    LocalMux I__4743 (
            .O(N__20527),
            .I(N__20502));
    LocalMux I__4742 (
            .O(N__20520),
            .I(N__20502));
    InMux I__4741 (
            .O(N__20519),
            .I(N__20497));
    InMux I__4740 (
            .O(N__20518),
            .I(N__20497));
    CascadeMux I__4739 (
            .O(N__20517),
            .I(N__20490));
    InMux I__4738 (
            .O(N__20516),
            .I(N__20487));
    Span4Mux_s3_v I__4737 (
            .O(N__20513),
            .I(N__20480));
    Span4Mux_v I__4736 (
            .O(N__20502),
            .I(N__20480));
    LocalMux I__4735 (
            .O(N__20497),
            .I(N__20480));
    InMux I__4734 (
            .O(N__20496),
            .I(N__20472));
    InMux I__4733 (
            .O(N__20495),
            .I(N__20472));
    InMux I__4732 (
            .O(N__20494),
            .I(N__20467));
    InMux I__4731 (
            .O(N__20493),
            .I(N__20467));
    InMux I__4730 (
            .O(N__20490),
            .I(N__20462));
    LocalMux I__4729 (
            .O(N__20487),
            .I(N__20457));
    Span4Mux_h I__4728 (
            .O(N__20480),
            .I(N__20457));
    InMux I__4727 (
            .O(N__20479),
            .I(N__20454));
    InMux I__4726 (
            .O(N__20478),
            .I(N__20448));
    InMux I__4725 (
            .O(N__20477),
            .I(N__20445));
    LocalMux I__4724 (
            .O(N__20472),
            .I(N__20442));
    LocalMux I__4723 (
            .O(N__20467),
            .I(N__20439));
    InMux I__4722 (
            .O(N__20466),
            .I(N__20433));
    InMux I__4721 (
            .O(N__20465),
            .I(N__20433));
    LocalMux I__4720 (
            .O(N__20462),
            .I(N__20430));
    Span4Mux_h I__4719 (
            .O(N__20457),
            .I(N__20425));
    LocalMux I__4718 (
            .O(N__20454),
            .I(N__20425));
    CascadeMux I__4717 (
            .O(N__20453),
            .I(N__20420));
    InMux I__4716 (
            .O(N__20452),
            .I(N__20415));
    InMux I__4715 (
            .O(N__20451),
            .I(N__20415));
    LocalMux I__4714 (
            .O(N__20448),
            .I(N__20412));
    LocalMux I__4713 (
            .O(N__20445),
            .I(N__20409));
    Span4Mux_v I__4712 (
            .O(N__20442),
            .I(N__20404));
    Span4Mux_v I__4711 (
            .O(N__20439),
            .I(N__20404));
    InMux I__4710 (
            .O(N__20438),
            .I(N__20401));
    LocalMux I__4709 (
            .O(N__20433),
            .I(N__20394));
    Span4Mux_h I__4708 (
            .O(N__20430),
            .I(N__20394));
    Span4Mux_s3_v I__4707 (
            .O(N__20425),
            .I(N__20394));
    InMux I__4706 (
            .O(N__20424),
            .I(N__20389));
    InMux I__4705 (
            .O(N__20423),
            .I(N__20389));
    InMux I__4704 (
            .O(N__20420),
            .I(N__20386));
    LocalMux I__4703 (
            .O(N__20415),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__4702 (
            .O(N__20412),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__4701 (
            .O(N__20409),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__4700 (
            .O(N__20404),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__4699 (
            .O(N__20401),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__4698 (
            .O(N__20394),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__4697 (
            .O(N__20389),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__4696 (
            .O(N__20386),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__4695 (
            .O(N__20369),
            .I(N__20366));
    LocalMux I__4694 (
            .O(N__20366),
            .I(N__20363));
    Odrv12 I__4693 (
            .O(N__20363),
            .I(\c0.n4765 ));
    InMux I__4692 (
            .O(N__20360),
            .I(N__20355));
    InMux I__4691 (
            .O(N__20359),
            .I(N__20350));
    InMux I__4690 (
            .O(N__20358),
            .I(N__20350));
    LocalMux I__4689 (
            .O(N__20355),
            .I(data_out_field_14));
    LocalMux I__4688 (
            .O(N__20350),
            .I(data_out_field_14));
    CascadeMux I__4687 (
            .O(N__20345),
            .I(N__20342));
    InMux I__4686 (
            .O(N__20342),
            .I(N__20338));
    InMux I__4685 (
            .O(N__20341),
            .I(N__20335));
    LocalMux I__4684 (
            .O(N__20338),
            .I(N__20332));
    LocalMux I__4683 (
            .O(N__20335),
            .I(N__20329));
    Span4Mux_s3_v I__4682 (
            .O(N__20332),
            .I(N__20322));
    Span4Mux_h I__4681 (
            .O(N__20329),
            .I(N__20322));
    InMux I__4680 (
            .O(N__20328),
            .I(N__20319));
    InMux I__4679 (
            .O(N__20327),
            .I(N__20316));
    Span4Mux_v I__4678 (
            .O(N__20322),
            .I(N__20313));
    LocalMux I__4677 (
            .O(N__20319),
            .I(\c0.data_out_field_47_N_682_42 ));
    LocalMux I__4676 (
            .O(N__20316),
            .I(\c0.data_out_field_47_N_682_42 ));
    Odrv4 I__4675 (
            .O(N__20313),
            .I(\c0.data_out_field_47_N_682_42 ));
    CascadeMux I__4674 (
            .O(N__20306),
            .I(N__20303));
    InMux I__4673 (
            .O(N__20303),
            .I(N__20300));
    LocalMux I__4672 (
            .O(N__20300),
            .I(N__20296));
    InMux I__4671 (
            .O(N__20299),
            .I(N__20293));
    Odrv4 I__4670 (
            .O(N__20296),
            .I(n1255));
    LocalMux I__4669 (
            .O(N__20293),
            .I(n1255));
    InMux I__4668 (
            .O(N__20288),
            .I(N__20285));
    LocalMux I__4667 (
            .O(N__20285),
            .I(N__20281));
    InMux I__4666 (
            .O(N__20284),
            .I(N__20278));
    Span4Mux_h I__4665 (
            .O(N__20281),
            .I(N__20275));
    LocalMux I__4664 (
            .O(N__20278),
            .I(N__20272));
    Span4Mux_h I__4663 (
            .O(N__20275),
            .I(N__20269));
    Odrv4 I__4662 (
            .O(N__20272),
            .I(data_out_6_4));
    Odrv4 I__4661 (
            .O(N__20269),
            .I(data_out_6_4));
    CascadeMux I__4660 (
            .O(N__20264),
            .I(N__20259));
    InMux I__4659 (
            .O(N__20263),
            .I(N__20252));
    InMux I__4658 (
            .O(N__20262),
            .I(N__20252));
    InMux I__4657 (
            .O(N__20259),
            .I(N__20247));
    InMux I__4656 (
            .O(N__20258),
            .I(N__20247));
    InMux I__4655 (
            .O(N__20257),
            .I(N__20244));
    LocalMux I__4654 (
            .O(N__20252),
            .I(data_out_field_5));
    LocalMux I__4653 (
            .O(N__20247),
            .I(data_out_field_5));
    LocalMux I__4652 (
            .O(N__20244),
            .I(data_out_field_5));
    CascadeMux I__4651 (
            .O(N__20237),
            .I(N__20231));
    InMux I__4650 (
            .O(N__20236),
            .I(N__20228));
    InMux I__4649 (
            .O(N__20235),
            .I(N__20225));
    InMux I__4648 (
            .O(N__20234),
            .I(N__20221));
    InMux I__4647 (
            .O(N__20231),
            .I(N__20218));
    LocalMux I__4646 (
            .O(N__20228),
            .I(N__20215));
    LocalMux I__4645 (
            .O(N__20225),
            .I(N__20212));
    InMux I__4644 (
            .O(N__20224),
            .I(N__20209));
    LocalMux I__4643 (
            .O(N__20221),
            .I(data_out_field_18));
    LocalMux I__4642 (
            .O(N__20218),
            .I(data_out_field_18));
    Odrv4 I__4641 (
            .O(N__20215),
            .I(data_out_field_18));
    Odrv4 I__4640 (
            .O(N__20212),
            .I(data_out_field_18));
    LocalMux I__4639 (
            .O(N__20209),
            .I(data_out_field_18));
    InMux I__4638 (
            .O(N__20198),
            .I(N__20195));
    LocalMux I__4637 (
            .O(N__20195),
            .I(N__20189));
    InMux I__4636 (
            .O(N__20194),
            .I(N__20186));
    InMux I__4635 (
            .O(N__20193),
            .I(N__20182));
    InMux I__4634 (
            .O(N__20192),
            .I(N__20179));
    Span4Mux_h I__4633 (
            .O(N__20189),
            .I(N__20174));
    LocalMux I__4632 (
            .O(N__20186),
            .I(N__20174));
    InMux I__4631 (
            .O(N__20185),
            .I(N__20171));
    LocalMux I__4630 (
            .O(N__20182),
            .I(data_out_field_20));
    LocalMux I__4629 (
            .O(N__20179),
            .I(data_out_field_20));
    Odrv4 I__4628 (
            .O(N__20174),
            .I(data_out_field_20));
    LocalMux I__4627 (
            .O(N__20171),
            .I(data_out_field_20));
    InMux I__4626 (
            .O(N__20162),
            .I(N__20158));
    InMux I__4625 (
            .O(N__20161),
            .I(N__20155));
    LocalMux I__4624 (
            .O(N__20158),
            .I(N__20152));
    LocalMux I__4623 (
            .O(N__20155),
            .I(N__20147));
    Span4Mux_h I__4622 (
            .O(N__20152),
            .I(N__20144));
    InMux I__4621 (
            .O(N__20151),
            .I(N__20139));
    InMux I__4620 (
            .O(N__20150),
            .I(N__20139));
    Span4Mux_h I__4619 (
            .O(N__20147),
            .I(N__20136));
    Odrv4 I__4618 (
            .O(N__20144),
            .I(data_out_field_12));
    LocalMux I__4617 (
            .O(N__20139),
            .I(data_out_field_12));
    Odrv4 I__4616 (
            .O(N__20136),
            .I(data_out_field_12));
    CascadeMux I__4615 (
            .O(N__20129),
            .I(\c0.n4432_cascade_ ));
    InMux I__4614 (
            .O(N__20126),
            .I(N__20123));
    LocalMux I__4613 (
            .O(N__20123),
            .I(\c0.n4417 ));
    InMux I__4612 (
            .O(N__20120),
            .I(N__20117));
    LocalMux I__4611 (
            .O(N__20117),
            .I(N__20114));
    Odrv4 I__4610 (
            .O(N__20114),
            .I(\c0.n4483 ));
    CascadeMux I__4609 (
            .O(N__20111),
            .I(\c0.n10_adj_900_cascade_ ));
    InMux I__4608 (
            .O(N__20108),
            .I(N__20104));
    InMux I__4607 (
            .O(N__20107),
            .I(N__20101));
    LocalMux I__4606 (
            .O(N__20104),
            .I(N__20096));
    LocalMux I__4605 (
            .O(N__20101),
            .I(N__20096));
    Odrv4 I__4604 (
            .O(N__20096),
            .I(n4438));
    InMux I__4603 (
            .O(N__20093),
            .I(N__20087));
    InMux I__4602 (
            .O(N__20092),
            .I(N__20087));
    LocalMux I__4601 (
            .O(N__20087),
            .I(\c0.n4489 ));
    InMux I__4600 (
            .O(N__20084),
            .I(N__20081));
    LocalMux I__4599 (
            .O(N__20081),
            .I(N__20078));
    Odrv12 I__4598 (
            .O(N__20078),
            .I(\c0.n4532 ));
    CascadeMux I__4597 (
            .O(N__20075),
            .I(N__20071));
    CascadeMux I__4596 (
            .O(N__20074),
            .I(N__20067));
    InMux I__4595 (
            .O(N__20071),
            .I(N__20064));
    InMux I__4594 (
            .O(N__20070),
            .I(N__20050));
    InMux I__4593 (
            .O(N__20067),
            .I(N__20047));
    LocalMux I__4592 (
            .O(N__20064),
            .I(N__20044));
    InMux I__4591 (
            .O(N__20063),
            .I(N__20041));
    InMux I__4590 (
            .O(N__20062),
            .I(N__20038));
    InMux I__4589 (
            .O(N__20061),
            .I(N__20035));
    InMux I__4588 (
            .O(N__20060),
            .I(N__20030));
    InMux I__4587 (
            .O(N__20059),
            .I(N__20030));
    InMux I__4586 (
            .O(N__20058),
            .I(N__20025));
    InMux I__4585 (
            .O(N__20057),
            .I(N__20025));
    InMux I__4584 (
            .O(N__20056),
            .I(N__20022));
    InMux I__4583 (
            .O(N__20055),
            .I(N__20019));
    InMux I__4582 (
            .O(N__20054),
            .I(N__20014));
    InMux I__4581 (
            .O(N__20053),
            .I(N__20014));
    LocalMux I__4580 (
            .O(N__20050),
            .I(n1677));
    LocalMux I__4579 (
            .O(N__20047),
            .I(n1677));
    Odrv4 I__4578 (
            .O(N__20044),
            .I(n1677));
    LocalMux I__4577 (
            .O(N__20041),
            .I(n1677));
    LocalMux I__4576 (
            .O(N__20038),
            .I(n1677));
    LocalMux I__4575 (
            .O(N__20035),
            .I(n1677));
    LocalMux I__4574 (
            .O(N__20030),
            .I(n1677));
    LocalMux I__4573 (
            .O(N__20025),
            .I(n1677));
    LocalMux I__4572 (
            .O(N__20022),
            .I(n1677));
    LocalMux I__4571 (
            .O(N__20019),
            .I(n1677));
    LocalMux I__4570 (
            .O(N__20014),
            .I(n1677));
    InMux I__4569 (
            .O(N__19991),
            .I(N__19988));
    LocalMux I__4568 (
            .O(N__19988),
            .I(N__19985));
    Span4Mux_h I__4567 (
            .O(N__19985),
            .I(N__19979));
    InMux I__4566 (
            .O(N__19984),
            .I(N__19972));
    InMux I__4565 (
            .O(N__19983),
            .I(N__19972));
    InMux I__4564 (
            .O(N__19982),
            .I(N__19972));
    Odrv4 I__4563 (
            .O(N__19979),
            .I(\c0.n4465 ));
    LocalMux I__4562 (
            .O(N__19972),
            .I(\c0.n4465 ));
    InMux I__4561 (
            .O(N__19967),
            .I(N__19963));
    InMux I__4560 (
            .O(N__19966),
            .I(N__19960));
    LocalMux I__4559 (
            .O(N__19963),
            .I(\c0.data_out_7_5 ));
    LocalMux I__4558 (
            .O(N__19960),
            .I(\c0.data_out_7_5 ));
    CascadeMux I__4557 (
            .O(N__19955),
            .I(N__19950));
    CascadeMux I__4556 (
            .O(N__19954),
            .I(N__19947));
    InMux I__4555 (
            .O(N__19953),
            .I(N__19940));
    InMux I__4554 (
            .O(N__19950),
            .I(N__19940));
    InMux I__4553 (
            .O(N__19947),
            .I(N__19935));
    InMux I__4552 (
            .O(N__19946),
            .I(N__19935));
    InMux I__4551 (
            .O(N__19945),
            .I(N__19932));
    LocalMux I__4550 (
            .O(N__19940),
            .I(N__19927));
    LocalMux I__4549 (
            .O(N__19935),
            .I(N__19927));
    LocalMux I__4548 (
            .O(N__19932),
            .I(\c0.data_out_field_47_N_682_45 ));
    Odrv4 I__4547 (
            .O(N__19927),
            .I(\c0.data_out_field_47_N_682_45 ));
    InMux I__4546 (
            .O(N__19922),
            .I(N__19919));
    LocalMux I__4545 (
            .O(N__19919),
            .I(\c0.n4615 ));
    InMux I__4544 (
            .O(N__19916),
            .I(N__19912));
    InMux I__4543 (
            .O(N__19915),
            .I(N__19909));
    LocalMux I__4542 (
            .O(N__19912),
            .I(data_out_6_6));
    LocalMux I__4541 (
            .O(N__19909),
            .I(data_out_6_6));
    InMux I__4540 (
            .O(N__19904),
            .I(N__19900));
    InMux I__4539 (
            .O(N__19903),
            .I(N__19897));
    LocalMux I__4538 (
            .O(N__19900),
            .I(N__19894));
    LocalMux I__4537 (
            .O(N__19897),
            .I(data_out_7_6));
    Odrv4 I__4536 (
            .O(N__19894),
            .I(data_out_7_6));
    CascadeMux I__4535 (
            .O(N__19889),
            .I(\c0.n4879_cascade_ ));
    InMux I__4534 (
            .O(N__19886),
            .I(N__19882));
    InMux I__4533 (
            .O(N__19885),
            .I(N__19879));
    LocalMux I__4532 (
            .O(N__19882),
            .I(N__19873));
    LocalMux I__4531 (
            .O(N__19879),
            .I(N__19870));
    InMux I__4530 (
            .O(N__19878),
            .I(N__19867));
    InMux I__4529 (
            .O(N__19877),
            .I(N__19864));
    InMux I__4528 (
            .O(N__19876),
            .I(N__19861));
    Span4Mux_s3_v I__4527 (
            .O(N__19873),
            .I(N__19854));
    Span4Mux_h I__4526 (
            .O(N__19870),
            .I(N__19854));
    LocalMux I__4525 (
            .O(N__19867),
            .I(N__19854));
    LocalMux I__4524 (
            .O(N__19864),
            .I(\c0.data_out_field_47_N_682_46 ));
    LocalMux I__4523 (
            .O(N__19861),
            .I(\c0.data_out_field_47_N_682_46 ));
    Odrv4 I__4522 (
            .O(N__19854),
            .I(\c0.data_out_field_47_N_682_46 ));
    InMux I__4521 (
            .O(N__19847),
            .I(N__19844));
    LocalMux I__4520 (
            .O(N__19844),
            .I(N__19841));
    Span4Mux_h I__4519 (
            .O(N__19841),
            .I(N__19838));
    Span4Mux_h I__4518 (
            .O(N__19838),
            .I(N__19834));
    InMux I__4517 (
            .O(N__19837),
            .I(N__19831));
    Odrv4 I__4516 (
            .O(N__19834),
            .I(\c0.tx_transmit_N_274_7 ));
    LocalMux I__4515 (
            .O(N__19831),
            .I(\c0.tx_transmit_N_274_7 ));
    InMux I__4514 (
            .O(N__19826),
            .I(N__19823));
    LocalMux I__4513 (
            .O(N__19823),
            .I(N__19818));
    InMux I__4512 (
            .O(N__19822),
            .I(N__19814));
    InMux I__4511 (
            .O(N__19821),
            .I(N__19810));
    Span4Mux_h I__4510 (
            .O(N__19818),
            .I(N__19807));
    InMux I__4509 (
            .O(N__19817),
            .I(N__19804));
    LocalMux I__4508 (
            .O(N__19814),
            .I(N__19801));
    InMux I__4507 (
            .O(N__19813),
            .I(N__19798));
    LocalMux I__4506 (
            .O(N__19810),
            .I(\c0.data_out_field_47_N_682_35 ));
    Odrv4 I__4505 (
            .O(N__19807),
            .I(\c0.data_out_field_47_N_682_35 ));
    LocalMux I__4504 (
            .O(N__19804),
            .I(\c0.data_out_field_47_N_682_35 ));
    Odrv12 I__4503 (
            .O(N__19801),
            .I(\c0.data_out_field_47_N_682_35 ));
    LocalMux I__4502 (
            .O(N__19798),
            .I(\c0.data_out_field_47_N_682_35 ));
    InMux I__4501 (
            .O(N__19787),
            .I(N__19784));
    LocalMux I__4500 (
            .O(N__19784),
            .I(N__19781));
    Span4Mux_h I__4499 (
            .O(N__19781),
            .I(N__19778));
    Odrv4 I__4498 (
            .O(N__19778),
            .I(n10_adj_947));
    CascadeMux I__4497 (
            .O(N__19775),
            .I(n9_adj_948_cascade_));
    InMux I__4496 (
            .O(N__19772),
            .I(N__19769));
    LocalMux I__4495 (
            .O(N__19769),
            .I(N__19764));
    InMux I__4494 (
            .O(N__19768),
            .I(N__19759));
    InMux I__4493 (
            .O(N__19767),
            .I(N__19759));
    Span4Mux_h I__4492 (
            .O(N__19764),
            .I(N__19755));
    LocalMux I__4491 (
            .O(N__19759),
            .I(N__19752));
    InMux I__4490 (
            .O(N__19758),
            .I(N__19749));
    Span4Mux_h I__4489 (
            .O(N__19755),
            .I(N__19746));
    Span4Mux_v I__4488 (
            .O(N__19752),
            .I(N__19743));
    LocalMux I__4487 (
            .O(N__19749),
            .I(data_out_field_27));
    Odrv4 I__4486 (
            .O(N__19746),
            .I(data_out_field_27));
    Odrv4 I__4485 (
            .O(N__19743),
            .I(data_out_field_27));
    CascadeMux I__4484 (
            .O(N__19736),
            .I(N__19733));
    InMux I__4483 (
            .O(N__19733),
            .I(N__19730));
    LocalMux I__4482 (
            .O(N__19730),
            .I(N__19727));
    Span12Mux_h I__4481 (
            .O(N__19727),
            .I(N__19724));
    Odrv12 I__4480 (
            .O(N__19724),
            .I(n4_adj_942));
    CascadeMux I__4479 (
            .O(N__19721),
            .I(N__19718));
    InMux I__4478 (
            .O(N__19718),
            .I(N__19715));
    LocalMux I__4477 (
            .O(N__19715),
            .I(N__19712));
    Span4Mux_v I__4476 (
            .O(N__19712),
            .I(N__19709));
    Odrv4 I__4475 (
            .O(N__19709),
            .I(\c0.n4531 ));
    InMux I__4474 (
            .O(N__19706),
            .I(N__19703));
    LocalMux I__4473 (
            .O(N__19703),
            .I(N__19700));
    Odrv4 I__4472 (
            .O(N__19700),
            .I(n8_adj_968));
    InMux I__4471 (
            .O(N__19697),
            .I(N__19693));
    InMux I__4470 (
            .O(N__19696),
            .I(N__19690));
    LocalMux I__4469 (
            .O(N__19693),
            .I(data_out_7_0));
    LocalMux I__4468 (
            .O(N__19690),
            .I(data_out_7_0));
    InMux I__4467 (
            .O(N__19685),
            .I(N__19679));
    InMux I__4466 (
            .O(N__19684),
            .I(N__19679));
    LocalMux I__4465 (
            .O(N__19679),
            .I(data_out_6_0));
    CascadeMux I__4464 (
            .O(N__19676),
            .I(N__19673));
    InMux I__4463 (
            .O(N__19673),
            .I(N__19670));
    LocalMux I__4462 (
            .O(N__19670),
            .I(N__19667));
    Odrv12 I__4461 (
            .O(N__19667),
            .I(\c0.n4577 ));
    InMux I__4460 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__4459 (
            .O(N__19661),
            .I(N__19658));
    Span4Mux_h I__4458 (
            .O(N__19658),
            .I(N__19652));
    InMux I__4457 (
            .O(N__19657),
            .I(N__19649));
    InMux I__4456 (
            .O(N__19656),
            .I(N__19644));
    InMux I__4455 (
            .O(N__19655),
            .I(N__19644));
    Odrv4 I__4454 (
            .O(N__19652),
            .I(data_out_field_6));
    LocalMux I__4453 (
            .O(N__19649),
            .I(data_out_field_6));
    LocalMux I__4452 (
            .O(N__19644),
            .I(data_out_field_6));
    CascadeMux I__4451 (
            .O(N__19637),
            .I(n1246_cascade_));
    CascadeMux I__4450 (
            .O(N__19634),
            .I(N__19629));
    InMux I__4449 (
            .O(N__19633),
            .I(N__19625));
    InMux I__4448 (
            .O(N__19632),
            .I(N__19622));
    InMux I__4447 (
            .O(N__19629),
            .I(N__19619));
    InMux I__4446 (
            .O(N__19628),
            .I(N__19616));
    LocalMux I__4445 (
            .O(N__19625),
            .I(data_out_field_22));
    LocalMux I__4444 (
            .O(N__19622),
            .I(data_out_field_22));
    LocalMux I__4443 (
            .O(N__19619),
            .I(data_out_field_22));
    LocalMux I__4442 (
            .O(N__19616),
            .I(data_out_field_22));
    InMux I__4441 (
            .O(N__19607),
            .I(\c0.n3844 ));
    CascadeMux I__4440 (
            .O(N__19604),
            .I(N__19598));
    InMux I__4439 (
            .O(N__19603),
            .I(N__19591));
    InMux I__4438 (
            .O(N__19602),
            .I(N__19591));
    InMux I__4437 (
            .O(N__19601),
            .I(N__19586));
    InMux I__4436 (
            .O(N__19598),
            .I(N__19582));
    InMux I__4435 (
            .O(N__19597),
            .I(N__19577));
    InMux I__4434 (
            .O(N__19596),
            .I(N__19577));
    LocalMux I__4433 (
            .O(N__19591),
            .I(N__19574));
    InMux I__4432 (
            .O(N__19590),
            .I(N__19569));
    InMux I__4431 (
            .O(N__19589),
            .I(N__19569));
    LocalMux I__4430 (
            .O(N__19586),
            .I(N__19562));
    InMux I__4429 (
            .O(N__19585),
            .I(N__19558));
    LocalMux I__4428 (
            .O(N__19582),
            .I(N__19549));
    LocalMux I__4427 (
            .O(N__19577),
            .I(N__19549));
    Span4Mux_v I__4426 (
            .O(N__19574),
            .I(N__19549));
    LocalMux I__4425 (
            .O(N__19569),
            .I(N__19549));
    CascadeMux I__4424 (
            .O(N__19568),
            .I(N__19546));
    InMux I__4423 (
            .O(N__19567),
            .I(N__19541));
    InMux I__4422 (
            .O(N__19566),
            .I(N__19541));
    InMux I__4421 (
            .O(N__19565),
            .I(N__19538));
    Span4Mux_v I__4420 (
            .O(N__19562),
            .I(N__19535));
    InMux I__4419 (
            .O(N__19561),
            .I(N__19532));
    LocalMux I__4418 (
            .O(N__19558),
            .I(N__19529));
    Span4Mux_v I__4417 (
            .O(N__19549),
            .I(N__19526));
    InMux I__4416 (
            .O(N__19546),
            .I(N__19523));
    LocalMux I__4415 (
            .O(N__19541),
            .I(N__19517));
    LocalMux I__4414 (
            .O(N__19538),
            .I(N__19517));
    Span4Mux_h I__4413 (
            .O(N__19535),
            .I(N__19512));
    LocalMux I__4412 (
            .O(N__19532),
            .I(N__19512));
    Span4Mux_h I__4411 (
            .O(N__19529),
            .I(N__19505));
    Span4Mux_h I__4410 (
            .O(N__19526),
            .I(N__19505));
    LocalMux I__4409 (
            .O(N__19523),
            .I(N__19505));
    InMux I__4408 (
            .O(N__19522),
            .I(N__19502));
    Odrv12 I__4407 (
            .O(N__19517),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__4406 (
            .O(N__19512),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__4405 (
            .O(N__19505),
            .I(\c0.byte_transmit_counter_2 ));
    LocalMux I__4404 (
            .O(N__19502),
            .I(\c0.byte_transmit_counter_2 ));
    InMux I__4403 (
            .O(N__19493),
            .I(\c0.n3845 ));
    InMux I__4402 (
            .O(N__19490),
            .I(N__19487));
    LocalMux I__4401 (
            .O(N__19487),
            .I(\c0.byte_transmit_counter_3 ));
    InMux I__4400 (
            .O(N__19484),
            .I(N__19480));
    InMux I__4399 (
            .O(N__19483),
            .I(N__19477));
    LocalMux I__4398 (
            .O(N__19480),
            .I(\c0.tx_transmit_N_274_3 ));
    LocalMux I__4397 (
            .O(N__19477),
            .I(\c0.tx_transmit_N_274_3 ));
    InMux I__4396 (
            .O(N__19472),
            .I(\c0.n3846 ));
    InMux I__4395 (
            .O(N__19469),
            .I(N__19466));
    LocalMux I__4394 (
            .O(N__19466),
            .I(N__19463));
    Span12Mux_s7_v I__4393 (
            .O(N__19463),
            .I(N__19460));
    Odrv12 I__4392 (
            .O(N__19460),
            .I(\c0.byte_transmit_counter_4 ));
    InMux I__4391 (
            .O(N__19457),
            .I(N__19454));
    LocalMux I__4390 (
            .O(N__19454),
            .I(N__19451));
    Span4Mux_h I__4389 (
            .O(N__19451),
            .I(N__19448));
    Span4Mux_h I__4388 (
            .O(N__19448),
            .I(N__19444));
    InMux I__4387 (
            .O(N__19447),
            .I(N__19441));
    Odrv4 I__4386 (
            .O(N__19444),
            .I(\c0.tx_transmit_N_274_4 ));
    LocalMux I__4385 (
            .O(N__19441),
            .I(\c0.tx_transmit_N_274_4 ));
    InMux I__4384 (
            .O(N__19436),
            .I(\c0.n3847 ));
    InMux I__4383 (
            .O(N__19433),
            .I(N__19430));
    LocalMux I__4382 (
            .O(N__19430),
            .I(N__19427));
    Span4Mux_h I__4381 (
            .O(N__19427),
            .I(N__19424));
    Span4Mux_h I__4380 (
            .O(N__19424),
            .I(N__19421));
    Odrv4 I__4379 (
            .O(N__19421),
            .I(\c0.byte_transmit_counter_5 ));
    InMux I__4378 (
            .O(N__19418),
            .I(N__19415));
    LocalMux I__4377 (
            .O(N__19415),
            .I(N__19412));
    Span4Mux_h I__4376 (
            .O(N__19412),
            .I(N__19409));
    Span4Mux_h I__4375 (
            .O(N__19409),
            .I(N__19405));
    InMux I__4374 (
            .O(N__19408),
            .I(N__19402));
    Odrv4 I__4373 (
            .O(N__19405),
            .I(\c0.tx_transmit_N_274_5 ));
    LocalMux I__4372 (
            .O(N__19402),
            .I(\c0.tx_transmit_N_274_5 ));
    InMux I__4371 (
            .O(N__19397),
            .I(\c0.n3848 ));
    InMux I__4370 (
            .O(N__19394),
            .I(N__19391));
    LocalMux I__4369 (
            .O(N__19391),
            .I(N__19388));
    Span4Mux_h I__4368 (
            .O(N__19388),
            .I(N__19385));
    Span4Mux_h I__4367 (
            .O(N__19385),
            .I(N__19382));
    Odrv4 I__4366 (
            .O(N__19382),
            .I(\c0.byte_transmit_counter_6 ));
    InMux I__4365 (
            .O(N__19379),
            .I(N__19376));
    LocalMux I__4364 (
            .O(N__19376),
            .I(N__19373));
    Span4Mux_h I__4363 (
            .O(N__19373),
            .I(N__19370));
    Span4Mux_h I__4362 (
            .O(N__19370),
            .I(N__19366));
    InMux I__4361 (
            .O(N__19369),
            .I(N__19363));
    Odrv4 I__4360 (
            .O(N__19366),
            .I(\c0.tx_transmit_N_274_6 ));
    LocalMux I__4359 (
            .O(N__19363),
            .I(\c0.tx_transmit_N_274_6 ));
    InMux I__4358 (
            .O(N__19358),
            .I(\c0.n3849 ));
    InMux I__4357 (
            .O(N__19355),
            .I(N__19352));
    LocalMux I__4356 (
            .O(N__19352),
            .I(N__19349));
    Span4Mux_v I__4355 (
            .O(N__19349),
            .I(N__19346));
    Span4Mux_h I__4354 (
            .O(N__19346),
            .I(N__19343));
    Odrv4 I__4353 (
            .O(N__19343),
            .I(\c0.byte_transmit_counter_7 ));
    InMux I__4352 (
            .O(N__19340),
            .I(\c0.n3850 ));
    CascadeMux I__4351 (
            .O(N__19337),
            .I(\c0.n4774_cascade_ ));
    InMux I__4350 (
            .O(N__19334),
            .I(N__19331));
    LocalMux I__4349 (
            .O(N__19331),
            .I(N__19328));
    Span4Mux_v I__4348 (
            .O(N__19328),
            .I(N__19325));
    Odrv4 I__4347 (
            .O(N__19325),
            .I(tx_data_6_keep));
    CascadeMux I__4346 (
            .O(N__19322),
            .I(N__19319));
    InMux I__4345 (
            .O(N__19319),
            .I(N__19316));
    LocalMux I__4344 (
            .O(N__19316),
            .I(N__19313));
    Span4Mux_h I__4343 (
            .O(N__19313),
            .I(N__19310));
    Odrv4 I__4342 (
            .O(N__19310),
            .I(n10_adj_971));
    CascadeMux I__4341 (
            .O(N__19307),
            .I(N__19304));
    InMux I__4340 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__4339 (
            .O(N__19301),
            .I(N__19298));
    Span4Mux_h I__4338 (
            .O(N__19298),
            .I(N__19294));
    InMux I__4337 (
            .O(N__19297),
            .I(N__19291));
    Odrv4 I__4336 (
            .O(N__19294),
            .I(\c0.data_12 ));
    LocalMux I__4335 (
            .O(N__19291),
            .I(\c0.data_12 ));
    InMux I__4334 (
            .O(N__19286),
            .I(N__19282));
    CascadeMux I__4333 (
            .O(N__19285),
            .I(N__19278));
    LocalMux I__4332 (
            .O(N__19282),
            .I(N__19275));
    InMux I__4331 (
            .O(N__19281),
            .I(N__19270));
    InMux I__4330 (
            .O(N__19278),
            .I(N__19270));
    Odrv12 I__4329 (
            .O(N__19275),
            .I(data_out_field_7));
    LocalMux I__4328 (
            .O(N__19270),
            .I(data_out_field_7));
    InMux I__4327 (
            .O(N__19265),
            .I(N__19262));
    LocalMux I__4326 (
            .O(N__19262),
            .I(N__19258));
    CascadeMux I__4325 (
            .O(N__19261),
            .I(N__19253));
    Span4Mux_h I__4324 (
            .O(N__19258),
            .I(N__19250));
    InMux I__4323 (
            .O(N__19257),
            .I(N__19247));
    InMux I__4322 (
            .O(N__19256),
            .I(N__19242));
    InMux I__4321 (
            .O(N__19253),
            .I(N__19242));
    Odrv4 I__4320 (
            .O(N__19250),
            .I(\c0.tx.r_Bit_Index_2 ));
    LocalMux I__4319 (
            .O(N__19247),
            .I(\c0.tx.r_Bit_Index_2 ));
    LocalMux I__4318 (
            .O(N__19242),
            .I(\c0.tx.r_Bit_Index_2 ));
    InMux I__4317 (
            .O(N__19235),
            .I(N__19232));
    LocalMux I__4316 (
            .O(N__19232),
            .I(N__19229));
    Span12Mux_s3_v I__4315 (
            .O(N__19229),
            .I(N__19223));
    InMux I__4314 (
            .O(N__19228),
            .I(N__19216));
    InMux I__4313 (
            .O(N__19227),
            .I(N__19216));
    InMux I__4312 (
            .O(N__19226),
            .I(N__19216));
    Odrv12 I__4311 (
            .O(N__19223),
            .I(\c0.tx.r_Bit_Index_1 ));
    LocalMux I__4310 (
            .O(N__19216),
            .I(\c0.tx.r_Bit_Index_1 ));
    InMux I__4309 (
            .O(N__19211),
            .I(N__19203));
    CascadeMux I__4308 (
            .O(N__19210),
            .I(N__19200));
    InMux I__4307 (
            .O(N__19209),
            .I(N__19194));
    InMux I__4306 (
            .O(N__19208),
            .I(N__19194));
    InMux I__4305 (
            .O(N__19207),
            .I(N__19189));
    InMux I__4304 (
            .O(N__19206),
            .I(N__19189));
    LocalMux I__4303 (
            .O(N__19203),
            .I(N__19186));
    InMux I__4302 (
            .O(N__19200),
            .I(N__19182));
    InMux I__4301 (
            .O(N__19199),
            .I(N__19179));
    LocalMux I__4300 (
            .O(N__19194),
            .I(N__19172));
    LocalMux I__4299 (
            .O(N__19189),
            .I(N__19172));
    Span4Mux_h I__4298 (
            .O(N__19186),
            .I(N__19172));
    InMux I__4297 (
            .O(N__19185),
            .I(N__19169));
    LocalMux I__4296 (
            .O(N__19182),
            .I(\c0.tx.r_Bit_Index_0 ));
    LocalMux I__4295 (
            .O(N__19179),
            .I(\c0.tx.r_Bit_Index_0 ));
    Odrv4 I__4294 (
            .O(N__19172),
            .I(\c0.tx.r_Bit_Index_0 ));
    LocalMux I__4293 (
            .O(N__19169),
            .I(\c0.tx.r_Bit_Index_0 ));
    InMux I__4292 (
            .O(N__19160),
            .I(N__19156));
    InMux I__4291 (
            .O(N__19159),
            .I(N__19153));
    LocalMux I__4290 (
            .O(N__19156),
            .I(data_out_6_5));
    LocalMux I__4289 (
            .O(N__19153),
            .I(data_out_6_5));
    InMux I__4288 (
            .O(N__19148),
            .I(N__19145));
    LocalMux I__4287 (
            .O(N__19145),
            .I(\c0.n4616 ));
    InMux I__4286 (
            .O(N__19142),
            .I(N__19136));
    InMux I__4285 (
            .O(N__19141),
            .I(N__19133));
    InMux I__4284 (
            .O(N__19140),
            .I(N__19127));
    InMux I__4283 (
            .O(N__19139),
            .I(N__19127));
    LocalMux I__4282 (
            .O(N__19136),
            .I(N__19122));
    LocalMux I__4281 (
            .O(N__19133),
            .I(N__19122));
    InMux I__4280 (
            .O(N__19132),
            .I(N__19119));
    LocalMux I__4279 (
            .O(N__19127),
            .I(data_out_field_25));
    Odrv12 I__4278 (
            .O(N__19122),
            .I(data_out_field_25));
    LocalMux I__4277 (
            .O(N__19119),
            .I(data_out_field_25));
    InMux I__4276 (
            .O(N__19112),
            .I(N__19107));
    InMux I__4275 (
            .O(N__19111),
            .I(N__19102));
    InMux I__4274 (
            .O(N__19110),
            .I(N__19099));
    LocalMux I__4273 (
            .O(N__19107),
            .I(N__19096));
    InMux I__4272 (
            .O(N__19106),
            .I(N__19091));
    InMux I__4271 (
            .O(N__19105),
            .I(N__19091));
    LocalMux I__4270 (
            .O(N__19102),
            .I(\c0.data_out_field_47_N_682_40 ));
    LocalMux I__4269 (
            .O(N__19099),
            .I(\c0.data_out_field_47_N_682_40 ));
    Odrv4 I__4268 (
            .O(N__19096),
            .I(\c0.data_out_field_47_N_682_40 ));
    LocalMux I__4267 (
            .O(N__19091),
            .I(\c0.data_out_field_47_N_682_40 ));
    InMux I__4266 (
            .O(N__19082),
            .I(N__19079));
    LocalMux I__4265 (
            .O(N__19079),
            .I(N__19076));
    Span4Mux_v I__4264 (
            .O(N__19076),
            .I(N__19073));
    Span4Mux_h I__4263 (
            .O(N__19073),
            .I(N__19070));
    Odrv4 I__4262 (
            .O(N__19070),
            .I(\c0.n4561 ));
    CascadeMux I__4261 (
            .O(N__19067),
            .I(N__19064));
    InMux I__4260 (
            .O(N__19064),
            .I(N__19061));
    LocalMux I__4259 (
            .O(N__19061),
            .I(N__19057));
    InMux I__4258 (
            .O(N__19060),
            .I(N__19054));
    Odrv12 I__4257 (
            .O(N__19057),
            .I(\c0.data_2 ));
    LocalMux I__4256 (
            .O(N__19054),
            .I(\c0.data_2 ));
    CascadeMux I__4255 (
            .O(N__19049),
            .I(\c0.n4771_cascade_ ));
    InMux I__4254 (
            .O(N__19046),
            .I(N__19043));
    LocalMux I__4253 (
            .O(N__19043),
            .I(n7_adj_935));
    CascadeMux I__4252 (
            .O(N__19040),
            .I(n8_adj_934_cascade_));
    CascadeMux I__4251 (
            .O(N__19037),
            .I(N__19034));
    InMux I__4250 (
            .O(N__19034),
            .I(N__19030));
    InMux I__4249 (
            .O(N__19033),
            .I(N__19027));
    LocalMux I__4248 (
            .O(N__19030),
            .I(N__19024));
    LocalMux I__4247 (
            .O(N__19027),
            .I(data_out_7_7));
    Odrv4 I__4246 (
            .O(N__19024),
            .I(data_out_7_7));
    InMux I__4245 (
            .O(N__19019),
            .I(N__19016));
    LocalMux I__4244 (
            .O(N__19016),
            .I(N__19013));
    Span4Mux_h I__4243 (
            .O(N__19013),
            .I(N__19010));
    Odrv4 I__4242 (
            .O(N__19010),
            .I(\c0.n1333 ));
    CascadeMux I__4241 (
            .O(N__19007),
            .I(\c0.n4447_cascade_ ));
    InMux I__4240 (
            .O(N__19004),
            .I(N__19001));
    LocalMux I__4239 (
            .O(N__19001),
            .I(n9_adj_972));
    InMux I__4238 (
            .O(N__18998),
            .I(N__18995));
    LocalMux I__4237 (
            .O(N__18995),
            .I(N__18992));
    Odrv4 I__4236 (
            .O(N__18992),
            .I(\c0.n4795 ));
    InMux I__4235 (
            .O(N__18989),
            .I(N__18986));
    LocalMux I__4234 (
            .O(N__18986),
            .I(N__18983));
    Odrv4 I__4233 (
            .O(N__18983),
            .I(n11_adj_945));
    InMux I__4232 (
            .O(N__18980),
            .I(N__18977));
    LocalMux I__4231 (
            .O(N__18977),
            .I(N__18974));
    Span4Mux_v I__4230 (
            .O(N__18974),
            .I(N__18971));
    Odrv4 I__4229 (
            .O(N__18971),
            .I(n4_adj_970));
    InMux I__4228 (
            .O(N__18968),
            .I(N__18961));
    InMux I__4227 (
            .O(N__18967),
            .I(N__18958));
    InMux I__4226 (
            .O(N__18966),
            .I(N__18955));
    InMux I__4225 (
            .O(N__18965),
            .I(N__18952));
    InMux I__4224 (
            .O(N__18964),
            .I(N__18949));
    LocalMux I__4223 (
            .O(N__18961),
            .I(N__18946));
    LocalMux I__4222 (
            .O(N__18958),
            .I(data_out_field_16));
    LocalMux I__4221 (
            .O(N__18955),
            .I(data_out_field_16));
    LocalMux I__4220 (
            .O(N__18952),
            .I(data_out_field_16));
    LocalMux I__4219 (
            .O(N__18949),
            .I(data_out_field_16));
    Odrv4 I__4218 (
            .O(N__18946),
            .I(data_out_field_16));
    InMux I__4217 (
            .O(N__18935),
            .I(N__18932));
    LocalMux I__4216 (
            .O(N__18932),
            .I(\c0.n4447 ));
    CascadeMux I__4215 (
            .O(N__18929),
            .I(n7_adj_969_cascade_));
    InMux I__4214 (
            .O(N__18926),
            .I(N__18922));
    InMux I__4213 (
            .O(N__18925),
            .I(N__18919));
    LocalMux I__4212 (
            .O(N__18922),
            .I(N__18916));
    LocalMux I__4211 (
            .O(N__18919),
            .I(N__18913));
    Span4Mux_h I__4210 (
            .O(N__18916),
            .I(N__18910));
    Odrv12 I__4209 (
            .O(N__18913),
            .I(\c0.n4380 ));
    Odrv4 I__4208 (
            .O(N__18910),
            .I(\c0.n4380 ));
    InMux I__4207 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__4206 (
            .O(N__18902),
            .I(N__18898));
    InMux I__4205 (
            .O(N__18901),
            .I(N__18895));
    Span4Mux_v I__4204 (
            .O(N__18898),
            .I(N__18889));
    LocalMux I__4203 (
            .O(N__18895),
            .I(N__18889));
    InMux I__4202 (
            .O(N__18894),
            .I(N__18884));
    Span4Mux_h I__4201 (
            .O(N__18889),
            .I(N__18881));
    InMux I__4200 (
            .O(N__18888),
            .I(N__18878));
    InMux I__4199 (
            .O(N__18887),
            .I(N__18875));
    LocalMux I__4198 (
            .O(N__18884),
            .I(\c0.data_out_field_47_N_682_33 ));
    Odrv4 I__4197 (
            .O(N__18881),
            .I(\c0.data_out_field_47_N_682_33 ));
    LocalMux I__4196 (
            .O(N__18878),
            .I(\c0.data_out_field_47_N_682_33 ));
    LocalMux I__4195 (
            .O(N__18875),
            .I(\c0.data_out_field_47_N_682_33 ));
    CascadeMux I__4194 (
            .O(N__18866),
            .I(N__18863));
    InMux I__4193 (
            .O(N__18863),
            .I(N__18860));
    LocalMux I__4192 (
            .O(N__18860),
            .I(\c0.n4393 ));
    InMux I__4191 (
            .O(N__18857),
            .I(N__18854));
    LocalMux I__4190 (
            .O(N__18854),
            .I(N__18851));
    Odrv4 I__4189 (
            .O(N__18851),
            .I(n12_adj_966));
    CascadeMux I__4188 (
            .O(N__18848),
            .I(n1677_cascade_));
    InMux I__4187 (
            .O(N__18845),
            .I(N__18841));
    InMux I__4186 (
            .O(N__18844),
            .I(N__18838));
    LocalMux I__4185 (
            .O(N__18841),
            .I(N__18835));
    LocalMux I__4184 (
            .O(N__18838),
            .I(data_out_6_7));
    Odrv4 I__4183 (
            .O(N__18835),
            .I(data_out_6_7));
    CascadeMux I__4182 (
            .O(N__18830),
            .I(N__18827));
    InMux I__4181 (
            .O(N__18827),
            .I(N__18824));
    LocalMux I__4180 (
            .O(N__18824),
            .I(\c0.n4885 ));
    InMux I__4179 (
            .O(N__18821),
            .I(N__18818));
    LocalMux I__4178 (
            .O(N__18818),
            .I(N__18815));
    Span4Mux_h I__4177 (
            .O(N__18815),
            .I(N__18811));
    InMux I__4176 (
            .O(N__18814),
            .I(N__18808));
    Odrv4 I__4175 (
            .O(N__18811),
            .I(\c0.data_5 ));
    LocalMux I__4174 (
            .O(N__18808),
            .I(\c0.data_5 ));
    CascadeMux I__4173 (
            .O(N__18803),
            .I(\c0.n6_adj_904_cascade_ ));
    CascadeMux I__4172 (
            .O(N__18800),
            .I(n7_adj_938_cascade_));
    InMux I__4171 (
            .O(N__18797),
            .I(N__18794));
    LocalMux I__4170 (
            .O(N__18794),
            .I(N__18790));
    InMux I__4169 (
            .O(N__18793),
            .I(N__18787));
    Span4Mux_v I__4168 (
            .O(N__18790),
            .I(N__18782));
    LocalMux I__4167 (
            .O(N__18787),
            .I(N__18782));
    Span4Mux_h I__4166 (
            .O(N__18782),
            .I(N__18779));
    Odrv4 I__4165 (
            .O(N__18779),
            .I(data_out_6_3));
    InMux I__4164 (
            .O(N__18776),
            .I(N__18772));
    InMux I__4163 (
            .O(N__18775),
            .I(N__18769));
    LocalMux I__4162 (
            .O(N__18772),
            .I(\c0.delay_counter_6 ));
    LocalMux I__4161 (
            .O(N__18769),
            .I(\c0.delay_counter_6 ));
    CascadeMux I__4160 (
            .O(N__18764),
            .I(N__18761));
    InMux I__4159 (
            .O(N__18761),
            .I(N__18757));
    InMux I__4158 (
            .O(N__18760),
            .I(N__18754));
    LocalMux I__4157 (
            .O(N__18757),
            .I(\c0.delay_counter_0 ));
    LocalMux I__4156 (
            .O(N__18754),
            .I(\c0.delay_counter_0 ));
    CascadeMux I__4155 (
            .O(N__18749),
            .I(N__18745));
    InMux I__4154 (
            .O(N__18748),
            .I(N__18742));
    InMux I__4153 (
            .O(N__18745),
            .I(N__18739));
    LocalMux I__4152 (
            .O(N__18742),
            .I(\c0.delay_counter_2 ));
    LocalMux I__4151 (
            .O(N__18739),
            .I(\c0.delay_counter_2 ));
    InMux I__4150 (
            .O(N__18734),
            .I(N__18730));
    InMux I__4149 (
            .O(N__18733),
            .I(N__18727));
    LocalMux I__4148 (
            .O(N__18730),
            .I(\c0.delay_counter_4 ));
    LocalMux I__4147 (
            .O(N__18727),
            .I(\c0.delay_counter_4 ));
    InMux I__4146 (
            .O(N__18722),
            .I(N__18718));
    InMux I__4145 (
            .O(N__18721),
            .I(N__18715));
    LocalMux I__4144 (
            .O(N__18718),
            .I(\c0.delay_counter_5 ));
    LocalMux I__4143 (
            .O(N__18715),
            .I(\c0.delay_counter_5 ));
    InMux I__4142 (
            .O(N__18710),
            .I(N__18706));
    InMux I__4141 (
            .O(N__18709),
            .I(N__18703));
    LocalMux I__4140 (
            .O(N__18706),
            .I(\c0.delay_counter_1 ));
    LocalMux I__4139 (
            .O(N__18703),
            .I(\c0.delay_counter_1 ));
    CascadeMux I__4138 (
            .O(N__18698),
            .I(N__18694));
    InMux I__4137 (
            .O(N__18697),
            .I(N__18691));
    InMux I__4136 (
            .O(N__18694),
            .I(N__18688));
    LocalMux I__4135 (
            .O(N__18691),
            .I(\c0.delay_counter_7 ));
    LocalMux I__4134 (
            .O(N__18688),
            .I(\c0.delay_counter_7 ));
    InMux I__4133 (
            .O(N__18683),
            .I(N__18679));
    InMux I__4132 (
            .O(N__18682),
            .I(N__18676));
    LocalMux I__4131 (
            .O(N__18679),
            .I(\c0.delay_counter_3 ));
    LocalMux I__4130 (
            .O(N__18676),
            .I(\c0.delay_counter_3 ));
    InMux I__4129 (
            .O(N__18671),
            .I(N__18668));
    LocalMux I__4128 (
            .O(N__18668),
            .I(\c0.n13 ));
    CascadeMux I__4127 (
            .O(N__18665),
            .I(\c0.n14_adj_902_cascade_ ));
    InMux I__4126 (
            .O(N__18662),
            .I(N__18659));
    LocalMux I__4125 (
            .O(N__18659),
            .I(N__18655));
    InMux I__4124 (
            .O(N__18658),
            .I(N__18652));
    Odrv12 I__4123 (
            .O(N__18655),
            .I(\c0.data_4 ));
    LocalMux I__4122 (
            .O(N__18652),
            .I(\c0.data_4 ));
    CascadeMux I__4121 (
            .O(N__18647),
            .I(n3580_cascade_));
    CascadeMux I__4120 (
            .O(N__18644),
            .I(N__18641));
    InMux I__4119 (
            .O(N__18641),
            .I(N__18638));
    LocalMux I__4118 (
            .O(N__18638),
            .I(N__18635));
    Span4Mux_h I__4117 (
            .O(N__18635),
            .I(N__18631));
    InMux I__4116 (
            .O(N__18634),
            .I(N__18628));
    Odrv4 I__4115 (
            .O(N__18631),
            .I(\c0.data_11 ));
    LocalMux I__4114 (
            .O(N__18628),
            .I(\c0.data_11 ));
    CascadeMux I__4113 (
            .O(N__18623),
            .I(N__18620));
    InMux I__4112 (
            .O(N__18620),
            .I(N__18617));
    LocalMux I__4111 (
            .O(N__18617),
            .I(N__18614));
    Span4Mux_h I__4110 (
            .O(N__18614),
            .I(N__18610));
    InMux I__4109 (
            .O(N__18613),
            .I(N__18607));
    Odrv4 I__4108 (
            .O(N__18610),
            .I(\c0.data_3 ));
    LocalMux I__4107 (
            .O(N__18607),
            .I(\c0.data_3 ));
    InMux I__4106 (
            .O(N__18602),
            .I(N__18599));
    LocalMux I__4105 (
            .O(N__18599),
            .I(n7_adj_933));
    InMux I__4104 (
            .O(N__18596),
            .I(N__18593));
    LocalMux I__4103 (
            .O(N__18593),
            .I(N__18589));
    InMux I__4102 (
            .O(N__18592),
            .I(N__18586));
    Span4Mux_s3_v I__4101 (
            .O(N__18589),
            .I(N__18579));
    LocalMux I__4100 (
            .O(N__18586),
            .I(N__18579));
    InMux I__4099 (
            .O(N__18585),
            .I(N__18576));
    InMux I__4098 (
            .O(N__18584),
            .I(N__18573));
    Span4Mux_h I__4097 (
            .O(N__18579),
            .I(N__18570));
    LocalMux I__4096 (
            .O(N__18576),
            .I(\c0.data_out_field_47_N_682_41 ));
    LocalMux I__4095 (
            .O(N__18573),
            .I(\c0.data_out_field_47_N_682_41 ));
    Odrv4 I__4094 (
            .O(N__18570),
            .I(\c0.data_out_field_47_N_682_41 ));
    InMux I__4093 (
            .O(N__18563),
            .I(N__18559));
    InMux I__4092 (
            .O(N__18562),
            .I(N__18553));
    LocalMux I__4091 (
            .O(N__18559),
            .I(N__18550));
    InMux I__4090 (
            .O(N__18558),
            .I(N__18547));
    CascadeMux I__4089 (
            .O(N__18557),
            .I(N__18544));
    InMux I__4088 (
            .O(N__18556),
            .I(N__18541));
    LocalMux I__4087 (
            .O(N__18553),
            .I(N__18538));
    Span4Mux_v I__4086 (
            .O(N__18550),
            .I(N__18533));
    LocalMux I__4085 (
            .O(N__18547),
            .I(N__18533));
    InMux I__4084 (
            .O(N__18544),
            .I(N__18530));
    LocalMux I__4083 (
            .O(N__18541),
            .I(N__18523));
    Span4Mux_h I__4082 (
            .O(N__18538),
            .I(N__18523));
    Span4Mux_h I__4081 (
            .O(N__18533),
            .I(N__18523));
    LocalMux I__4080 (
            .O(N__18530),
            .I(\c0.data_out_field_47_N_682_34 ));
    Odrv4 I__4079 (
            .O(N__18523),
            .I(\c0.data_out_field_47_N_682_34 ));
    CascadeMux I__4078 (
            .O(N__18518),
            .I(\c0.n1384_cascade_ ));
    InMux I__4077 (
            .O(N__18515),
            .I(N__18512));
    LocalMux I__4076 (
            .O(N__18512),
            .I(N__18505));
    InMux I__4075 (
            .O(N__18511),
            .I(N__18502));
    InMux I__4074 (
            .O(N__18510),
            .I(N__18497));
    InMux I__4073 (
            .O(N__18509),
            .I(N__18497));
    InMux I__4072 (
            .O(N__18508),
            .I(N__18494));
    Span4Mux_v I__4071 (
            .O(N__18505),
            .I(N__18491));
    LocalMux I__4070 (
            .O(N__18502),
            .I(N__18486));
    LocalMux I__4069 (
            .O(N__18497),
            .I(N__18486));
    LocalMux I__4068 (
            .O(N__18494),
            .I(\c0.data_out_field_47_N_682_32 ));
    Odrv4 I__4067 (
            .O(N__18491),
            .I(\c0.data_out_field_47_N_682_32 ));
    Odrv4 I__4066 (
            .O(N__18486),
            .I(\c0.data_out_field_47_N_682_32 ));
    InMux I__4065 (
            .O(N__18479),
            .I(N__18476));
    LocalMux I__4064 (
            .O(N__18476),
            .I(N__18472));
    InMux I__4063 (
            .O(N__18475),
            .I(N__18467));
    Span4Mux_h I__4062 (
            .O(N__18472),
            .I(N__18464));
    InMux I__4061 (
            .O(N__18471),
            .I(N__18459));
    InMux I__4060 (
            .O(N__18470),
            .I(N__18459));
    LocalMux I__4059 (
            .O(N__18467),
            .I(data_out_field_3));
    Odrv4 I__4058 (
            .O(N__18464),
            .I(data_out_field_3));
    LocalMux I__4057 (
            .O(N__18459),
            .I(data_out_field_3));
    InMux I__4056 (
            .O(N__18452),
            .I(N__18447));
    CascadeMux I__4055 (
            .O(N__18451),
            .I(N__18443));
    InMux I__4054 (
            .O(N__18450),
            .I(N__18440));
    LocalMux I__4053 (
            .O(N__18447),
            .I(N__18437));
    InMux I__4052 (
            .O(N__18446),
            .I(N__18432));
    InMux I__4051 (
            .O(N__18443),
            .I(N__18432));
    LocalMux I__4050 (
            .O(N__18440),
            .I(N__18427));
    Span4Mux_v I__4049 (
            .O(N__18437),
            .I(N__18427));
    LocalMux I__4048 (
            .O(N__18432),
            .I(N__18424));
    Odrv4 I__4047 (
            .O(N__18427),
            .I(data_out_field_4));
    Odrv4 I__4046 (
            .O(N__18424),
            .I(data_out_field_4));
    InMux I__4045 (
            .O(N__18419),
            .I(N__18416));
    LocalMux I__4044 (
            .O(N__18416),
            .I(N__18413));
    Span4Mux_h I__4043 (
            .O(N__18413),
            .I(N__18410));
    Odrv4 I__4042 (
            .O(N__18410),
            .I(\c0.n4529 ));
    InMux I__4041 (
            .O(N__18407),
            .I(N__18404));
    LocalMux I__4040 (
            .O(N__18404),
            .I(N__18401));
    Span4Mux_v I__4039 (
            .O(N__18401),
            .I(N__18398));
    Odrv4 I__4038 (
            .O(N__18398),
            .I(n7_adj_937));
    InMux I__4037 (
            .O(N__18395),
            .I(N__18392));
    LocalMux I__4036 (
            .O(N__18392),
            .I(N__18389));
    Odrv4 I__4035 (
            .O(N__18389),
            .I(\c0.n4565 ));
    CascadeMux I__4034 (
            .O(N__18386),
            .I(n11_adj_967_cascade_));
    InMux I__4033 (
            .O(N__18383),
            .I(N__18380));
    LocalMux I__4032 (
            .O(N__18380),
            .I(N__18376));
    InMux I__4031 (
            .O(N__18379),
            .I(N__18373));
    Span4Mux_v I__4030 (
            .O(N__18376),
            .I(N__18370));
    LocalMux I__4029 (
            .O(N__18373),
            .I(data_out_7_4));
    Odrv4 I__4028 (
            .O(N__18370),
            .I(data_out_7_4));
    InMux I__4027 (
            .O(N__18365),
            .I(N__18361));
    InMux I__4026 (
            .O(N__18364),
            .I(N__18358));
    LocalMux I__4025 (
            .O(N__18361),
            .I(N__18353));
    LocalMux I__4024 (
            .O(N__18358),
            .I(N__18350));
    InMux I__4023 (
            .O(N__18357),
            .I(N__18347));
    InMux I__4022 (
            .O(N__18356),
            .I(N__18344));
    Span4Mux_h I__4021 (
            .O(N__18353),
            .I(N__18337));
    Span4Mux_h I__4020 (
            .O(N__18350),
            .I(N__18337));
    LocalMux I__4019 (
            .O(N__18347),
            .I(N__18337));
    LocalMux I__4018 (
            .O(N__18344),
            .I(data_out_field_11));
    Odrv4 I__4017 (
            .O(N__18337),
            .I(data_out_field_11));
    CascadeMux I__4016 (
            .O(N__18332),
            .I(\c0.n6_cascade_ ));
    InMux I__4015 (
            .O(N__18329),
            .I(N__18324));
    InMux I__4014 (
            .O(N__18328),
            .I(N__18321));
    InMux I__4013 (
            .O(N__18327),
            .I(N__18318));
    LocalMux I__4012 (
            .O(N__18324),
            .I(N__18315));
    LocalMux I__4011 (
            .O(N__18321),
            .I(N__18309));
    LocalMux I__4010 (
            .O(N__18318),
            .I(N__18309));
    Span4Mux_h I__4009 (
            .O(N__18315),
            .I(N__18306));
    InMux I__4008 (
            .O(N__18314),
            .I(N__18303));
    Span4Mux_v I__4007 (
            .O(N__18309),
            .I(N__18300));
    Span4Mux_v I__4006 (
            .O(N__18306),
            .I(N__18297));
    LocalMux I__4005 (
            .O(N__18303),
            .I(data_out_field_24));
    Odrv4 I__4004 (
            .O(N__18300),
            .I(data_out_field_24));
    Odrv4 I__4003 (
            .O(N__18297),
            .I(data_out_field_24));
    CascadeMux I__4002 (
            .O(N__18290),
            .I(\c0.n4456_cascade_ ));
    CascadeMux I__4001 (
            .O(N__18287),
            .I(N__18284));
    InMux I__4000 (
            .O(N__18284),
            .I(N__18281));
    LocalMux I__3999 (
            .O(N__18281),
            .I(N__18278));
    Span4Mux_v I__3998 (
            .O(N__18278),
            .I(N__18274));
    InMux I__3997 (
            .O(N__18277),
            .I(N__18271));
    Odrv4 I__3996 (
            .O(N__18274),
            .I(\c0.data_0 ));
    LocalMux I__3995 (
            .O(N__18271),
            .I(\c0.data_0 ));
    InMux I__3994 (
            .O(N__18266),
            .I(N__18262));
    InMux I__3993 (
            .O(N__18265),
            .I(N__18258));
    LocalMux I__3992 (
            .O(N__18262),
            .I(N__18255));
    InMux I__3991 (
            .O(N__18261),
            .I(N__18252));
    LocalMux I__3990 (
            .O(N__18258),
            .I(data_out_field_17));
    Odrv4 I__3989 (
            .O(N__18255),
            .I(data_out_field_17));
    LocalMux I__3988 (
            .O(N__18252),
            .I(data_out_field_17));
    InMux I__3987 (
            .O(N__18245),
            .I(N__18242));
    LocalMux I__3986 (
            .O(N__18242),
            .I(N__18239));
    Span4Mux_h I__3985 (
            .O(N__18239),
            .I(N__18236));
    Odrv4 I__3984 (
            .O(N__18236),
            .I(\c0.n4562 ));
    InMux I__3983 (
            .O(N__18233),
            .I(N__18230));
    LocalMux I__3982 (
            .O(N__18230),
            .I(N__18226));
    InMux I__3981 (
            .O(N__18229),
            .I(N__18223));
    Span4Mux_v I__3980 (
            .O(N__18226),
            .I(N__18220));
    LocalMux I__3979 (
            .O(N__18223),
            .I(data_out_7_2));
    Odrv4 I__3978 (
            .O(N__18220),
            .I(data_out_7_2));
    InMux I__3977 (
            .O(N__18215),
            .I(N__18211));
    InMux I__3976 (
            .O(N__18214),
            .I(N__18208));
    LocalMux I__3975 (
            .O(N__18211),
            .I(N__18203));
    LocalMux I__3974 (
            .O(N__18208),
            .I(N__18203));
    Odrv12 I__3973 (
            .O(N__18203),
            .I(data_out_7_1));
    InMux I__3972 (
            .O(N__18200),
            .I(N__18197));
    LocalMux I__3971 (
            .O(N__18197),
            .I(N__18194));
    Odrv12 I__3970 (
            .O(N__18194),
            .I(\c0.n4574 ));
    InMux I__3969 (
            .O(N__18191),
            .I(N__18188));
    LocalMux I__3968 (
            .O(N__18188),
            .I(N__18185));
    Span12Mux_h I__3967 (
            .O(N__18185),
            .I(N__18181));
    InMux I__3966 (
            .O(N__18184),
            .I(N__18178));
    Odrv12 I__3965 (
            .O(N__18181),
            .I(\c0.data_10 ));
    LocalMux I__3964 (
            .O(N__18178),
            .I(\c0.data_10 ));
    InMux I__3963 (
            .O(N__18173),
            .I(N__18169));
    InMux I__3962 (
            .O(N__18172),
            .I(N__18166));
    LocalMux I__3961 (
            .O(N__18169),
            .I(N__18162));
    LocalMux I__3960 (
            .O(N__18166),
            .I(N__18159));
    InMux I__3959 (
            .O(N__18165),
            .I(N__18156));
    Span4Mux_v I__3958 (
            .O(N__18162),
            .I(N__18153));
    Span4Mux_h I__3957 (
            .O(N__18159),
            .I(N__18150));
    LocalMux I__3956 (
            .O(N__18156),
            .I(data_out_field_19));
    Odrv4 I__3955 (
            .O(N__18153),
            .I(data_out_field_19));
    Odrv4 I__3954 (
            .O(N__18150),
            .I(data_out_field_19));
    InMux I__3953 (
            .O(N__18143),
            .I(N__18140));
    LocalMux I__3952 (
            .O(N__18140),
            .I(n8_adj_936));
    InMux I__3951 (
            .O(N__18137),
            .I(N__18133));
    InMux I__3950 (
            .O(N__18136),
            .I(N__18130));
    LocalMux I__3949 (
            .O(N__18133),
            .I(N__18127));
    LocalMux I__3948 (
            .O(N__18130),
            .I(data_out_6_2));
    Odrv4 I__3947 (
            .O(N__18127),
            .I(data_out_6_2));
    InMux I__3946 (
            .O(N__18122),
            .I(N__18119));
    LocalMux I__3945 (
            .O(N__18119),
            .I(\c0.n2429 ));
    CascadeMux I__3944 (
            .O(N__18116),
            .I(N__18113));
    InMux I__3943 (
            .O(N__18113),
            .I(N__18110));
    LocalMux I__3942 (
            .O(N__18110),
            .I(N__18107));
    Span4Mux_h I__3941 (
            .O(N__18107),
            .I(N__18103));
    InMux I__3940 (
            .O(N__18106),
            .I(N__18100));
    Odrv4 I__3939 (
            .O(N__18103),
            .I(\c0.data_6 ));
    LocalMux I__3938 (
            .O(N__18100),
            .I(\c0.data_6 ));
    InMux I__3937 (
            .O(N__18095),
            .I(N__18092));
    LocalMux I__3936 (
            .O(N__18092),
            .I(N__18089));
    Span4Mux_h I__3935 (
            .O(N__18089),
            .I(N__18085));
    InMux I__3934 (
            .O(N__18088),
            .I(N__18082));
    Odrv4 I__3933 (
            .O(N__18085),
            .I(\c0.data_7 ));
    LocalMux I__3932 (
            .O(N__18082),
            .I(\c0.data_7 ));
    CascadeMux I__3931 (
            .O(N__18077),
            .I(N__18074));
    InMux I__3930 (
            .O(N__18074),
            .I(N__18071));
    LocalMux I__3929 (
            .O(N__18071),
            .I(N__18068));
    Span4Mux_h I__3928 (
            .O(N__18068),
            .I(N__18064));
    InMux I__3927 (
            .O(N__18067),
            .I(N__18061));
    Odrv4 I__3926 (
            .O(N__18064),
            .I(\c0.data_14 ));
    LocalMux I__3925 (
            .O(N__18061),
            .I(\c0.data_14 ));
    InMux I__3924 (
            .O(N__18056),
            .I(N__18052));
    InMux I__3923 (
            .O(N__18055),
            .I(N__18049));
    LocalMux I__3922 (
            .O(N__18052),
            .I(N__18046));
    LocalMux I__3921 (
            .O(N__18049),
            .I(N__18041));
    Span4Mux_v I__3920 (
            .O(N__18046),
            .I(N__18041));
    Odrv4 I__3919 (
            .O(N__18041),
            .I(data_out_7_3));
    CascadeMux I__3918 (
            .O(N__18038),
            .I(N__18035));
    InMux I__3917 (
            .O(N__18035),
            .I(N__18032));
    LocalMux I__3916 (
            .O(N__18032),
            .I(N__18029));
    Span4Mux_h I__3915 (
            .O(N__18029),
            .I(N__18025));
    InMux I__3914 (
            .O(N__18028),
            .I(N__18022));
    Odrv4 I__3913 (
            .O(N__18025),
            .I(\c0.data_8 ));
    LocalMux I__3912 (
            .O(N__18022),
            .I(\c0.data_8 ));
    CascadeMux I__3911 (
            .O(N__18017),
            .I(n8_adj_932_cascade_));
    InMux I__3910 (
            .O(N__18014),
            .I(\c0.n3901 ));
    InMux I__3909 (
            .O(N__18011),
            .I(\c0.n3902 ));
    InMux I__3908 (
            .O(N__18008),
            .I(\c0.n3903 ));
    InMux I__3907 (
            .O(N__18005),
            .I(\c0.n3904 ));
    InMux I__3906 (
            .O(N__18002),
            .I(\c0.n3905 ));
    InMux I__3905 (
            .O(N__17999),
            .I(N__17996));
    LocalMux I__3904 (
            .O(N__17996),
            .I(N__17992));
    InMux I__3903 (
            .O(N__17995),
            .I(N__17989));
    Span4Mux_h I__3902 (
            .O(N__17992),
            .I(N__17986));
    LocalMux I__3901 (
            .O(N__17989),
            .I(data_out_6_1));
    Odrv4 I__3900 (
            .O(N__17986),
            .I(data_out_6_1));
    InMux I__3899 (
            .O(N__17981),
            .I(N__17978));
    LocalMux I__3898 (
            .O(N__17978),
            .I(N__17974));
    InMux I__3897 (
            .O(N__17977),
            .I(N__17971));
    Span4Mux_h I__3896 (
            .O(N__17974),
            .I(N__17968));
    LocalMux I__3895 (
            .O(N__17971),
            .I(\c0.data_15 ));
    Odrv4 I__3894 (
            .O(N__17968),
            .I(\c0.data_15 ));
    InMux I__3893 (
            .O(N__17963),
            .I(N__17960));
    LocalMux I__3892 (
            .O(N__17960),
            .I(N__17957));
    Odrv12 I__3891 (
            .O(N__17957),
            .I(\c0.n4888 ));
    InMux I__3890 (
            .O(N__17954),
            .I(N__17951));
    LocalMux I__3889 (
            .O(N__17951),
            .I(\c0.rx.n4093 ));
    InMux I__3888 (
            .O(N__17948),
            .I(N__17945));
    LocalMux I__3887 (
            .O(N__17945),
            .I(\c0.rx.n4378 ));
    CascadeMux I__3886 (
            .O(N__17942),
            .I(\c0.rx.n13_cascade_ ));
    InMux I__3885 (
            .O(N__17939),
            .I(N__17936));
    LocalMux I__3884 (
            .O(N__17936),
            .I(\c0.rx.n6 ));
    CascadeMux I__3883 (
            .O(N__17933),
            .I(N__17926));
    InMux I__3882 (
            .O(N__17932),
            .I(N__17921));
    InMux I__3881 (
            .O(N__17931),
            .I(N__17914));
    InMux I__3880 (
            .O(N__17930),
            .I(N__17914));
    InMux I__3879 (
            .O(N__17929),
            .I(N__17914));
    InMux I__3878 (
            .O(N__17926),
            .I(N__17907));
    InMux I__3877 (
            .O(N__17925),
            .I(N__17907));
    InMux I__3876 (
            .O(N__17924),
            .I(N__17907));
    LocalMux I__3875 (
            .O(N__17921),
            .I(n1554));
    LocalMux I__3874 (
            .O(N__17914),
            .I(n1554));
    LocalMux I__3873 (
            .O(N__17907),
            .I(n1554));
    InMux I__3872 (
            .O(N__17900),
            .I(N__17897));
    LocalMux I__3871 (
            .O(N__17897),
            .I(N__17894));
    Odrv4 I__3870 (
            .O(N__17894),
            .I(n220));
    InMux I__3869 (
            .O(N__17891),
            .I(N__17883));
    InMux I__3868 (
            .O(N__17890),
            .I(N__17880));
    InMux I__3867 (
            .O(N__17889),
            .I(N__17875));
    InMux I__3866 (
            .O(N__17888),
            .I(N__17875));
    InMux I__3865 (
            .O(N__17887),
            .I(N__17870));
    InMux I__3864 (
            .O(N__17886),
            .I(N__17870));
    LocalMux I__3863 (
            .O(N__17883),
            .I(n573));
    LocalMux I__3862 (
            .O(N__17880),
            .I(n573));
    LocalMux I__3861 (
            .O(N__17875),
            .I(n573));
    LocalMux I__3860 (
            .O(N__17870),
            .I(n573));
    CascadeMux I__3859 (
            .O(N__17861),
            .I(n1554_cascade_));
    InMux I__3858 (
            .O(N__17858),
            .I(N__17852));
    InMux I__3857 (
            .O(N__17857),
            .I(N__17847));
    InMux I__3856 (
            .O(N__17856),
            .I(N__17847));
    InMux I__3855 (
            .O(N__17855),
            .I(N__17843));
    LocalMux I__3854 (
            .O(N__17852),
            .I(N__17838));
    LocalMux I__3853 (
            .O(N__17847),
            .I(N__17838));
    InMux I__3852 (
            .O(N__17846),
            .I(N__17834));
    LocalMux I__3851 (
            .O(N__17843),
            .I(N__17831));
    Span4Mux_v I__3850 (
            .O(N__17838),
            .I(N__17828));
    InMux I__3849 (
            .O(N__17837),
            .I(N__17825));
    LocalMux I__3848 (
            .O(N__17834),
            .I(r_Clock_Count_6));
    Odrv4 I__3847 (
            .O(N__17831),
            .I(r_Clock_Count_6));
    Odrv4 I__3846 (
            .O(N__17828),
            .I(r_Clock_Count_6));
    LocalMux I__3845 (
            .O(N__17825),
            .I(r_Clock_Count_6));
    InMux I__3844 (
            .O(N__17816),
            .I(N__17813));
    LocalMux I__3843 (
            .O(N__17813),
            .I(N__17810));
    Span4Mux_s1_v I__3842 (
            .O(N__17810),
            .I(N__17804));
    InMux I__3841 (
            .O(N__17809),
            .I(N__17801));
    InMux I__3840 (
            .O(N__17808),
            .I(N__17796));
    InMux I__3839 (
            .O(N__17807),
            .I(N__17796));
    Odrv4 I__3838 (
            .O(N__17804),
            .I(\c0.rx.n2179 ));
    LocalMux I__3837 (
            .O(N__17801),
            .I(\c0.rx.n2179 ));
    LocalMux I__3836 (
            .O(N__17796),
            .I(\c0.rx.n2179 ));
    CascadeMux I__3835 (
            .O(N__17789),
            .I(N__17785));
    CascadeMux I__3834 (
            .O(N__17788),
            .I(N__17782));
    InMux I__3833 (
            .O(N__17785),
            .I(N__17773));
    InMux I__3832 (
            .O(N__17782),
            .I(N__17773));
    InMux I__3831 (
            .O(N__17781),
            .I(N__17768));
    InMux I__3830 (
            .O(N__17780),
            .I(N__17768));
    CascadeMux I__3829 (
            .O(N__17779),
            .I(N__17763));
    CascadeMux I__3828 (
            .O(N__17778),
            .I(N__17757));
    LocalMux I__3827 (
            .O(N__17773),
            .I(N__17753));
    LocalMux I__3826 (
            .O(N__17768),
            .I(N__17750));
    InMux I__3825 (
            .O(N__17767),
            .I(N__17745));
    InMux I__3824 (
            .O(N__17766),
            .I(N__17745));
    InMux I__3823 (
            .O(N__17763),
            .I(N__17736));
    InMux I__3822 (
            .O(N__17762),
            .I(N__17736));
    InMux I__3821 (
            .O(N__17761),
            .I(N__17736));
    InMux I__3820 (
            .O(N__17760),
            .I(N__17736));
    InMux I__3819 (
            .O(N__17757),
            .I(N__17733));
    InMux I__3818 (
            .O(N__17756),
            .I(N__17730));
    Span4Mux_h I__3817 (
            .O(N__17753),
            .I(N__17727));
    Span4Mux_v I__3816 (
            .O(N__17750),
            .I(N__17720));
    LocalMux I__3815 (
            .O(N__17745),
            .I(N__17720));
    LocalMux I__3814 (
            .O(N__17736),
            .I(N__17720));
    LocalMux I__3813 (
            .O(N__17733),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__3812 (
            .O(N__17730),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv4 I__3811 (
            .O(N__17727),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv4 I__3810 (
            .O(N__17720),
            .I(\c0.rx.r_SM_Main_0 ));
    InMux I__3809 (
            .O(N__17711),
            .I(N__17702));
    InMux I__3808 (
            .O(N__17710),
            .I(N__17697));
    InMux I__3807 (
            .O(N__17709),
            .I(N__17697));
    InMux I__3806 (
            .O(N__17708),
            .I(N__17688));
    InMux I__3805 (
            .O(N__17707),
            .I(N__17688));
    InMux I__3804 (
            .O(N__17706),
            .I(N__17688));
    InMux I__3803 (
            .O(N__17705),
            .I(N__17688));
    LocalMux I__3802 (
            .O(N__17702),
            .I(N__17680));
    LocalMux I__3801 (
            .O(N__17697),
            .I(N__17675));
    LocalMux I__3800 (
            .O(N__17688),
            .I(N__17675));
    InMux I__3799 (
            .O(N__17687),
            .I(N__17672));
    InMux I__3798 (
            .O(N__17686),
            .I(N__17669));
    InMux I__3797 (
            .O(N__17685),
            .I(N__17666));
    InMux I__3796 (
            .O(N__17684),
            .I(N__17663));
    InMux I__3795 (
            .O(N__17683),
            .I(N__17660));
    Span4Mux_h I__3794 (
            .O(N__17680),
            .I(N__17655));
    Span4Mux_h I__3793 (
            .O(N__17675),
            .I(N__17655));
    LocalMux I__3792 (
            .O(N__17672),
            .I(N__17646));
    LocalMux I__3791 (
            .O(N__17669),
            .I(N__17646));
    LocalMux I__3790 (
            .O(N__17666),
            .I(N__17646));
    LocalMux I__3789 (
            .O(N__17663),
            .I(N__17646));
    LocalMux I__3788 (
            .O(N__17660),
            .I(r_Rx_Data));
    Odrv4 I__3787 (
            .O(N__17655),
            .I(r_Rx_Data));
    Odrv12 I__3786 (
            .O(N__17646),
            .I(r_Rx_Data));
    InMux I__3785 (
            .O(N__17639),
            .I(N__17634));
    InMux I__3784 (
            .O(N__17638),
            .I(N__17622));
    InMux I__3783 (
            .O(N__17637),
            .I(N__17622));
    LocalMux I__3782 (
            .O(N__17634),
            .I(N__17615));
    InMux I__3781 (
            .O(N__17633),
            .I(N__17612));
    InMux I__3780 (
            .O(N__17632),
            .I(N__17607));
    InMux I__3779 (
            .O(N__17631),
            .I(N__17607));
    InMux I__3778 (
            .O(N__17630),
            .I(N__17598));
    InMux I__3777 (
            .O(N__17629),
            .I(N__17598));
    InMux I__3776 (
            .O(N__17628),
            .I(N__17598));
    InMux I__3775 (
            .O(N__17627),
            .I(N__17598));
    LocalMux I__3774 (
            .O(N__17622),
            .I(N__17595));
    InMux I__3773 (
            .O(N__17621),
            .I(N__17588));
    InMux I__3772 (
            .O(N__17620),
            .I(N__17588));
    InMux I__3771 (
            .O(N__17619),
            .I(N__17588));
    InMux I__3770 (
            .O(N__17618),
            .I(N__17585));
    Span4Mux_h I__3769 (
            .O(N__17615),
            .I(N__17576));
    LocalMux I__3768 (
            .O(N__17612),
            .I(N__17576));
    LocalMux I__3767 (
            .O(N__17607),
            .I(N__17576));
    LocalMux I__3766 (
            .O(N__17598),
            .I(N__17576));
    Odrv4 I__3765 (
            .O(N__17595),
            .I(\c0.rx.r_SM_Main_2 ));
    LocalMux I__3764 (
            .O(N__17588),
            .I(\c0.rx.r_SM_Main_2 ));
    LocalMux I__3763 (
            .O(N__17585),
            .I(\c0.rx.r_SM_Main_2 ));
    Odrv4 I__3762 (
            .O(N__17576),
            .I(\c0.rx.r_SM_Main_2 ));
    CascadeMux I__3761 (
            .O(N__17567),
            .I(\c0.rx.n4666_cascade_ ));
    InMux I__3760 (
            .O(N__17564),
            .I(N__17561));
    LocalMux I__3759 (
            .O(N__17561),
            .I(\c0.rx.n4667 ));
    InMux I__3758 (
            .O(N__17558),
            .I(N__17545));
    InMux I__3757 (
            .O(N__17557),
            .I(N__17545));
    InMux I__3756 (
            .O(N__17556),
            .I(N__17537));
    InMux I__3755 (
            .O(N__17555),
            .I(N__17537));
    InMux I__3754 (
            .O(N__17554),
            .I(N__17528));
    InMux I__3753 (
            .O(N__17553),
            .I(N__17528));
    InMux I__3752 (
            .O(N__17552),
            .I(N__17528));
    InMux I__3751 (
            .O(N__17551),
            .I(N__17528));
    CascadeMux I__3750 (
            .O(N__17550),
            .I(N__17525));
    LocalMux I__3749 (
            .O(N__17545),
            .I(N__17521));
    CascadeMux I__3748 (
            .O(N__17544),
            .I(N__17518));
    InMux I__3747 (
            .O(N__17543),
            .I(N__17513));
    InMux I__3746 (
            .O(N__17542),
            .I(N__17510));
    LocalMux I__3745 (
            .O(N__17537),
            .I(N__17507));
    LocalMux I__3744 (
            .O(N__17528),
            .I(N__17504));
    InMux I__3743 (
            .O(N__17525),
            .I(N__17499));
    InMux I__3742 (
            .O(N__17524),
            .I(N__17499));
    Span4Mux_h I__3741 (
            .O(N__17521),
            .I(N__17496));
    InMux I__3740 (
            .O(N__17518),
            .I(N__17489));
    InMux I__3739 (
            .O(N__17517),
            .I(N__17489));
    InMux I__3738 (
            .O(N__17516),
            .I(N__17489));
    LocalMux I__3737 (
            .O(N__17513),
            .I(\c0.rx.r_SM_Main_1 ));
    LocalMux I__3736 (
            .O(N__17510),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv12 I__3735 (
            .O(N__17507),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv4 I__3734 (
            .O(N__17504),
            .I(\c0.rx.r_SM_Main_1 ));
    LocalMux I__3733 (
            .O(N__17499),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv4 I__3732 (
            .O(N__17496),
            .I(\c0.rx.r_SM_Main_1 ));
    LocalMux I__3731 (
            .O(N__17489),
            .I(\c0.rx.r_SM_Main_1 ));
    InMux I__3730 (
            .O(N__17474),
            .I(\c0.n3899 ));
    InMux I__3729 (
            .O(N__17471),
            .I(\c0.n3900 ));
    CascadeMux I__3728 (
            .O(N__17468),
            .I(N__17465));
    InMux I__3727 (
            .O(N__17465),
            .I(N__17462));
    LocalMux I__3726 (
            .O(N__17462),
            .I(N__17459));
    Span4Mux_v I__3725 (
            .O(N__17459),
            .I(N__17455));
    InMux I__3724 (
            .O(N__17458),
            .I(N__17452));
    Sp12to4 I__3723 (
            .O(N__17455),
            .I(N__17446));
    LocalMux I__3722 (
            .O(N__17452),
            .I(N__17446));
    InMux I__3721 (
            .O(N__17451),
            .I(N__17443));
    Odrv12 I__3720 (
            .O(N__17446),
            .I(data_in_5_1));
    LocalMux I__3719 (
            .O(N__17443),
            .I(data_in_5_1));
    CascadeMux I__3718 (
            .O(N__17438),
            .I(N__17435));
    InMux I__3717 (
            .O(N__17435),
            .I(N__17432));
    LocalMux I__3716 (
            .O(N__17432),
            .I(N__17429));
    Span4Mux_h I__3715 (
            .O(N__17429),
            .I(N__17426));
    Odrv4 I__3714 (
            .O(N__17426),
            .I(n224));
    InMux I__3713 (
            .O(N__17423),
            .I(N__17420));
    LocalMux I__3712 (
            .O(N__17420),
            .I(N__17413));
    InMux I__3711 (
            .O(N__17419),
            .I(N__17410));
    InMux I__3710 (
            .O(N__17418),
            .I(N__17407));
    InMux I__3709 (
            .O(N__17417),
            .I(N__17404));
    InMux I__3708 (
            .O(N__17416),
            .I(N__17401));
    Span4Mux_h I__3707 (
            .O(N__17413),
            .I(N__17396));
    LocalMux I__3706 (
            .O(N__17410),
            .I(N__17396));
    LocalMux I__3705 (
            .O(N__17407),
            .I(r_Clock_Count_2));
    LocalMux I__3704 (
            .O(N__17404),
            .I(r_Clock_Count_2));
    LocalMux I__3703 (
            .O(N__17401),
            .I(r_Clock_Count_2));
    Odrv4 I__3702 (
            .O(N__17396),
            .I(r_Clock_Count_2));
    InMux I__3701 (
            .O(N__17387),
            .I(N__17384));
    LocalMux I__3700 (
            .O(N__17384),
            .I(N__17381));
    Odrv12 I__3699 (
            .O(N__17381),
            .I(\c0.n4528 ));
    InMux I__3698 (
            .O(N__17378),
            .I(N__17375));
    LocalMux I__3697 (
            .O(N__17375),
            .I(N__17369));
    InMux I__3696 (
            .O(N__17374),
            .I(N__17364));
    InMux I__3695 (
            .O(N__17373),
            .I(N__17360));
    InMux I__3694 (
            .O(N__17372),
            .I(N__17357));
    Span4Mux_s2_v I__3693 (
            .O(N__17369),
            .I(N__17354));
    InMux I__3692 (
            .O(N__17368),
            .I(N__17349));
    InMux I__3691 (
            .O(N__17367),
            .I(N__17349));
    LocalMux I__3690 (
            .O(N__17364),
            .I(N__17346));
    InMux I__3689 (
            .O(N__17363),
            .I(N__17343));
    LocalMux I__3688 (
            .O(N__17360),
            .I(\c0.rx.r_SM_Main_2_N_816_2 ));
    LocalMux I__3687 (
            .O(N__17357),
            .I(\c0.rx.r_SM_Main_2_N_816_2 ));
    Odrv4 I__3686 (
            .O(N__17354),
            .I(\c0.rx.r_SM_Main_2_N_816_2 ));
    LocalMux I__3685 (
            .O(N__17349),
            .I(\c0.rx.r_SM_Main_2_N_816_2 ));
    Odrv4 I__3684 (
            .O(N__17346),
            .I(\c0.rx.r_SM_Main_2_N_816_2 ));
    LocalMux I__3683 (
            .O(N__17343),
            .I(\c0.rx.r_SM_Main_2_N_816_2 ));
    SRMux I__3682 (
            .O(N__17330),
            .I(N__17327));
    LocalMux I__3681 (
            .O(N__17327),
            .I(N__17324));
    Odrv4 I__3680 (
            .O(N__17324),
            .I(\c0.rx.n1024 ));
    InMux I__3679 (
            .O(N__17321),
            .I(N__17318));
    LocalMux I__3678 (
            .O(N__17318),
            .I(\c0.tx.o_Tx_Serial_N_790 ));
    InMux I__3677 (
            .O(N__17315),
            .I(N__17312));
    LocalMux I__3676 (
            .O(N__17312),
            .I(\c0.tx.n12 ));
    CascadeMux I__3675 (
            .O(N__17309),
            .I(\c0.rx.n6_cascade_ ));
    InMux I__3674 (
            .O(N__17306),
            .I(N__17297));
    InMux I__3673 (
            .O(N__17305),
            .I(N__17297));
    InMux I__3672 (
            .O(N__17304),
            .I(N__17297));
    LocalMux I__3671 (
            .O(N__17297),
            .I(\c0.rx.n357 ));
    InMux I__3670 (
            .O(N__17294),
            .I(N__17291));
    LocalMux I__3669 (
            .O(N__17291),
            .I(N__17288));
    Span4Mux_h I__3668 (
            .O(N__17288),
            .I(N__17284));
    InMux I__3667 (
            .O(N__17287),
            .I(N__17281));
    Odrv4 I__3666 (
            .O(N__17284),
            .I(rx_data_1));
    LocalMux I__3665 (
            .O(N__17281),
            .I(rx_data_1));
    CascadeMux I__3664 (
            .O(N__17276),
            .I(N__17273));
    InMux I__3663 (
            .O(N__17273),
            .I(N__17269));
    InMux I__3662 (
            .O(N__17272),
            .I(N__17266));
    LocalMux I__3661 (
            .O(N__17269),
            .I(N__17262));
    LocalMux I__3660 (
            .O(N__17266),
            .I(N__17258));
    InMux I__3659 (
            .O(N__17265),
            .I(N__17255));
    Span4Mux_v I__3658 (
            .O(N__17262),
            .I(N__17252));
    InMux I__3657 (
            .O(N__17261),
            .I(N__17249));
    Span4Mux_h I__3656 (
            .O(N__17258),
            .I(N__17242));
    LocalMux I__3655 (
            .O(N__17255),
            .I(N__17242));
    Span4Mux_s2_v I__3654 (
            .O(N__17252),
            .I(N__17242));
    LocalMux I__3653 (
            .O(N__17249),
            .I(data_in_7_1));
    Odrv4 I__3652 (
            .O(N__17242),
            .I(data_in_7_1));
    InMux I__3651 (
            .O(N__17237),
            .I(N__17233));
    InMux I__3650 (
            .O(N__17236),
            .I(N__17230));
    LocalMux I__3649 (
            .O(N__17233),
            .I(N__17227));
    LocalMux I__3648 (
            .O(N__17230),
            .I(r_Tx_Data_1));
    Odrv4 I__3647 (
            .O(N__17227),
            .I(r_Tx_Data_1));
    InMux I__3646 (
            .O(N__17222),
            .I(N__17218));
    InMux I__3645 (
            .O(N__17221),
            .I(N__17215));
    LocalMux I__3644 (
            .O(N__17218),
            .I(N__17212));
    LocalMux I__3643 (
            .O(N__17215),
            .I(r_Tx_Data_0));
    Odrv4 I__3642 (
            .O(N__17212),
            .I(r_Tx_Data_0));
    InMux I__3641 (
            .O(N__17207),
            .I(N__17203));
    InMux I__3640 (
            .O(N__17206),
            .I(N__17200));
    LocalMux I__3639 (
            .O(N__17203),
            .I(N__17197));
    LocalMux I__3638 (
            .O(N__17200),
            .I(r_Tx_Data_3));
    Odrv12 I__3637 (
            .O(N__17197),
            .I(r_Tx_Data_3));
    InMux I__3636 (
            .O(N__17192),
            .I(N__17188));
    InMux I__3635 (
            .O(N__17191),
            .I(N__17185));
    LocalMux I__3634 (
            .O(N__17188),
            .I(N__17182));
    LocalMux I__3633 (
            .O(N__17185),
            .I(r_Tx_Data_2));
    Odrv4 I__3632 (
            .O(N__17182),
            .I(r_Tx_Data_2));
    InMux I__3631 (
            .O(N__17177),
            .I(N__17174));
    LocalMux I__3630 (
            .O(N__17174),
            .I(\c0.tx.n4558 ));
    CascadeMux I__3629 (
            .O(N__17171),
            .I(\c0.tx.n4559_cascade_ ));
    InMux I__3628 (
            .O(N__17168),
            .I(N__17165));
    LocalMux I__3627 (
            .O(N__17165),
            .I(\c0.tx.n4837 ));
    IoInMux I__3626 (
            .O(N__17162),
            .I(N__17159));
    LocalMux I__3625 (
            .O(N__17159),
            .I(N__17155));
    InMux I__3624 (
            .O(N__17158),
            .I(N__17152));
    Span4Mux_s1_v I__3623 (
            .O(N__17155),
            .I(N__17149));
    LocalMux I__3622 (
            .O(N__17152),
            .I(N__17146));
    Sp12to4 I__3621 (
            .O(N__17149),
            .I(N__17142));
    Span4Mux_s1_v I__3620 (
            .O(N__17146),
            .I(N__17139));
    InMux I__3619 (
            .O(N__17145),
            .I(N__17136));
    Odrv12 I__3618 (
            .O(N__17142),
            .I(tx_o));
    Odrv4 I__3617 (
            .O(N__17139),
            .I(tx_o));
    LocalMux I__3616 (
            .O(N__17136),
            .I(tx_o));
    InMux I__3615 (
            .O(N__17129),
            .I(N__17121));
    InMux I__3614 (
            .O(N__17128),
            .I(N__17121));
    CascadeMux I__3613 (
            .O(N__17127),
            .I(N__17117));
    InMux I__3612 (
            .O(N__17126),
            .I(N__17113));
    LocalMux I__3611 (
            .O(N__17121),
            .I(N__17110));
    InMux I__3610 (
            .O(N__17120),
            .I(N__17103));
    InMux I__3609 (
            .O(N__17117),
            .I(N__17103));
    InMux I__3608 (
            .O(N__17116),
            .I(N__17103));
    LocalMux I__3607 (
            .O(N__17113),
            .I(N__17080));
    Span4Mux_h I__3606 (
            .O(N__17110),
            .I(N__17080));
    LocalMux I__3605 (
            .O(N__17103),
            .I(N__17080));
    InMux I__3604 (
            .O(N__17102),
            .I(N__17075));
    InMux I__3603 (
            .O(N__17101),
            .I(N__17075));
    InMux I__3602 (
            .O(N__17100),
            .I(N__17070));
    InMux I__3601 (
            .O(N__17099),
            .I(N__17070));
    CascadeMux I__3600 (
            .O(N__17098),
            .I(N__17066));
    InMux I__3599 (
            .O(N__17097),
            .I(N__17053));
    InMux I__3598 (
            .O(N__17096),
            .I(N__17050));
    InMux I__3597 (
            .O(N__17095),
            .I(N__17046));
    InMux I__3596 (
            .O(N__17094),
            .I(N__17041));
    InMux I__3595 (
            .O(N__17093),
            .I(N__17041));
    InMux I__3594 (
            .O(N__17092),
            .I(N__17038));
    InMux I__3593 (
            .O(N__17091),
            .I(N__17033));
    InMux I__3592 (
            .O(N__17090),
            .I(N__17033));
    InMux I__3591 (
            .O(N__17089),
            .I(N__17028));
    InMux I__3590 (
            .O(N__17088),
            .I(N__17028));
    InMux I__3589 (
            .O(N__17087),
            .I(N__17025));
    Span4Mux_v I__3588 (
            .O(N__17080),
            .I(N__17012));
    LocalMux I__3587 (
            .O(N__17075),
            .I(N__17012));
    LocalMux I__3586 (
            .O(N__17070),
            .I(N__17012));
    InMux I__3585 (
            .O(N__17069),
            .I(N__17003));
    InMux I__3584 (
            .O(N__17066),
            .I(N__17003));
    InMux I__3583 (
            .O(N__17065),
            .I(N__17003));
    InMux I__3582 (
            .O(N__17064),
            .I(N__17003));
    InMux I__3581 (
            .O(N__17063),
            .I(N__16989));
    InMux I__3580 (
            .O(N__17062),
            .I(N__16989));
    InMux I__3579 (
            .O(N__17061),
            .I(N__16989));
    InMux I__3578 (
            .O(N__17060),
            .I(N__16974));
    InMux I__3577 (
            .O(N__17059),
            .I(N__16974));
    InMux I__3576 (
            .O(N__17058),
            .I(N__16974));
    InMux I__3575 (
            .O(N__17057),
            .I(N__16974));
    InMux I__3574 (
            .O(N__17056),
            .I(N__16974));
    LocalMux I__3573 (
            .O(N__17053),
            .I(N__16965));
    LocalMux I__3572 (
            .O(N__17050),
            .I(N__16965));
    InMux I__3571 (
            .O(N__17049),
            .I(N__16962));
    LocalMux I__3570 (
            .O(N__17046),
            .I(N__16957));
    LocalMux I__3569 (
            .O(N__17041),
            .I(N__16957));
    LocalMux I__3568 (
            .O(N__17038),
            .I(N__16954));
    LocalMux I__3567 (
            .O(N__17033),
            .I(N__16951));
    LocalMux I__3566 (
            .O(N__17028),
            .I(N__16946));
    LocalMux I__3565 (
            .O(N__17025),
            .I(N__16946));
    InMux I__3564 (
            .O(N__17024),
            .I(N__16943));
    InMux I__3563 (
            .O(N__17023),
            .I(N__16940));
    InMux I__3562 (
            .O(N__17022),
            .I(N__16937));
    InMux I__3561 (
            .O(N__17021),
            .I(N__16932));
    InMux I__3560 (
            .O(N__17020),
            .I(N__16932));
    InMux I__3559 (
            .O(N__17019),
            .I(N__16929));
    Span4Mux_s1_v I__3558 (
            .O(N__17012),
            .I(N__16924));
    LocalMux I__3557 (
            .O(N__17003),
            .I(N__16924));
    InMux I__3556 (
            .O(N__17002),
            .I(N__16908));
    InMux I__3555 (
            .O(N__17001),
            .I(N__16908));
    InMux I__3554 (
            .O(N__17000),
            .I(N__16908));
    InMux I__3553 (
            .O(N__16999),
            .I(N__16908));
    InMux I__3552 (
            .O(N__16998),
            .I(N__16902));
    InMux I__3551 (
            .O(N__16997),
            .I(N__16899));
    InMux I__3550 (
            .O(N__16996),
            .I(N__16896));
    LocalMux I__3549 (
            .O(N__16989),
            .I(N__16893));
    InMux I__3548 (
            .O(N__16988),
            .I(N__16884));
    InMux I__3547 (
            .O(N__16987),
            .I(N__16884));
    InMux I__3546 (
            .O(N__16986),
            .I(N__16884));
    InMux I__3545 (
            .O(N__16985),
            .I(N__16884));
    LocalMux I__3544 (
            .O(N__16974),
            .I(N__16881));
    InMux I__3543 (
            .O(N__16973),
            .I(N__16874));
    InMux I__3542 (
            .O(N__16972),
            .I(N__16874));
    InMux I__3541 (
            .O(N__16971),
            .I(N__16874));
    InMux I__3540 (
            .O(N__16970),
            .I(N__16871));
    Span4Mux_v I__3539 (
            .O(N__16965),
            .I(N__16866));
    LocalMux I__3538 (
            .O(N__16962),
            .I(N__16866));
    Span4Mux_s2_v I__3537 (
            .O(N__16957),
            .I(N__16863));
    Span4Mux_h I__3536 (
            .O(N__16954),
            .I(N__16856));
    Span4Mux_h I__3535 (
            .O(N__16951),
            .I(N__16856));
    Span4Mux_v I__3534 (
            .O(N__16946),
            .I(N__16856));
    LocalMux I__3533 (
            .O(N__16943),
            .I(N__16843));
    LocalMux I__3532 (
            .O(N__16940),
            .I(N__16843));
    LocalMux I__3531 (
            .O(N__16937),
            .I(N__16843));
    LocalMux I__3530 (
            .O(N__16932),
            .I(N__16843));
    LocalMux I__3529 (
            .O(N__16929),
            .I(N__16843));
    Sp12to4 I__3528 (
            .O(N__16924),
            .I(N__16843));
    InMux I__3527 (
            .O(N__16923),
            .I(N__16832));
    InMux I__3526 (
            .O(N__16922),
            .I(N__16832));
    InMux I__3525 (
            .O(N__16921),
            .I(N__16832));
    InMux I__3524 (
            .O(N__16920),
            .I(N__16832));
    InMux I__3523 (
            .O(N__16919),
            .I(N__16832));
    InMux I__3522 (
            .O(N__16918),
            .I(N__16827));
    InMux I__3521 (
            .O(N__16917),
            .I(N__16827));
    LocalMux I__3520 (
            .O(N__16908),
            .I(N__16824));
    InMux I__3519 (
            .O(N__16907),
            .I(N__16821));
    InMux I__3518 (
            .O(N__16906),
            .I(N__16816));
    InMux I__3517 (
            .O(N__16905),
            .I(N__16816));
    LocalMux I__3516 (
            .O(N__16902),
            .I(N__16811));
    LocalMux I__3515 (
            .O(N__16899),
            .I(N__16811));
    LocalMux I__3514 (
            .O(N__16896),
            .I(N__16806));
    Span4Mux_v I__3513 (
            .O(N__16893),
            .I(N__16806));
    LocalMux I__3512 (
            .O(N__16884),
            .I(N__16801));
    Span4Mux_h I__3511 (
            .O(N__16881),
            .I(N__16801));
    LocalMux I__3510 (
            .O(N__16874),
            .I(N__16790));
    LocalMux I__3509 (
            .O(N__16871),
            .I(N__16790));
    Span4Mux_s2_v I__3508 (
            .O(N__16866),
            .I(N__16790));
    Span4Mux_h I__3507 (
            .O(N__16863),
            .I(N__16790));
    Span4Mux_v I__3506 (
            .O(N__16856),
            .I(N__16790));
    Span12Mux_s5_h I__3505 (
            .O(N__16843),
            .I(N__16787));
    LocalMux I__3504 (
            .O(N__16832),
            .I(N__16780));
    LocalMux I__3503 (
            .O(N__16827),
            .I(N__16780));
    Span12Mux_v I__3502 (
            .O(N__16824),
            .I(N__16780));
    LocalMux I__3501 (
            .O(N__16821),
            .I(rx_data_ready_keep));
    LocalMux I__3500 (
            .O(N__16816),
            .I(rx_data_ready_keep));
    Odrv4 I__3499 (
            .O(N__16811),
            .I(rx_data_ready_keep));
    Odrv4 I__3498 (
            .O(N__16806),
            .I(rx_data_ready_keep));
    Odrv4 I__3497 (
            .O(N__16801),
            .I(rx_data_ready_keep));
    Odrv4 I__3496 (
            .O(N__16790),
            .I(rx_data_ready_keep));
    Odrv12 I__3495 (
            .O(N__16787),
            .I(rx_data_ready_keep));
    Odrv12 I__3494 (
            .O(N__16780),
            .I(rx_data_ready_keep));
    InMux I__3493 (
            .O(N__16763),
            .I(N__16759));
    InMux I__3492 (
            .O(N__16762),
            .I(N__16756));
    LocalMux I__3491 (
            .O(N__16759),
            .I(N__16753));
    LocalMux I__3490 (
            .O(N__16756),
            .I(N__16746));
    Span4Mux_s2_v I__3489 (
            .O(N__16753),
            .I(N__16746));
    InMux I__3488 (
            .O(N__16752),
            .I(N__16743));
    InMux I__3487 (
            .O(N__16751),
            .I(N__16740));
    Odrv4 I__3486 (
            .O(N__16746),
            .I(data_in_6_1));
    LocalMux I__3485 (
            .O(N__16743),
            .I(data_in_6_1));
    LocalMux I__3484 (
            .O(N__16740),
            .I(data_in_6_1));
    InMux I__3483 (
            .O(N__16733),
            .I(N__16730));
    LocalMux I__3482 (
            .O(N__16730),
            .I(\c0.n4789 ));
    CascadeMux I__3481 (
            .O(N__16727),
            .I(tx_data_4_keep_cascade_));
    InMux I__3480 (
            .O(N__16724),
            .I(N__16720));
    InMux I__3479 (
            .O(N__16723),
            .I(N__16717));
    LocalMux I__3478 (
            .O(N__16720),
            .I(r_Tx_Data_4));
    LocalMux I__3477 (
            .O(N__16717),
            .I(r_Tx_Data_4));
    InMux I__3476 (
            .O(N__16712),
            .I(N__16709));
    LocalMux I__3475 (
            .O(N__16709),
            .I(\c0.n4576 ));
    InMux I__3474 (
            .O(N__16706),
            .I(N__16703));
    LocalMux I__3473 (
            .O(N__16703),
            .I(N__16700));
    Odrv4 I__3472 (
            .O(N__16700),
            .I(\c0.tx.n4589 ));
    InMux I__3471 (
            .O(N__16697),
            .I(N__16694));
    LocalMux I__3470 (
            .O(N__16694),
            .I(\c0.tx.n4588 ));
    CascadeMux I__3469 (
            .O(N__16691),
            .I(tx_data_5_keep_cascade_));
    InMux I__3468 (
            .O(N__16688),
            .I(N__16684));
    InMux I__3467 (
            .O(N__16687),
            .I(N__16681));
    LocalMux I__3466 (
            .O(N__16684),
            .I(r_Tx_Data_5));
    LocalMux I__3465 (
            .O(N__16681),
            .I(r_Tx_Data_5));
    CascadeMux I__3464 (
            .O(N__16676),
            .I(N__16672));
    InMux I__3463 (
            .O(N__16675),
            .I(N__16667));
    InMux I__3462 (
            .O(N__16672),
            .I(N__16667));
    LocalMux I__3461 (
            .O(N__16667),
            .I(N__16664));
    Odrv12 I__3460 (
            .O(N__16664),
            .I(\c0.tx.n1588 ));
    CascadeMux I__3459 (
            .O(N__16661),
            .I(\c0.tx.n4715_cascade_ ));
    InMux I__3458 (
            .O(N__16658),
            .I(N__16654));
    InMux I__3457 (
            .O(N__16657),
            .I(N__16651));
    LocalMux I__3456 (
            .O(N__16654),
            .I(r_Tx_Data_7));
    LocalMux I__3455 (
            .O(N__16651),
            .I(r_Tx_Data_7));
    InMux I__3454 (
            .O(N__16646),
            .I(N__16643));
    LocalMux I__3453 (
            .O(N__16643),
            .I(\c0.n4585 ));
    InMux I__3452 (
            .O(N__16640),
            .I(N__16634));
    InMux I__3451 (
            .O(N__16639),
            .I(N__16634));
    LocalMux I__3450 (
            .O(N__16634),
            .I(r_Tx_Data_6));
    CascadeMux I__3449 (
            .O(N__16631),
            .I(\c0.n4861_cascade_ ));
    CascadeMux I__3448 (
            .O(N__16628),
            .I(tx_data_0_keep_cascade_));
    CascadeMux I__3447 (
            .O(N__16625),
            .I(N__16622));
    InMux I__3446 (
            .O(N__16622),
            .I(N__16619));
    LocalMux I__3445 (
            .O(N__16619),
            .I(\c0.n4586 ));
    InMux I__3444 (
            .O(N__16616),
            .I(N__16613));
    LocalMux I__3443 (
            .O(N__16613),
            .I(N__16610));
    Odrv4 I__3442 (
            .O(N__16610),
            .I(\c0.n4573 ));
    InMux I__3441 (
            .O(N__16607),
            .I(N__16604));
    LocalMux I__3440 (
            .O(N__16604),
            .I(\c0.n4621 ));
    InMux I__3439 (
            .O(N__16601),
            .I(N__16598));
    LocalMux I__3438 (
            .O(N__16598),
            .I(\c0.n4525 ));
    InMux I__3437 (
            .O(N__16595),
            .I(N__16592));
    LocalMux I__3436 (
            .O(N__16592),
            .I(N__16588));
    InMux I__3435 (
            .O(N__16591),
            .I(N__16585));
    Span4Mux_s2_v I__3434 (
            .O(N__16588),
            .I(N__16582));
    LocalMux I__3433 (
            .O(N__16585),
            .I(N__16579));
    Span4Mux_h I__3432 (
            .O(N__16582),
            .I(N__16572));
    Span4Mux_h I__3431 (
            .O(N__16579),
            .I(N__16572));
    InMux I__3430 (
            .O(N__16578),
            .I(N__16567));
    InMux I__3429 (
            .O(N__16577),
            .I(N__16567));
    Odrv4 I__3428 (
            .O(N__16572),
            .I(data_in_6_3));
    LocalMux I__3427 (
            .O(N__16567),
            .I(data_in_6_3));
    InMux I__3426 (
            .O(N__16562),
            .I(N__16558));
    InMux I__3425 (
            .O(N__16561),
            .I(N__16555));
    LocalMux I__3424 (
            .O(N__16558),
            .I(N__16552));
    LocalMux I__3423 (
            .O(N__16555),
            .I(N__16549));
    Span12Mux_s6_h I__3422 (
            .O(N__16552),
            .I(N__16545));
    Span4Mux_h I__3421 (
            .O(N__16549),
            .I(N__16542));
    InMux I__3420 (
            .O(N__16548),
            .I(N__16539));
    Odrv12 I__3419 (
            .O(N__16545),
            .I(data_in_5_3));
    Odrv4 I__3418 (
            .O(N__16542),
            .I(data_in_5_3));
    LocalMux I__3417 (
            .O(N__16539),
            .I(data_in_5_3));
    CascadeMux I__3416 (
            .O(N__16532),
            .I(\c0.n4768_cascade_ ));
    CascadeMux I__3415 (
            .O(N__16529),
            .I(tx_data_7_keep_cascade_));
    CascadeMux I__3414 (
            .O(N__16526),
            .I(\c0.n4843_cascade_ ));
    CascadeMux I__3413 (
            .O(N__16523),
            .I(tx_data_1_keep_cascade_));
    CascadeMux I__3412 (
            .O(N__16520),
            .I(\c0.rx.n4641_cascade_ ));
    InMux I__3411 (
            .O(N__16517),
            .I(N__16514));
    LocalMux I__3410 (
            .O(N__16514),
            .I(\c0.rx.n8 ));
    InMux I__3409 (
            .O(N__16511),
            .I(N__16508));
    LocalMux I__3408 (
            .O(N__16508),
            .I(\c0.rx.n4 ));
    CascadeMux I__3407 (
            .O(N__16505),
            .I(N__16502));
    InMux I__3406 (
            .O(N__16502),
            .I(N__16499));
    LocalMux I__3405 (
            .O(N__16499),
            .I(N__16496));
    Odrv12 I__3404 (
            .O(N__16496),
            .I(\c0.rx.n7 ));
    CascadeMux I__3403 (
            .O(N__16493),
            .I(\c0.rx.n4093_cascade_ ));
    InMux I__3402 (
            .O(N__16490),
            .I(N__16487));
    LocalMux I__3401 (
            .O(N__16487),
            .I(\c0.rx.n2246 ));
    CascadeMux I__3400 (
            .O(N__16484),
            .I(N__16481));
    InMux I__3399 (
            .O(N__16481),
            .I(N__16478));
    LocalMux I__3398 (
            .O(N__16478),
            .I(n221));
    InMux I__3397 (
            .O(N__16475),
            .I(N__16470));
    InMux I__3396 (
            .O(N__16474),
            .I(N__16467));
    InMux I__3395 (
            .O(N__16473),
            .I(N__16464));
    LocalMux I__3394 (
            .O(N__16470),
            .I(r_Clock_Count_5));
    LocalMux I__3393 (
            .O(N__16467),
            .I(r_Clock_Count_5));
    LocalMux I__3392 (
            .O(N__16464),
            .I(r_Clock_Count_5));
    CascadeMux I__3391 (
            .O(N__16457),
            .I(\c0.n4783_cascade_ ));
    InMux I__3390 (
            .O(N__16454),
            .I(N__16451));
    LocalMux I__3389 (
            .O(N__16451),
            .I(N__16448));
    Span4Mux_v I__3388 (
            .O(N__16448),
            .I(N__16445));
    Odrv4 I__3387 (
            .O(N__16445),
            .I(\c0.n4526 ));
    CascadeMux I__3386 (
            .O(N__16442),
            .I(tx_data_3_keep_cascade_));
    CascadeMux I__3385 (
            .O(N__16439),
            .I(N__16436));
    InMux I__3384 (
            .O(N__16436),
            .I(N__16433));
    LocalMux I__3383 (
            .O(N__16433),
            .I(\c0.n4622 ));
    InMux I__3382 (
            .O(N__16430),
            .I(N__16425));
    InMux I__3381 (
            .O(N__16429),
            .I(N__16421));
    InMux I__3380 (
            .O(N__16428),
            .I(N__16418));
    LocalMux I__3379 (
            .O(N__16425),
            .I(N__16415));
    InMux I__3378 (
            .O(N__16424),
            .I(N__16412));
    LocalMux I__3377 (
            .O(N__16421),
            .I(r_Clock_Count_3));
    LocalMux I__3376 (
            .O(N__16418),
            .I(r_Clock_Count_3));
    Odrv4 I__3375 (
            .O(N__16415),
            .I(r_Clock_Count_3));
    LocalMux I__3374 (
            .O(N__16412),
            .I(r_Clock_Count_3));
    CascadeMux I__3373 (
            .O(N__16403),
            .I(\c0.rx.n214_cascade_ ));
    CascadeMux I__3372 (
            .O(N__16400),
            .I(\c0.rx.n4_cascade_ ));
    InMux I__3371 (
            .O(N__16397),
            .I(N__16388));
    InMux I__3370 (
            .O(N__16396),
            .I(N__16383));
    InMux I__3369 (
            .O(N__16395),
            .I(N__16383));
    InMux I__3368 (
            .O(N__16394),
            .I(N__16378));
    InMux I__3367 (
            .O(N__16393),
            .I(N__16378));
    InMux I__3366 (
            .O(N__16392),
            .I(N__16373));
    InMux I__3365 (
            .O(N__16391),
            .I(N__16373));
    LocalMux I__3364 (
            .O(N__16388),
            .I(r_Bit_Index_2));
    LocalMux I__3363 (
            .O(N__16383),
            .I(r_Bit_Index_2));
    LocalMux I__3362 (
            .O(N__16378),
            .I(r_Bit_Index_2));
    LocalMux I__3361 (
            .O(N__16373),
            .I(r_Bit_Index_2));
    InMux I__3360 (
            .O(N__16364),
            .I(N__16355));
    InMux I__3359 (
            .O(N__16363),
            .I(N__16352));
    InMux I__3358 (
            .O(N__16362),
            .I(N__16349));
    InMux I__3357 (
            .O(N__16361),
            .I(N__16344));
    InMux I__3356 (
            .O(N__16360),
            .I(N__16344));
    InMux I__3355 (
            .O(N__16359),
            .I(N__16339));
    InMux I__3354 (
            .O(N__16358),
            .I(N__16339));
    LocalMux I__3353 (
            .O(N__16355),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__3352 (
            .O(N__16352),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__3351 (
            .O(N__16349),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__3350 (
            .O(N__16344),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__3349 (
            .O(N__16339),
            .I(\c0.rx.r_Bit_Index_1 ));
    InMux I__3348 (
            .O(N__16328),
            .I(N__16322));
    InMux I__3347 (
            .O(N__16327),
            .I(N__16322));
    LocalMux I__3346 (
            .O(N__16322),
            .I(N__16319));
    Odrv4 I__3345 (
            .O(N__16319),
            .I(n4_adj_951));
    InMux I__3344 (
            .O(N__16316),
            .I(N__16313));
    LocalMux I__3343 (
            .O(N__16313),
            .I(\c0.rx.n4679 ));
    CascadeMux I__3342 (
            .O(N__16310),
            .I(N__16307));
    InMux I__3341 (
            .O(N__16307),
            .I(N__16301));
    InMux I__3340 (
            .O(N__16306),
            .I(N__16298));
    InMux I__3339 (
            .O(N__16305),
            .I(N__16293));
    InMux I__3338 (
            .O(N__16304),
            .I(N__16293));
    LocalMux I__3337 (
            .O(N__16301),
            .I(N__16290));
    LocalMux I__3336 (
            .O(N__16298),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__3335 (
            .O(N__16293),
            .I(\c0.rx.r_Clock_Count_1 ));
    Odrv12 I__3334 (
            .O(N__16290),
            .I(\c0.rx.r_Clock_Count_1 ));
    InMux I__3333 (
            .O(N__16283),
            .I(N__16280));
    LocalMux I__3332 (
            .O(N__16280),
            .I(n219));
    InMux I__3331 (
            .O(N__16277),
            .I(N__16274));
    LocalMux I__3330 (
            .O(N__16274),
            .I(N__16267));
    InMux I__3329 (
            .O(N__16273),
            .I(N__16264));
    InMux I__3328 (
            .O(N__16272),
            .I(N__16261));
    InMux I__3327 (
            .O(N__16271),
            .I(N__16256));
    InMux I__3326 (
            .O(N__16270),
            .I(N__16256));
    Odrv4 I__3325 (
            .O(N__16267),
            .I(r_Clock_Count_7));
    LocalMux I__3324 (
            .O(N__16264),
            .I(r_Clock_Count_7));
    LocalMux I__3323 (
            .O(N__16261),
            .I(r_Clock_Count_7));
    LocalMux I__3322 (
            .O(N__16256),
            .I(r_Clock_Count_7));
    InMux I__3321 (
            .O(N__16247),
            .I(N__16244));
    LocalMux I__3320 (
            .O(N__16244),
            .I(N__16241));
    Odrv12 I__3319 (
            .O(N__16241),
            .I(\c0.rx.n4677 ));
    InMux I__3318 (
            .O(N__16238),
            .I(N__16235));
    LocalMux I__3317 (
            .O(N__16235),
            .I(N__16232));
    Odrv4 I__3316 (
            .O(N__16232),
            .I(n226));
    CascadeMux I__3315 (
            .O(N__16229),
            .I(n573_cascade_));
    CascadeMux I__3314 (
            .O(N__16226),
            .I(N__16221));
    InMux I__3313 (
            .O(N__16225),
            .I(N__16218));
    InMux I__3312 (
            .O(N__16224),
            .I(N__16214));
    InMux I__3311 (
            .O(N__16221),
            .I(N__16211));
    LocalMux I__3310 (
            .O(N__16218),
            .I(N__16208));
    InMux I__3309 (
            .O(N__16217),
            .I(N__16205));
    LocalMux I__3308 (
            .O(N__16214),
            .I(r_Clock_Count_0));
    LocalMux I__3307 (
            .O(N__16211),
            .I(r_Clock_Count_0));
    Odrv4 I__3306 (
            .O(N__16208),
            .I(r_Clock_Count_0));
    LocalMux I__3305 (
            .O(N__16205),
            .I(r_Clock_Count_0));
    CascadeMux I__3304 (
            .O(N__16196),
            .I(N__16193));
    InMux I__3303 (
            .O(N__16193),
            .I(N__16190));
    LocalMux I__3302 (
            .O(N__16190),
            .I(N__16187));
    Odrv4 I__3301 (
            .O(N__16187),
            .I(n222));
    InMux I__3300 (
            .O(N__16184),
            .I(N__16181));
    LocalMux I__3299 (
            .O(N__16181),
            .I(N__16176));
    InMux I__3298 (
            .O(N__16180),
            .I(N__16173));
    InMux I__3297 (
            .O(N__16179),
            .I(N__16170));
    Odrv4 I__3296 (
            .O(N__16176),
            .I(r_Clock_Count_4));
    LocalMux I__3295 (
            .O(N__16173),
            .I(r_Clock_Count_4));
    LocalMux I__3294 (
            .O(N__16170),
            .I(r_Clock_Count_4));
    CascadeMux I__3293 (
            .O(N__16163),
            .I(N__16159));
    InMux I__3292 (
            .O(N__16162),
            .I(N__16151));
    InMux I__3291 (
            .O(N__16159),
            .I(N__16151));
    InMux I__3290 (
            .O(N__16158),
            .I(N__16151));
    LocalMux I__3289 (
            .O(N__16151),
            .I(n1527));
    CascadeMux I__3288 (
            .O(N__16148),
            .I(n1527_cascade_));
    InMux I__3287 (
            .O(N__16145),
            .I(N__16136));
    InMux I__3286 (
            .O(N__16144),
            .I(N__16136));
    InMux I__3285 (
            .O(N__16143),
            .I(N__16136));
    LocalMux I__3284 (
            .O(N__16136),
            .I(n2142));
    CascadeMux I__3283 (
            .O(N__16133),
            .I(N__16128));
    CascadeMux I__3282 (
            .O(N__16132),
            .I(N__16125));
    InMux I__3281 (
            .O(N__16131),
            .I(N__16122));
    InMux I__3280 (
            .O(N__16128),
            .I(N__16119));
    InMux I__3279 (
            .O(N__16125),
            .I(N__16115));
    LocalMux I__3278 (
            .O(N__16122),
            .I(N__16112));
    LocalMux I__3277 (
            .O(N__16119),
            .I(N__16109));
    InMux I__3276 (
            .O(N__16118),
            .I(N__16106));
    LocalMux I__3275 (
            .O(N__16115),
            .I(N__16103));
    Span4Mux_h I__3274 (
            .O(N__16112),
            .I(N__16100));
    Span4Mux_h I__3273 (
            .O(N__16109),
            .I(N__16097));
    LocalMux I__3272 (
            .O(N__16106),
            .I(data_in_7_0));
    Odrv4 I__3271 (
            .O(N__16103),
            .I(data_in_7_0));
    Odrv4 I__3270 (
            .O(N__16100),
            .I(data_in_7_0));
    Odrv4 I__3269 (
            .O(N__16097),
            .I(data_in_7_0));
    InMux I__3268 (
            .O(N__16088),
            .I(N__16082));
    InMux I__3267 (
            .O(N__16087),
            .I(N__16079));
    InMux I__3266 (
            .O(N__16086),
            .I(N__16076));
    InMux I__3265 (
            .O(N__16085),
            .I(N__16073));
    LocalMux I__3264 (
            .O(N__16082),
            .I(N__16070));
    LocalMux I__3263 (
            .O(N__16079),
            .I(N__16067));
    LocalMux I__3262 (
            .O(N__16076),
            .I(data_in_6_0));
    LocalMux I__3261 (
            .O(N__16073),
            .I(data_in_6_0));
    Odrv12 I__3260 (
            .O(N__16070),
            .I(data_in_6_0));
    Odrv4 I__3259 (
            .O(N__16067),
            .I(data_in_6_0));
    CascadeMux I__3258 (
            .O(N__16058),
            .I(N__16055));
    InMux I__3257 (
            .O(N__16055),
            .I(N__16052));
    LocalMux I__3256 (
            .O(N__16052),
            .I(\c0.rx.n232 ));
    CascadeMux I__3255 (
            .O(N__16049),
            .I(\c0.rx.r_SM_Main_2_N_816_2_cascade_ ));
    InMux I__3254 (
            .O(N__16046),
            .I(N__16043));
    LocalMux I__3253 (
            .O(N__16043),
            .I(N__16040));
    Span4Mux_s2_v I__3252 (
            .O(N__16040),
            .I(N__16037));
    Odrv4 I__3251 (
            .O(N__16037),
            .I(\c0.rx.n4678 ));
    CascadeMux I__3250 (
            .O(N__16034),
            .I(N__16028));
    InMux I__3249 (
            .O(N__16033),
            .I(N__16021));
    InMux I__3248 (
            .O(N__16032),
            .I(N__16021));
    InMux I__3247 (
            .O(N__16031),
            .I(N__16016));
    InMux I__3246 (
            .O(N__16028),
            .I(N__16016));
    InMux I__3245 (
            .O(N__16027),
            .I(N__16011));
    InMux I__3244 (
            .O(N__16026),
            .I(N__16011));
    LocalMux I__3243 (
            .O(N__16021),
            .I(r_Bit_Index_0));
    LocalMux I__3242 (
            .O(N__16016),
            .I(r_Bit_Index_0));
    LocalMux I__3241 (
            .O(N__16011),
            .I(r_Bit_Index_0));
    CascadeMux I__3240 (
            .O(N__16004),
            .I(N__16001));
    InMux I__3239 (
            .O(N__16001),
            .I(N__15997));
    InMux I__3238 (
            .O(N__16000),
            .I(N__15994));
    LocalMux I__3237 (
            .O(N__15997),
            .I(n4_adj_943));
    LocalMux I__3236 (
            .O(N__15994),
            .I(n4_adj_943));
    CascadeMux I__3235 (
            .O(N__15989),
            .I(N__15986));
    InMux I__3234 (
            .O(N__15986),
            .I(N__15983));
    LocalMux I__3233 (
            .O(N__15983),
            .I(N__15980));
    Odrv4 I__3232 (
            .O(N__15980),
            .I(n223));
    InMux I__3231 (
            .O(N__15977),
            .I(N__15974));
    LocalMux I__3230 (
            .O(N__15974),
            .I(N__15970));
    InMux I__3229 (
            .O(N__15973),
            .I(N__15967));
    Odrv4 I__3228 (
            .O(N__15970),
            .I(\c0.rx.n214 ));
    LocalMux I__3227 (
            .O(N__15967),
            .I(\c0.rx.n214 ));
    InMux I__3226 (
            .O(N__15962),
            .I(N__15959));
    LocalMux I__3225 (
            .O(N__15959),
            .I(N__15956));
    Span4Mux_h I__3224 (
            .O(N__15956),
            .I(N__15953));
    Odrv4 I__3223 (
            .O(N__15953),
            .I(\c0.n4408 ));
    InMux I__3222 (
            .O(N__15950),
            .I(N__15947));
    LocalMux I__3221 (
            .O(N__15947),
            .I(N__15944));
    Span4Mux_h I__3220 (
            .O(N__15944),
            .I(N__15940));
    InMux I__3219 (
            .O(N__15943),
            .I(N__15937));
    Odrv4 I__3218 (
            .O(N__15940),
            .I(\c0.n1271 ));
    LocalMux I__3217 (
            .O(N__15937),
            .I(\c0.n1271 ));
    InMux I__3216 (
            .O(N__15932),
            .I(N__15929));
    LocalMux I__3215 (
            .O(N__15929),
            .I(N__15926));
    Span4Mux_h I__3214 (
            .O(N__15926),
            .I(N__15923));
    Odrv4 I__3213 (
            .O(N__15923),
            .I(\c0.n4409 ));
    CascadeMux I__3212 (
            .O(N__15920),
            .I(\c0.rx.n232_cascade_ ));
    InMux I__3211 (
            .O(N__15917),
            .I(N__15914));
    LocalMux I__3210 (
            .O(N__15914),
            .I(N__15911));
    Odrv4 I__3209 (
            .O(N__15911),
            .I(\c0.n4516 ));
    CascadeMux I__3208 (
            .O(N__15908),
            .I(\c0.rx.n1464_cascade_ ));
    CascadeMux I__3207 (
            .O(N__15905),
            .I(N__15902));
    InMux I__3206 (
            .O(N__15902),
            .I(N__15899));
    LocalMux I__3205 (
            .O(N__15899),
            .I(N__15895));
    InMux I__3204 (
            .O(N__15898),
            .I(N__15892));
    Odrv4 I__3203 (
            .O(N__15895),
            .I(\c0.data_1 ));
    LocalMux I__3202 (
            .O(N__15892),
            .I(\c0.data_1 ));
    InMux I__3201 (
            .O(N__15887),
            .I(N__15884));
    LocalMux I__3200 (
            .O(N__15884),
            .I(N__15879));
    CascadeMux I__3199 (
            .O(N__15883),
            .I(N__15875));
    InMux I__3198 (
            .O(N__15882),
            .I(N__15872));
    Span4Mux_h I__3197 (
            .O(N__15879),
            .I(N__15869));
    InMux I__3196 (
            .O(N__15878),
            .I(N__15866));
    InMux I__3195 (
            .O(N__15875),
            .I(N__15863));
    LocalMux I__3194 (
            .O(N__15872),
            .I(data_in_7_2));
    Odrv4 I__3193 (
            .O(N__15869),
            .I(data_in_7_2));
    LocalMux I__3192 (
            .O(N__15866),
            .I(data_in_7_2));
    LocalMux I__3191 (
            .O(N__15863),
            .I(data_in_7_2));
    InMux I__3190 (
            .O(N__15854),
            .I(N__15849));
    InMux I__3189 (
            .O(N__15853),
            .I(N__15846));
    CascadeMux I__3188 (
            .O(N__15852),
            .I(N__15842));
    LocalMux I__3187 (
            .O(N__15849),
            .I(N__15839));
    LocalMux I__3186 (
            .O(N__15846),
            .I(N__15836));
    InMux I__3185 (
            .O(N__15845),
            .I(N__15833));
    InMux I__3184 (
            .O(N__15842),
            .I(N__15830));
    Span4Mux_h I__3183 (
            .O(N__15839),
            .I(N__15825));
    Span4Mux_h I__3182 (
            .O(N__15836),
            .I(N__15825));
    LocalMux I__3181 (
            .O(N__15833),
            .I(data_in_6_2));
    LocalMux I__3180 (
            .O(N__15830),
            .I(data_in_6_2));
    Odrv4 I__3179 (
            .O(N__15825),
            .I(data_in_6_2));
    CascadeMux I__3178 (
            .O(N__15818),
            .I(\c0.n4517_cascade_ ));
    CascadeMux I__3177 (
            .O(N__15815),
            .I(\c0.n4867_cascade_ ));
    CascadeMux I__3176 (
            .O(N__15812),
            .I(tx_data_2_keep_cascade_));
    InMux I__3175 (
            .O(N__15809),
            .I(N__15806));
    LocalMux I__3174 (
            .O(N__15806),
            .I(\c0.n4564 ));
    InMux I__3173 (
            .O(N__15803),
            .I(\c0.n3916 ));
    InMux I__3172 (
            .O(N__15800),
            .I(\c0.n3917 ));
    InMux I__3171 (
            .O(N__15797),
            .I(\c0.n3918 ));
    InMux I__3170 (
            .O(N__15794),
            .I(\c0.n3919 ));
    InMux I__3169 (
            .O(N__15791),
            .I(\c0.n3920 ));
    CascadeMux I__3168 (
            .O(N__15788),
            .I(N__15779));
    CascadeMux I__3167 (
            .O(N__15787),
            .I(N__15774));
    CascadeMux I__3166 (
            .O(N__15786),
            .I(N__15771));
    CascadeMux I__3165 (
            .O(N__15785),
            .I(N__15768));
    CascadeMux I__3164 (
            .O(N__15784),
            .I(N__15762));
    CascadeMux I__3163 (
            .O(N__15783),
            .I(N__15757));
    CascadeMux I__3162 (
            .O(N__15782),
            .I(N__15754));
    InMux I__3161 (
            .O(N__15779),
            .I(N__15751));
    InMux I__3160 (
            .O(N__15778),
            .I(N__15748));
    CascadeMux I__3159 (
            .O(N__15777),
            .I(N__15743));
    InMux I__3158 (
            .O(N__15774),
            .I(N__15740));
    InMux I__3157 (
            .O(N__15771),
            .I(N__15735));
    InMux I__3156 (
            .O(N__15768),
            .I(N__15735));
    InMux I__3155 (
            .O(N__15767),
            .I(N__15732));
    InMux I__3154 (
            .O(N__15766),
            .I(N__15728));
    InMux I__3153 (
            .O(N__15765),
            .I(N__15723));
    InMux I__3152 (
            .O(N__15762),
            .I(N__15723));
    InMux I__3151 (
            .O(N__15761),
            .I(N__15720));
    InMux I__3150 (
            .O(N__15760),
            .I(N__15717));
    InMux I__3149 (
            .O(N__15757),
            .I(N__15714));
    InMux I__3148 (
            .O(N__15754),
            .I(N__15711));
    LocalMux I__3147 (
            .O(N__15751),
            .I(N__15706));
    LocalMux I__3146 (
            .O(N__15748),
            .I(N__15706));
    InMux I__3145 (
            .O(N__15747),
            .I(N__15698));
    InMux I__3144 (
            .O(N__15746),
            .I(N__15698));
    InMux I__3143 (
            .O(N__15743),
            .I(N__15698));
    LocalMux I__3142 (
            .O(N__15740),
            .I(N__15693));
    LocalMux I__3141 (
            .O(N__15735),
            .I(N__15693));
    LocalMux I__3140 (
            .O(N__15732),
            .I(N__15690));
    InMux I__3139 (
            .O(N__15731),
            .I(N__15687));
    LocalMux I__3138 (
            .O(N__15728),
            .I(N__15672));
    LocalMux I__3137 (
            .O(N__15723),
            .I(N__15672));
    LocalMux I__3136 (
            .O(N__15720),
            .I(N__15672));
    LocalMux I__3135 (
            .O(N__15717),
            .I(N__15672));
    LocalMux I__3134 (
            .O(N__15714),
            .I(N__15672));
    LocalMux I__3133 (
            .O(N__15711),
            .I(N__15672));
    Span4Mux_s1_h I__3132 (
            .O(N__15706),
            .I(N__15672));
    InMux I__3131 (
            .O(N__15705),
            .I(N__15669));
    LocalMux I__3130 (
            .O(N__15698),
            .I(N__15664));
    Span4Mux_h I__3129 (
            .O(N__15693),
            .I(N__15664));
    Span4Mux_h I__3128 (
            .O(N__15690),
            .I(N__15661));
    LocalMux I__3127 (
            .O(N__15687),
            .I(N__15656));
    Span4Mux_v I__3126 (
            .O(N__15672),
            .I(N__15656));
    LocalMux I__3125 (
            .O(N__15669),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__3124 (
            .O(N__15664),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__3123 (
            .O(N__15661),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__3122 (
            .O(N__15656),
            .I(\c0.byte_transmit_counter2_2 ));
    InMux I__3121 (
            .O(N__15647),
            .I(N__15641));
    InMux I__3120 (
            .O(N__15646),
            .I(N__15641));
    LocalMux I__3119 (
            .O(N__15641),
            .I(N__15632));
    InMux I__3118 (
            .O(N__15640),
            .I(N__15629));
    InMux I__3117 (
            .O(N__15639),
            .I(N__15626));
    InMux I__3116 (
            .O(N__15638),
            .I(N__15623));
    InMux I__3115 (
            .O(N__15637),
            .I(N__15620));
    InMux I__3114 (
            .O(N__15636),
            .I(N__15617));
    InMux I__3113 (
            .O(N__15635),
            .I(N__15614));
    Span4Mux_s2_h I__3112 (
            .O(N__15632),
            .I(N__15609));
    LocalMux I__3111 (
            .O(N__15629),
            .I(N__15609));
    LocalMux I__3110 (
            .O(N__15626),
            .I(N__15605));
    LocalMux I__3109 (
            .O(N__15623),
            .I(N__15601));
    LocalMux I__3108 (
            .O(N__15620),
            .I(N__15598));
    LocalMux I__3107 (
            .O(N__15617),
            .I(N__15595));
    LocalMux I__3106 (
            .O(N__15614),
            .I(N__15590));
    Span4Mux_v I__3105 (
            .O(N__15609),
            .I(N__15590));
    InMux I__3104 (
            .O(N__15608),
            .I(N__15587));
    Span4Mux_h I__3103 (
            .O(N__15605),
            .I(N__15584));
    InMux I__3102 (
            .O(N__15604),
            .I(N__15581));
    Span4Mux_h I__3101 (
            .O(N__15601),
            .I(N__15578));
    Span4Mux_v I__3100 (
            .O(N__15598),
            .I(N__15571));
    Span4Mux_v I__3099 (
            .O(N__15595),
            .I(N__15571));
    Span4Mux_s2_h I__3098 (
            .O(N__15590),
            .I(N__15571));
    LocalMux I__3097 (
            .O(N__15587),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__3096 (
            .O(N__15584),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__3095 (
            .O(N__15581),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__3094 (
            .O(N__15578),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__3093 (
            .O(N__15571),
            .I(\c0.byte_transmit_counter2_1 ));
    InMux I__3092 (
            .O(N__15560),
            .I(N__15555));
    InMux I__3091 (
            .O(N__15559),
            .I(N__15552));
    InMux I__3090 (
            .O(N__15558),
            .I(N__15549));
    LocalMux I__3089 (
            .O(N__15555),
            .I(N__15537));
    LocalMux I__3088 (
            .O(N__15552),
            .I(N__15537));
    LocalMux I__3087 (
            .O(N__15549),
            .I(N__15537));
    InMux I__3086 (
            .O(N__15548),
            .I(N__15532));
    InMux I__3085 (
            .O(N__15547),
            .I(N__15532));
    CascadeMux I__3084 (
            .O(N__15546),
            .I(N__15529));
    InMux I__3083 (
            .O(N__15545),
            .I(N__15522));
    InMux I__3082 (
            .O(N__15544),
            .I(N__15507));
    Span4Mux_v I__3081 (
            .O(N__15537),
            .I(N__15502));
    LocalMux I__3080 (
            .O(N__15532),
            .I(N__15502));
    InMux I__3079 (
            .O(N__15529),
            .I(N__15499));
    InMux I__3078 (
            .O(N__15528),
            .I(N__15496));
    InMux I__3077 (
            .O(N__15527),
            .I(N__15492));
    InMux I__3076 (
            .O(N__15526),
            .I(N__15487));
    InMux I__3075 (
            .O(N__15525),
            .I(N__15487));
    LocalMux I__3074 (
            .O(N__15522),
            .I(N__15484));
    InMux I__3073 (
            .O(N__15521),
            .I(N__15481));
    InMux I__3072 (
            .O(N__15520),
            .I(N__15478));
    InMux I__3071 (
            .O(N__15519),
            .I(N__15475));
    InMux I__3070 (
            .O(N__15518),
            .I(N__15472));
    InMux I__3069 (
            .O(N__15517),
            .I(N__15461));
    InMux I__3068 (
            .O(N__15516),
            .I(N__15461));
    InMux I__3067 (
            .O(N__15515),
            .I(N__15454));
    InMux I__3066 (
            .O(N__15514),
            .I(N__15454));
    InMux I__3065 (
            .O(N__15513),
            .I(N__15454));
    InMux I__3064 (
            .O(N__15512),
            .I(N__15449));
    InMux I__3063 (
            .O(N__15511),
            .I(N__15449));
    InMux I__3062 (
            .O(N__15510),
            .I(N__15446));
    LocalMux I__3061 (
            .O(N__15507),
            .I(N__15443));
    Span4Mux_s3_v I__3060 (
            .O(N__15502),
            .I(N__15436));
    LocalMux I__3059 (
            .O(N__15499),
            .I(N__15436));
    LocalMux I__3058 (
            .O(N__15496),
            .I(N__15436));
    CascadeMux I__3057 (
            .O(N__15495),
            .I(N__15433));
    LocalMux I__3056 (
            .O(N__15492),
            .I(N__15427));
    LocalMux I__3055 (
            .O(N__15487),
            .I(N__15418));
    Span4Mux_v I__3054 (
            .O(N__15484),
            .I(N__15418));
    LocalMux I__3053 (
            .O(N__15481),
            .I(N__15418));
    LocalMux I__3052 (
            .O(N__15478),
            .I(N__15418));
    LocalMux I__3051 (
            .O(N__15475),
            .I(N__15413));
    LocalMux I__3050 (
            .O(N__15472),
            .I(N__15413));
    InMux I__3049 (
            .O(N__15471),
            .I(N__15410));
    InMux I__3048 (
            .O(N__15470),
            .I(N__15407));
    InMux I__3047 (
            .O(N__15469),
            .I(N__15402));
    InMux I__3046 (
            .O(N__15468),
            .I(N__15402));
    InMux I__3045 (
            .O(N__15467),
            .I(N__15397));
    InMux I__3044 (
            .O(N__15466),
            .I(N__15397));
    LocalMux I__3043 (
            .O(N__15461),
            .I(N__15390));
    LocalMux I__3042 (
            .O(N__15454),
            .I(N__15390));
    LocalMux I__3041 (
            .O(N__15449),
            .I(N__15390));
    LocalMux I__3040 (
            .O(N__15446),
            .I(N__15383));
    Span4Mux_s3_v I__3039 (
            .O(N__15443),
            .I(N__15383));
    Span4Mux_h I__3038 (
            .O(N__15436),
            .I(N__15383));
    InMux I__3037 (
            .O(N__15433),
            .I(N__15380));
    InMux I__3036 (
            .O(N__15432),
            .I(N__15377));
    InMux I__3035 (
            .O(N__15431),
            .I(N__15374));
    InMux I__3034 (
            .O(N__15430),
            .I(N__15371));
    Span4Mux_v I__3033 (
            .O(N__15427),
            .I(N__15364));
    Span4Mux_v I__3032 (
            .O(N__15418),
            .I(N__15364));
    Span4Mux_v I__3031 (
            .O(N__15413),
            .I(N__15364));
    LocalMux I__3030 (
            .O(N__15410),
            .I(N__15355));
    LocalMux I__3029 (
            .O(N__15407),
            .I(N__15355));
    LocalMux I__3028 (
            .O(N__15402),
            .I(N__15355));
    LocalMux I__3027 (
            .O(N__15397),
            .I(N__15355));
    Span4Mux_h I__3026 (
            .O(N__15390),
            .I(N__15352));
    Span4Mux_v I__3025 (
            .O(N__15383),
            .I(N__15349));
    LocalMux I__3024 (
            .O(N__15380),
            .I(\c0.byte_transmit_counter2_0 ));
    LocalMux I__3023 (
            .O(N__15377),
            .I(\c0.byte_transmit_counter2_0 ));
    LocalMux I__3022 (
            .O(N__15374),
            .I(\c0.byte_transmit_counter2_0 ));
    LocalMux I__3021 (
            .O(N__15371),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__3020 (
            .O(N__15364),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv12 I__3019 (
            .O(N__15355),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__3018 (
            .O(N__15352),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__3017 (
            .O(N__15349),
            .I(\c0.byte_transmit_counter2_0 ));
    InMux I__3016 (
            .O(N__15332),
            .I(N__15329));
    LocalMux I__3015 (
            .O(N__15329),
            .I(N__15324));
    InMux I__3014 (
            .O(N__15328),
            .I(N__15321));
    InMux I__3013 (
            .O(N__15327),
            .I(N__15318));
    Span4Mux_h I__3012 (
            .O(N__15324),
            .I(N__15315));
    LocalMux I__3011 (
            .O(N__15321),
            .I(N__15310));
    LocalMux I__3010 (
            .O(N__15318),
            .I(N__15310));
    Odrv4 I__3009 (
            .O(N__15315),
            .I(\c0.FRAME_MATCHER_wait_for_transmission_N_423 ));
    Odrv4 I__3008 (
            .O(N__15310),
            .I(\c0.FRAME_MATCHER_wait_for_transmission_N_423 ));
    CascadeMux I__3007 (
            .O(N__15305),
            .I(N__15302));
    InMux I__3006 (
            .O(N__15302),
            .I(N__15298));
    InMux I__3005 (
            .O(N__15301),
            .I(N__15295));
    LocalMux I__3004 (
            .O(N__15298),
            .I(\c0.data_9 ));
    LocalMux I__3003 (
            .O(N__15295),
            .I(\c0.data_9 ));
    CascadeMux I__3002 (
            .O(N__15290),
            .I(\c0.n4619_cascade_ ));
    InMux I__3001 (
            .O(N__15287),
            .I(\c0.n3907 ));
    InMux I__3000 (
            .O(N__15284),
            .I(\c0.n3908 ));
    InMux I__2999 (
            .O(N__15281),
            .I(\c0.n3909 ));
    InMux I__2998 (
            .O(N__15278),
            .I(\c0.n3910 ));
    InMux I__2997 (
            .O(N__15275),
            .I(\c0.n3911 ));
    InMux I__2996 (
            .O(N__15272),
            .I(\c0.n3912 ));
    InMux I__2995 (
            .O(N__15269),
            .I(bfn_6_26_0_));
    InMux I__2994 (
            .O(N__15266),
            .I(\c0.n3914 ));
    InMux I__2993 (
            .O(N__15263),
            .I(\c0.n3915 ));
    InMux I__2992 (
            .O(N__15260),
            .I(\c0.rx.n3886 ));
    InMux I__2991 (
            .O(N__15257),
            .I(\c0.rx.n3887 ));
    InMux I__2990 (
            .O(N__15254),
            .I(\c0.rx.n3888 ));
    InMux I__2989 (
            .O(N__15251),
            .I(\c0.rx.n3889 ));
    InMux I__2988 (
            .O(N__15248),
            .I(\c0.rx.n3890 ));
    InMux I__2987 (
            .O(N__15245),
            .I(N__15242));
    LocalMux I__2986 (
            .O(N__15242),
            .I(N__15239));
    Span4Mux_h I__2985 (
            .O(N__15239),
            .I(N__15236));
    Odrv4 I__2984 (
            .O(N__15236),
            .I(n1695));
    InMux I__2983 (
            .O(N__15233),
            .I(N__15230));
    LocalMux I__2982 (
            .O(N__15230),
            .I(N__15219));
    InMux I__2981 (
            .O(N__15229),
            .I(N__15208));
    InMux I__2980 (
            .O(N__15228),
            .I(N__15208));
    InMux I__2979 (
            .O(N__15227),
            .I(N__15208));
    InMux I__2978 (
            .O(N__15226),
            .I(N__15208));
    InMux I__2977 (
            .O(N__15225),
            .I(N__15208));
    InMux I__2976 (
            .O(N__15224),
            .I(N__15201));
    InMux I__2975 (
            .O(N__15223),
            .I(N__15201));
    InMux I__2974 (
            .O(N__15222),
            .I(N__15201));
    Odrv12 I__2973 (
            .O(N__15219),
            .I(n6_adj_940));
    LocalMux I__2972 (
            .O(N__15208),
            .I(n6_adj_940));
    LocalMux I__2971 (
            .O(N__15201),
            .I(n6_adj_940));
    InMux I__2970 (
            .O(N__15194),
            .I(N__15189));
    InMux I__2969 (
            .O(N__15193),
            .I(N__15186));
    InMux I__2968 (
            .O(N__15192),
            .I(N__15183));
    LocalMux I__2967 (
            .O(N__15189),
            .I(N__15178));
    LocalMux I__2966 (
            .O(N__15186),
            .I(N__15178));
    LocalMux I__2965 (
            .O(N__15183),
            .I(N__15175));
    Span4Mux_h I__2964 (
            .O(N__15178),
            .I(N__15172));
    Span4Mux_h I__2963 (
            .O(N__15175),
            .I(N__15169));
    Odrv4 I__2962 (
            .O(N__15172),
            .I(\c0.tx2.r_Clock_Count_6 ));
    Odrv4 I__2961 (
            .O(N__15169),
            .I(\c0.tx2.r_Clock_Count_6 ));
    InMux I__2960 (
            .O(N__15164),
            .I(bfn_6_25_0_));
    InMux I__2959 (
            .O(N__15161),
            .I(\c0.n3906 ));
    CascadeMux I__2958 (
            .O(N__15158),
            .I(n1222_cascade_));
    InMux I__2957 (
            .O(N__15155),
            .I(N__15151));
    InMux I__2956 (
            .O(N__15154),
            .I(N__15148));
    LocalMux I__2955 (
            .O(N__15151),
            .I(rx_data_0));
    LocalMux I__2954 (
            .O(N__15148),
            .I(rx_data_0));
    InMux I__2953 (
            .O(N__15143),
            .I(N__15139));
    InMux I__2952 (
            .O(N__15142),
            .I(N__15136));
    LocalMux I__2951 (
            .O(N__15139),
            .I(N__15131));
    LocalMux I__2950 (
            .O(N__15136),
            .I(N__15131));
    Odrv12 I__2949 (
            .O(N__15131),
            .I(n4_adj_950));
    InMux I__2948 (
            .O(N__15128),
            .I(N__15122));
    InMux I__2947 (
            .O(N__15127),
            .I(N__15122));
    LocalMux I__2946 (
            .O(N__15122),
            .I(n4));
    InMux I__2945 (
            .O(N__15119),
            .I(N__15116));
    LocalMux I__2944 (
            .O(N__15116),
            .I(\c0.rx.n2269 ));
    CascadeMux I__2943 (
            .O(N__15113),
            .I(\c0.rx.n2269_cascade_ ));
    InMux I__2942 (
            .O(N__15110),
            .I(N__15107));
    LocalMux I__2941 (
            .O(N__15107),
            .I(N__15102));
    InMux I__2940 (
            .O(N__15106),
            .I(N__15097));
    InMux I__2939 (
            .O(N__15105),
            .I(N__15097));
    Odrv4 I__2938 (
            .O(N__15102),
            .I(n1227));
    LocalMux I__2937 (
            .O(N__15097),
            .I(n1227));
    CascadeMux I__2936 (
            .O(N__15092),
            .I(n1227_cascade_));
    InMux I__2935 (
            .O(N__15089),
            .I(bfn_5_32_0_));
    InMux I__2934 (
            .O(N__15086),
            .I(\c0.rx.n3884 ));
    InMux I__2933 (
            .O(N__15083),
            .I(\c0.rx.n3885 ));
    InMux I__2932 (
            .O(N__15080),
            .I(N__15075));
    InMux I__2931 (
            .O(N__15079),
            .I(N__15072));
    InMux I__2930 (
            .O(N__15078),
            .I(N__15068));
    LocalMux I__2929 (
            .O(N__15075),
            .I(N__15065));
    LocalMux I__2928 (
            .O(N__15072),
            .I(N__15062));
    InMux I__2927 (
            .O(N__15071),
            .I(N__15059));
    LocalMux I__2926 (
            .O(N__15068),
            .I(N__15056));
    Odrv12 I__2925 (
            .O(N__15065),
            .I(data_in_1_2));
    Odrv4 I__2924 (
            .O(N__15062),
            .I(data_in_1_2));
    LocalMux I__2923 (
            .O(N__15059),
            .I(data_in_1_2));
    Odrv4 I__2922 (
            .O(N__15056),
            .I(data_in_1_2));
    CascadeMux I__2921 (
            .O(N__15047),
            .I(N__15039));
    InMux I__2920 (
            .O(N__15046),
            .I(N__15006));
    InMux I__2919 (
            .O(N__15045),
            .I(N__15001));
    InMux I__2918 (
            .O(N__15044),
            .I(N__15001));
    CascadeMux I__2917 (
            .O(N__15043),
            .I(N__14998));
    InMux I__2916 (
            .O(N__15042),
            .I(N__14994));
    InMux I__2915 (
            .O(N__15039),
            .I(N__14989));
    InMux I__2914 (
            .O(N__15038),
            .I(N__14989));
    InMux I__2913 (
            .O(N__15037),
            .I(N__14984));
    InMux I__2912 (
            .O(N__15036),
            .I(N__14984));
    InMux I__2911 (
            .O(N__15035),
            .I(N__14979));
    InMux I__2910 (
            .O(N__15034),
            .I(N__14979));
    InMux I__2909 (
            .O(N__15033),
            .I(N__14974));
    InMux I__2908 (
            .O(N__15032),
            .I(N__14965));
    InMux I__2907 (
            .O(N__15031),
            .I(N__14965));
    InMux I__2906 (
            .O(N__15030),
            .I(N__14965));
    InMux I__2905 (
            .O(N__15029),
            .I(N__14965));
    InMux I__2904 (
            .O(N__15028),
            .I(N__14953));
    InMux I__2903 (
            .O(N__15027),
            .I(N__14950));
    InMux I__2902 (
            .O(N__15026),
            .I(N__14947));
    CascadeMux I__2901 (
            .O(N__15025),
            .I(N__14941));
    InMux I__2900 (
            .O(N__15024),
            .I(N__14919));
    InMux I__2899 (
            .O(N__15023),
            .I(N__14919));
    InMux I__2898 (
            .O(N__15022),
            .I(N__14919));
    InMux I__2897 (
            .O(N__15021),
            .I(N__14919));
    InMux I__2896 (
            .O(N__15020),
            .I(N__14914));
    InMux I__2895 (
            .O(N__15019),
            .I(N__14914));
    InMux I__2894 (
            .O(N__15018),
            .I(N__14901));
    InMux I__2893 (
            .O(N__15017),
            .I(N__14901));
    InMux I__2892 (
            .O(N__15016),
            .I(N__14901));
    InMux I__2891 (
            .O(N__15015),
            .I(N__14901));
    InMux I__2890 (
            .O(N__15014),
            .I(N__14901));
    InMux I__2889 (
            .O(N__15013),
            .I(N__14901));
    InMux I__2888 (
            .O(N__15012),
            .I(N__14892));
    InMux I__2887 (
            .O(N__15011),
            .I(N__14892));
    InMux I__2886 (
            .O(N__15010),
            .I(N__14892));
    InMux I__2885 (
            .O(N__15009),
            .I(N__14892));
    LocalMux I__2884 (
            .O(N__15006),
            .I(N__14889));
    LocalMux I__2883 (
            .O(N__15001),
            .I(N__14886));
    InMux I__2882 (
            .O(N__14998),
            .I(N__14881));
    InMux I__2881 (
            .O(N__14997),
            .I(N__14881));
    LocalMux I__2880 (
            .O(N__14994),
            .I(N__14872));
    LocalMux I__2879 (
            .O(N__14989),
            .I(N__14872));
    LocalMux I__2878 (
            .O(N__14984),
            .I(N__14872));
    LocalMux I__2877 (
            .O(N__14979),
            .I(N__14872));
    InMux I__2876 (
            .O(N__14978),
            .I(N__14867));
    InMux I__2875 (
            .O(N__14977),
            .I(N__14867));
    LocalMux I__2874 (
            .O(N__14974),
            .I(N__14864));
    LocalMux I__2873 (
            .O(N__14965),
            .I(N__14861));
    InMux I__2872 (
            .O(N__14964),
            .I(N__14856));
    InMux I__2871 (
            .O(N__14963),
            .I(N__14856));
    InMux I__2870 (
            .O(N__14962),
            .I(N__14853));
    InMux I__2869 (
            .O(N__14961),
            .I(N__14850));
    InMux I__2868 (
            .O(N__14960),
            .I(N__14839));
    InMux I__2867 (
            .O(N__14959),
            .I(N__14839));
    InMux I__2866 (
            .O(N__14958),
            .I(N__14839));
    InMux I__2865 (
            .O(N__14957),
            .I(N__14839));
    InMux I__2864 (
            .O(N__14956),
            .I(N__14839));
    LocalMux I__2863 (
            .O(N__14953),
            .I(N__14836));
    LocalMux I__2862 (
            .O(N__14950),
            .I(N__14831));
    LocalMux I__2861 (
            .O(N__14947),
            .I(N__14831));
    InMux I__2860 (
            .O(N__14946),
            .I(N__14826));
    InMux I__2859 (
            .O(N__14945),
            .I(N__14826));
    InMux I__2858 (
            .O(N__14944),
            .I(N__14823));
    InMux I__2857 (
            .O(N__14941),
            .I(N__14818));
    InMux I__2856 (
            .O(N__14940),
            .I(N__14818));
    InMux I__2855 (
            .O(N__14939),
            .I(N__14811));
    InMux I__2854 (
            .O(N__14938),
            .I(N__14811));
    InMux I__2853 (
            .O(N__14937),
            .I(N__14811));
    InMux I__2852 (
            .O(N__14936),
            .I(N__14804));
    InMux I__2851 (
            .O(N__14935),
            .I(N__14804));
    InMux I__2850 (
            .O(N__14934),
            .I(N__14804));
    InMux I__2849 (
            .O(N__14933),
            .I(N__14791));
    InMux I__2848 (
            .O(N__14932),
            .I(N__14791));
    InMux I__2847 (
            .O(N__14931),
            .I(N__14791));
    InMux I__2846 (
            .O(N__14930),
            .I(N__14791));
    InMux I__2845 (
            .O(N__14929),
            .I(N__14791));
    InMux I__2844 (
            .O(N__14928),
            .I(N__14791));
    LocalMux I__2843 (
            .O(N__14919),
            .I(N__14786));
    LocalMux I__2842 (
            .O(N__14914),
            .I(N__14786));
    LocalMux I__2841 (
            .O(N__14901),
            .I(N__14777));
    LocalMux I__2840 (
            .O(N__14892),
            .I(N__14777));
    Span4Mux_s2_v I__2839 (
            .O(N__14889),
            .I(N__14777));
    Span4Mux_v I__2838 (
            .O(N__14886),
            .I(N__14777));
    LocalMux I__2837 (
            .O(N__14881),
            .I(N__14772));
    Span4Mux_h I__2836 (
            .O(N__14872),
            .I(N__14772));
    LocalMux I__2835 (
            .O(N__14867),
            .I(N__14765));
    Span4Mux_v I__2834 (
            .O(N__14864),
            .I(N__14765));
    Span4Mux_h I__2833 (
            .O(N__14861),
            .I(N__14765));
    LocalMux I__2832 (
            .O(N__14856),
            .I(N__14762));
    LocalMux I__2831 (
            .O(N__14853),
            .I(N__14751));
    LocalMux I__2830 (
            .O(N__14850),
            .I(N__14751));
    LocalMux I__2829 (
            .O(N__14839),
            .I(N__14751));
    Span4Mux_v I__2828 (
            .O(N__14836),
            .I(N__14751));
    Span4Mux_h I__2827 (
            .O(N__14831),
            .I(N__14751));
    LocalMux I__2826 (
            .O(N__14826),
            .I(\c0.n1197 ));
    LocalMux I__2825 (
            .O(N__14823),
            .I(\c0.n1197 ));
    LocalMux I__2824 (
            .O(N__14818),
            .I(\c0.n1197 ));
    LocalMux I__2823 (
            .O(N__14811),
            .I(\c0.n1197 ));
    LocalMux I__2822 (
            .O(N__14804),
            .I(\c0.n1197 ));
    LocalMux I__2821 (
            .O(N__14791),
            .I(\c0.n1197 ));
    Odrv12 I__2820 (
            .O(N__14786),
            .I(\c0.n1197 ));
    Odrv4 I__2819 (
            .O(N__14777),
            .I(\c0.n1197 ));
    Odrv4 I__2818 (
            .O(N__14772),
            .I(\c0.n1197 ));
    Odrv4 I__2817 (
            .O(N__14765),
            .I(\c0.n1197 ));
    Odrv12 I__2816 (
            .O(N__14762),
            .I(\c0.n1197 ));
    Odrv4 I__2815 (
            .O(N__14751),
            .I(\c0.n1197 ));
    CascadeMux I__2814 (
            .O(N__14726),
            .I(N__14717));
    CascadeMux I__2813 (
            .O(N__14725),
            .I(N__14708));
    CascadeMux I__2812 (
            .O(N__14724),
            .I(N__14699));
    CascadeMux I__2811 (
            .O(N__14723),
            .I(N__14696));
    CascadeMux I__2810 (
            .O(N__14722),
            .I(N__14690));
    CascadeMux I__2809 (
            .O(N__14721),
            .I(N__14681));
    InMux I__2808 (
            .O(N__14720),
            .I(N__14674));
    InMux I__2807 (
            .O(N__14717),
            .I(N__14674));
    InMux I__2806 (
            .O(N__14716),
            .I(N__14674));
    CascadeMux I__2805 (
            .O(N__14715),
            .I(N__14671));
    CascadeMux I__2804 (
            .O(N__14714),
            .I(N__14666));
    CascadeMux I__2803 (
            .O(N__14713),
            .I(N__14662));
    CascadeMux I__2802 (
            .O(N__14712),
            .I(N__14659));
    CascadeMux I__2801 (
            .O(N__14711),
            .I(N__14656));
    InMux I__2800 (
            .O(N__14708),
            .I(N__14647));
    InMux I__2799 (
            .O(N__14707),
            .I(N__14647));
    CascadeMux I__2798 (
            .O(N__14706),
            .I(N__14636));
    CascadeMux I__2797 (
            .O(N__14705),
            .I(N__14633));
    CascadeMux I__2796 (
            .O(N__14704),
            .I(N__14630));
    CascadeMux I__2795 (
            .O(N__14703),
            .I(N__14625));
    CascadeMux I__2794 (
            .O(N__14702),
            .I(N__14622));
    InMux I__2793 (
            .O(N__14699),
            .I(N__14612));
    InMux I__2792 (
            .O(N__14696),
            .I(N__14612));
    InMux I__2791 (
            .O(N__14695),
            .I(N__14612));
    InMux I__2790 (
            .O(N__14694),
            .I(N__14612));
    InMux I__2789 (
            .O(N__14693),
            .I(N__14607));
    InMux I__2788 (
            .O(N__14690),
            .I(N__14607));
    InMux I__2787 (
            .O(N__14689),
            .I(N__14598));
    InMux I__2786 (
            .O(N__14688),
            .I(N__14598));
    InMux I__2785 (
            .O(N__14687),
            .I(N__14598));
    InMux I__2784 (
            .O(N__14686),
            .I(N__14598));
    CascadeMux I__2783 (
            .O(N__14685),
            .I(N__14595));
    CascadeMux I__2782 (
            .O(N__14684),
            .I(N__14592));
    InMux I__2781 (
            .O(N__14681),
            .I(N__14586));
    LocalMux I__2780 (
            .O(N__14674),
            .I(N__14583));
    InMux I__2779 (
            .O(N__14671),
            .I(N__14580));
    CascadeMux I__2778 (
            .O(N__14670),
            .I(N__14575));
    CascadeMux I__2777 (
            .O(N__14669),
            .I(N__14571));
    InMux I__2776 (
            .O(N__14666),
            .I(N__14567));
    InMux I__2775 (
            .O(N__14665),
            .I(N__14562));
    InMux I__2774 (
            .O(N__14662),
            .I(N__14562));
    InMux I__2773 (
            .O(N__14659),
            .I(N__14555));
    InMux I__2772 (
            .O(N__14656),
            .I(N__14555));
    InMux I__2771 (
            .O(N__14655),
            .I(N__14555));
    InMux I__2770 (
            .O(N__14654),
            .I(N__14548));
    InMux I__2769 (
            .O(N__14653),
            .I(N__14548));
    InMux I__2768 (
            .O(N__14652),
            .I(N__14548));
    LocalMux I__2767 (
            .O(N__14647),
            .I(N__14545));
    InMux I__2766 (
            .O(N__14646),
            .I(N__14542));
    InMux I__2765 (
            .O(N__14645),
            .I(N__14531));
    InMux I__2764 (
            .O(N__14644),
            .I(N__14531));
    InMux I__2763 (
            .O(N__14643),
            .I(N__14531));
    InMux I__2762 (
            .O(N__14642),
            .I(N__14531));
    InMux I__2761 (
            .O(N__14641),
            .I(N__14531));
    InMux I__2760 (
            .O(N__14640),
            .I(N__14518));
    InMux I__2759 (
            .O(N__14639),
            .I(N__14518));
    InMux I__2758 (
            .O(N__14636),
            .I(N__14518));
    InMux I__2757 (
            .O(N__14633),
            .I(N__14518));
    InMux I__2756 (
            .O(N__14630),
            .I(N__14518));
    InMux I__2755 (
            .O(N__14629),
            .I(N__14518));
    InMux I__2754 (
            .O(N__14628),
            .I(N__14509));
    InMux I__2753 (
            .O(N__14625),
            .I(N__14509));
    InMux I__2752 (
            .O(N__14622),
            .I(N__14509));
    InMux I__2751 (
            .O(N__14621),
            .I(N__14509));
    LocalMux I__2750 (
            .O(N__14612),
            .I(N__14502));
    LocalMux I__2749 (
            .O(N__14607),
            .I(N__14502));
    LocalMux I__2748 (
            .O(N__14598),
            .I(N__14502));
    InMux I__2747 (
            .O(N__14595),
            .I(N__14496));
    InMux I__2746 (
            .O(N__14592),
            .I(N__14496));
    CascadeMux I__2745 (
            .O(N__14591),
            .I(N__14490));
    CascadeMux I__2744 (
            .O(N__14590),
            .I(N__14487));
    CascadeMux I__2743 (
            .O(N__14589),
            .I(N__14481));
    LocalMux I__2742 (
            .O(N__14586),
            .I(N__14474));
    Span4Mux_s3_v I__2741 (
            .O(N__14583),
            .I(N__14474));
    LocalMux I__2740 (
            .O(N__14580),
            .I(N__14474));
    CascadeMux I__2739 (
            .O(N__14579),
            .I(N__14469));
    CascadeMux I__2738 (
            .O(N__14578),
            .I(N__14466));
    InMux I__2737 (
            .O(N__14575),
            .I(N__14459));
    InMux I__2736 (
            .O(N__14574),
            .I(N__14459));
    InMux I__2735 (
            .O(N__14571),
            .I(N__14454));
    InMux I__2734 (
            .O(N__14570),
            .I(N__14454));
    LocalMux I__2733 (
            .O(N__14567),
            .I(N__14451));
    LocalMux I__2732 (
            .O(N__14562),
            .I(N__14432));
    LocalMux I__2731 (
            .O(N__14555),
            .I(N__14432));
    LocalMux I__2730 (
            .O(N__14548),
            .I(N__14432));
    Span4Mux_s2_h I__2729 (
            .O(N__14545),
            .I(N__14432));
    LocalMux I__2728 (
            .O(N__14542),
            .I(N__14432));
    LocalMux I__2727 (
            .O(N__14531),
            .I(N__14432));
    LocalMux I__2726 (
            .O(N__14518),
            .I(N__14432));
    LocalMux I__2725 (
            .O(N__14509),
            .I(N__14432));
    Span4Mux_s3_v I__2724 (
            .O(N__14502),
            .I(N__14432));
    CascadeMux I__2723 (
            .O(N__14501),
            .I(N__14429));
    LocalMux I__2722 (
            .O(N__14496),
            .I(N__14425));
    InMux I__2721 (
            .O(N__14495),
            .I(N__14420));
    InMux I__2720 (
            .O(N__14494),
            .I(N__14420));
    InMux I__2719 (
            .O(N__14493),
            .I(N__14407));
    InMux I__2718 (
            .O(N__14490),
            .I(N__14407));
    InMux I__2717 (
            .O(N__14487),
            .I(N__14407));
    InMux I__2716 (
            .O(N__14486),
            .I(N__14407));
    InMux I__2715 (
            .O(N__14485),
            .I(N__14407));
    InMux I__2714 (
            .O(N__14484),
            .I(N__14407));
    InMux I__2713 (
            .O(N__14481),
            .I(N__14401));
    Span4Mux_v I__2712 (
            .O(N__14474),
            .I(N__14398));
    InMux I__2711 (
            .O(N__14473),
            .I(N__14389));
    InMux I__2710 (
            .O(N__14472),
            .I(N__14389));
    InMux I__2709 (
            .O(N__14469),
            .I(N__14389));
    InMux I__2708 (
            .O(N__14466),
            .I(N__14389));
    InMux I__2707 (
            .O(N__14465),
            .I(N__14384));
    InMux I__2706 (
            .O(N__14464),
            .I(N__14384));
    LocalMux I__2705 (
            .O(N__14459),
            .I(N__14381));
    LocalMux I__2704 (
            .O(N__14454),
            .I(N__14376));
    Span4Mux_s3_h I__2703 (
            .O(N__14451),
            .I(N__14376));
    Span4Mux_v I__2702 (
            .O(N__14432),
            .I(N__14373));
    InMux I__2701 (
            .O(N__14429),
            .I(N__14370));
    InMux I__2700 (
            .O(N__14428),
            .I(N__14367));
    Span4Mux_v I__2699 (
            .O(N__14425),
            .I(N__14362));
    LocalMux I__2698 (
            .O(N__14420),
            .I(N__14362));
    LocalMux I__2697 (
            .O(N__14407),
            .I(N__14359));
    InMux I__2696 (
            .O(N__14406),
            .I(N__14354));
    InMux I__2695 (
            .O(N__14405),
            .I(N__14354));
    InMux I__2694 (
            .O(N__14404),
            .I(N__14351));
    LocalMux I__2693 (
            .O(N__14401),
            .I(N__14346));
    Span4Mux_s0_h I__2692 (
            .O(N__14398),
            .I(N__14346));
    LocalMux I__2691 (
            .O(N__14389),
            .I(N__14337));
    LocalMux I__2690 (
            .O(N__14384),
            .I(N__14337));
    Span4Mux_s3_h I__2689 (
            .O(N__14381),
            .I(N__14337));
    Span4Mux_v I__2688 (
            .O(N__14376),
            .I(N__14337));
    Span4Mux_s2_h I__2687 (
            .O(N__14373),
            .I(N__14334));
    LocalMux I__2686 (
            .O(N__14370),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    LocalMux I__2685 (
            .O(N__14367),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__2684 (
            .O(N__14362),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv12 I__2683 (
            .O(N__14359),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    LocalMux I__2682 (
            .O(N__14354),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    LocalMux I__2681 (
            .O(N__14351),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__2680 (
            .O(N__14346),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__2679 (
            .O(N__14337),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__2678 (
            .O(N__14334),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    InMux I__2677 (
            .O(N__14315),
            .I(N__14312));
    LocalMux I__2676 (
            .O(N__14312),
            .I(N__14307));
    CascadeMux I__2675 (
            .O(N__14311),
            .I(N__14304));
    InMux I__2674 (
            .O(N__14310),
            .I(N__14301));
    Span4Mux_v I__2673 (
            .O(N__14307),
            .I(N__14298));
    InMux I__2672 (
            .O(N__14304),
            .I(N__14295));
    LocalMux I__2671 (
            .O(N__14301),
            .I(\c0.data_in_field_10 ));
    Odrv4 I__2670 (
            .O(N__14298),
            .I(\c0.data_in_field_10 ));
    LocalMux I__2669 (
            .O(N__14295),
            .I(\c0.data_in_field_10 ));
    InMux I__2668 (
            .O(N__14288),
            .I(N__14284));
    InMux I__2667 (
            .O(N__14287),
            .I(N__14281));
    LocalMux I__2666 (
            .O(N__14284),
            .I(n2651));
    LocalMux I__2665 (
            .O(N__14281),
            .I(n2651));
    CascadeMux I__2664 (
            .O(N__14276),
            .I(N__14273));
    InMux I__2663 (
            .O(N__14273),
            .I(N__14268));
    InMux I__2662 (
            .O(N__14272),
            .I(N__14265));
    InMux I__2661 (
            .O(N__14271),
            .I(N__14262));
    LocalMux I__2660 (
            .O(N__14268),
            .I(data_in_5_0));
    LocalMux I__2659 (
            .O(N__14265),
            .I(data_in_5_0));
    LocalMux I__2658 (
            .O(N__14262),
            .I(data_in_5_0));
    InMux I__2657 (
            .O(N__14255),
            .I(N__14251));
    InMux I__2656 (
            .O(N__14254),
            .I(N__14248));
    LocalMux I__2655 (
            .O(N__14251),
            .I(N__14242));
    LocalMux I__2654 (
            .O(N__14248),
            .I(N__14242));
    InMux I__2653 (
            .O(N__14247),
            .I(N__14239));
    Odrv4 I__2652 (
            .O(N__14242),
            .I(data_in_4_0));
    LocalMux I__2651 (
            .O(N__14239),
            .I(data_in_4_0));
    InMux I__2650 (
            .O(N__14234),
            .I(N__14231));
    LocalMux I__2649 (
            .O(N__14231),
            .I(N__14228));
    Span4Mux_h I__2648 (
            .O(N__14228),
            .I(N__14223));
    InMux I__2647 (
            .O(N__14227),
            .I(N__14220));
    InMux I__2646 (
            .O(N__14226),
            .I(N__14217));
    Odrv4 I__2645 (
            .O(N__14223),
            .I(data_in_4_3));
    LocalMux I__2644 (
            .O(N__14220),
            .I(data_in_4_3));
    LocalMux I__2643 (
            .O(N__14217),
            .I(data_in_4_3));
    InMux I__2642 (
            .O(N__14210),
            .I(N__14206));
    InMux I__2641 (
            .O(N__14209),
            .I(N__14203));
    LocalMux I__2640 (
            .O(N__14206),
            .I(N__14198));
    LocalMux I__2639 (
            .O(N__14203),
            .I(N__14195));
    InMux I__2638 (
            .O(N__14202),
            .I(N__14192));
    InMux I__2637 (
            .O(N__14201),
            .I(N__14189));
    Span4Mux_v I__2636 (
            .O(N__14198),
            .I(N__14182));
    Span4Mux_s2_v I__2635 (
            .O(N__14195),
            .I(N__14182));
    LocalMux I__2634 (
            .O(N__14192),
            .I(N__14182));
    LocalMux I__2633 (
            .O(N__14189),
            .I(data_in_3_3));
    Odrv4 I__2632 (
            .O(N__14182),
            .I(data_in_3_3));
    CascadeMux I__2631 (
            .O(N__14177),
            .I(N__14174));
    InMux I__2630 (
            .O(N__14174),
            .I(N__14170));
    InMux I__2629 (
            .O(N__14173),
            .I(N__14167));
    LocalMux I__2628 (
            .O(N__14170),
            .I(N__14162));
    LocalMux I__2627 (
            .O(N__14167),
            .I(N__14162));
    Span4Mux_v I__2626 (
            .O(N__14162),
            .I(N__14158));
    InMux I__2625 (
            .O(N__14161),
            .I(N__14155));
    Odrv4 I__2624 (
            .O(N__14158),
            .I(data_in_5_2));
    LocalMux I__2623 (
            .O(N__14155),
            .I(data_in_5_2));
    InMux I__2622 (
            .O(N__14150),
            .I(N__14146));
    CascadeMux I__2621 (
            .O(N__14149),
            .I(N__14143));
    LocalMux I__2620 (
            .O(N__14146),
            .I(N__14139));
    InMux I__2619 (
            .O(N__14143),
            .I(N__14134));
    InMux I__2618 (
            .O(N__14142),
            .I(N__14134));
    Odrv12 I__2617 (
            .O(N__14139),
            .I(n1222));
    LocalMux I__2616 (
            .O(N__14134),
            .I(n1222));
    CascadeMux I__2615 (
            .O(N__14129),
            .I(N__14125));
    InMux I__2614 (
            .O(N__14128),
            .I(N__14122));
    InMux I__2613 (
            .O(N__14125),
            .I(N__14119));
    LocalMux I__2612 (
            .O(N__14122),
            .I(N__14115));
    LocalMux I__2611 (
            .O(N__14119),
            .I(N__14111));
    InMux I__2610 (
            .O(N__14118),
            .I(N__14108));
    Span4Mux_h I__2609 (
            .O(N__14115),
            .I(N__14105));
    InMux I__2608 (
            .O(N__14114),
            .I(N__14102));
    Span4Mux_h I__2607 (
            .O(N__14111),
            .I(N__14099));
    LocalMux I__2606 (
            .O(N__14108),
            .I(data_in_7_3));
    Odrv4 I__2605 (
            .O(N__14105),
            .I(data_in_7_3));
    LocalMux I__2604 (
            .O(N__14102),
            .I(data_in_7_3));
    Odrv4 I__2603 (
            .O(N__14099),
            .I(data_in_7_3));
    InMux I__2602 (
            .O(N__14090),
            .I(N__14087));
    LocalMux I__2601 (
            .O(N__14087),
            .I(N__14081));
    InMux I__2600 (
            .O(N__14086),
            .I(N__14078));
    InMux I__2599 (
            .O(N__14085),
            .I(N__14073));
    InMux I__2598 (
            .O(N__14084),
            .I(N__14073));
    Span4Mux_v I__2597 (
            .O(N__14081),
            .I(N__14070));
    LocalMux I__2596 (
            .O(N__14078),
            .I(N__14067));
    LocalMux I__2595 (
            .O(N__14073),
            .I(data_in_7_6));
    Odrv4 I__2594 (
            .O(N__14070),
            .I(data_in_7_6));
    Odrv4 I__2593 (
            .O(N__14067),
            .I(data_in_7_6));
    IoInMux I__2592 (
            .O(N__14060),
            .I(N__14057));
    LocalMux I__2591 (
            .O(N__14057),
            .I(N__14053));
    InMux I__2590 (
            .O(N__14056),
            .I(N__14050));
    Span4Mux_s3_h I__2589 (
            .O(N__14053),
            .I(N__14046));
    LocalMux I__2588 (
            .O(N__14050),
            .I(N__14043));
    InMux I__2587 (
            .O(N__14049),
            .I(N__14040));
    Odrv4 I__2586 (
            .O(N__14046),
            .I(tx2_o_adj_949));
    Odrv4 I__2585 (
            .O(N__14043),
            .I(tx2_o_adj_949));
    LocalMux I__2584 (
            .O(N__14040),
            .I(tx2_o_adj_949));
    IoInMux I__2583 (
            .O(N__14033),
            .I(N__14030));
    LocalMux I__2582 (
            .O(N__14030),
            .I(N__14027));
    Span4Mux_s0_h I__2581 (
            .O(N__14027),
            .I(N__14024));
    Span4Mux_h I__2580 (
            .O(N__14024),
            .I(N__14021));
    Odrv4 I__2579 (
            .O(N__14021),
            .I(tx2_enable));
    InMux I__2578 (
            .O(N__14018),
            .I(N__14015));
    LocalMux I__2577 (
            .O(N__14015),
            .I(N__14009));
    CascadeMux I__2576 (
            .O(N__14014),
            .I(N__14006));
    InMux I__2575 (
            .O(N__14013),
            .I(N__14002));
    InMux I__2574 (
            .O(N__14012),
            .I(N__13999));
    Span12Mux_h I__2573 (
            .O(N__14009),
            .I(N__13996));
    InMux I__2572 (
            .O(N__14006),
            .I(N__13993));
    InMux I__2571 (
            .O(N__14005),
            .I(N__13990));
    LocalMux I__2570 (
            .O(N__14002),
            .I(N__13987));
    LocalMux I__2569 (
            .O(N__13999),
            .I(\c0.data_in_field_12 ));
    Odrv12 I__2568 (
            .O(N__13996),
            .I(\c0.data_in_field_12 ));
    LocalMux I__2567 (
            .O(N__13993),
            .I(\c0.data_in_field_12 ));
    LocalMux I__2566 (
            .O(N__13990),
            .I(\c0.data_in_field_12 ));
    Odrv12 I__2565 (
            .O(N__13987),
            .I(\c0.data_in_field_12 ));
    InMux I__2564 (
            .O(N__13976),
            .I(N__13973));
    LocalMux I__2563 (
            .O(N__13973),
            .I(N__13968));
    InMux I__2562 (
            .O(N__13972),
            .I(N__13965));
    InMux I__2561 (
            .O(N__13971),
            .I(N__13960));
    Sp12to4 I__2560 (
            .O(N__13968),
            .I(N__13955));
    LocalMux I__2559 (
            .O(N__13965),
            .I(N__13955));
    InMux I__2558 (
            .O(N__13964),
            .I(N__13952));
    InMux I__2557 (
            .O(N__13963),
            .I(N__13949));
    LocalMux I__2556 (
            .O(N__13960),
            .I(\c0.data_in_field_40 ));
    Odrv12 I__2555 (
            .O(N__13955),
            .I(\c0.data_in_field_40 ));
    LocalMux I__2554 (
            .O(N__13952),
            .I(\c0.data_in_field_40 ));
    LocalMux I__2553 (
            .O(N__13949),
            .I(\c0.data_in_field_40 ));
    InMux I__2552 (
            .O(N__13940),
            .I(N__13936));
    InMux I__2551 (
            .O(N__13939),
            .I(N__13932));
    LocalMux I__2550 (
            .O(N__13936),
            .I(N__13929));
    CascadeMux I__2549 (
            .O(N__13935),
            .I(N__13925));
    LocalMux I__2548 (
            .O(N__13932),
            .I(N__13922));
    Span4Mux_h I__2547 (
            .O(N__13929),
            .I(N__13919));
    InMux I__2546 (
            .O(N__13928),
            .I(N__13914));
    InMux I__2545 (
            .O(N__13925),
            .I(N__13914));
    Odrv12 I__2544 (
            .O(N__13922),
            .I(data_in_6_6));
    Odrv4 I__2543 (
            .O(N__13919),
            .I(data_in_6_6));
    LocalMux I__2542 (
            .O(N__13914),
            .I(data_in_6_6));
    CascadeMux I__2541 (
            .O(N__13907),
            .I(N__13903));
    InMux I__2540 (
            .O(N__13906),
            .I(N__13900));
    InMux I__2539 (
            .O(N__13903),
            .I(N__13897));
    LocalMux I__2538 (
            .O(N__13900),
            .I(N__13890));
    LocalMux I__2537 (
            .O(N__13897),
            .I(N__13890));
    InMux I__2536 (
            .O(N__13896),
            .I(N__13887));
    InMux I__2535 (
            .O(N__13895),
            .I(N__13883));
    Span4Mux_h I__2534 (
            .O(N__13890),
            .I(N__13880));
    LocalMux I__2533 (
            .O(N__13887),
            .I(N__13877));
    InMux I__2532 (
            .O(N__13886),
            .I(N__13874));
    LocalMux I__2531 (
            .O(N__13883),
            .I(\c0.data_in_field_41 ));
    Odrv4 I__2530 (
            .O(N__13880),
            .I(\c0.data_in_field_41 ));
    Odrv12 I__2529 (
            .O(N__13877),
            .I(\c0.data_in_field_41 ));
    LocalMux I__2528 (
            .O(N__13874),
            .I(\c0.data_in_field_41 ));
    InMux I__2527 (
            .O(N__13865),
            .I(N__13862));
    LocalMux I__2526 (
            .O(N__13862),
            .I(N__13859));
    Odrv4 I__2525 (
            .O(N__13859),
            .I(\c0.n12_adj_878 ));
    InMux I__2524 (
            .O(N__13856),
            .I(N__13853));
    LocalMux I__2523 (
            .O(N__13853),
            .I(N__13849));
    CascadeMux I__2522 (
            .O(N__13852),
            .I(N__13846));
    Span4Mux_h I__2521 (
            .O(N__13849),
            .I(N__13843));
    InMux I__2520 (
            .O(N__13846),
            .I(N__13840));
    Odrv4 I__2519 (
            .O(N__13843),
            .I(rx_data_4));
    LocalMux I__2518 (
            .O(N__13840),
            .I(rx_data_4));
    InMux I__2517 (
            .O(N__13835),
            .I(N__13832));
    LocalMux I__2516 (
            .O(N__13832),
            .I(N__13828));
    CascadeMux I__2515 (
            .O(N__13831),
            .I(N__13825));
    Span4Mux_h I__2514 (
            .O(N__13828),
            .I(N__13822));
    InMux I__2513 (
            .O(N__13825),
            .I(N__13817));
    Span4Mux_v I__2512 (
            .O(N__13822),
            .I(N__13814));
    InMux I__2511 (
            .O(N__13821),
            .I(N__13811));
    InMux I__2510 (
            .O(N__13820),
            .I(N__13808));
    LocalMux I__2509 (
            .O(N__13817),
            .I(N__13805));
    Odrv4 I__2508 (
            .O(N__13814),
            .I(data_in_7_4));
    LocalMux I__2507 (
            .O(N__13811),
            .I(data_in_7_4));
    LocalMux I__2506 (
            .O(N__13808),
            .I(data_in_7_4));
    Odrv4 I__2505 (
            .O(N__13805),
            .I(data_in_7_4));
    InMux I__2504 (
            .O(N__13796),
            .I(N__13793));
    LocalMux I__2503 (
            .O(N__13793),
            .I(N__13789));
    InMux I__2502 (
            .O(N__13792),
            .I(N__13786));
    Span4Mux_h I__2501 (
            .O(N__13789),
            .I(N__13781));
    LocalMux I__2500 (
            .O(N__13786),
            .I(N__13778));
    InMux I__2499 (
            .O(N__13785),
            .I(N__13775));
    InMux I__2498 (
            .O(N__13784),
            .I(N__13772));
    Odrv4 I__2497 (
            .O(N__13781),
            .I(data_in_3_0));
    Odrv4 I__2496 (
            .O(N__13778),
            .I(data_in_3_0));
    LocalMux I__2495 (
            .O(N__13775),
            .I(data_in_3_0));
    LocalMux I__2494 (
            .O(N__13772),
            .I(data_in_3_0));
    InMux I__2493 (
            .O(N__13763),
            .I(N__13760));
    LocalMux I__2492 (
            .O(N__13760),
            .I(N__13756));
    InMux I__2491 (
            .O(N__13759),
            .I(N__13753));
    Span4Mux_v I__2490 (
            .O(N__13756),
            .I(N__13746));
    LocalMux I__2489 (
            .O(N__13753),
            .I(N__13746));
    InMux I__2488 (
            .O(N__13752),
            .I(N__13743));
    InMux I__2487 (
            .O(N__13751),
            .I(N__13739));
    Span4Mux_h I__2486 (
            .O(N__13746),
            .I(N__13734));
    LocalMux I__2485 (
            .O(N__13743),
            .I(N__13734));
    InMux I__2484 (
            .O(N__13742),
            .I(N__13731));
    LocalMux I__2483 (
            .O(N__13739),
            .I(\c0.data_in_field_24 ));
    Odrv4 I__2482 (
            .O(N__13734),
            .I(\c0.data_in_field_24 ));
    LocalMux I__2481 (
            .O(N__13731),
            .I(\c0.data_in_field_24 ));
    InMux I__2480 (
            .O(N__13724),
            .I(N__13719));
    InMux I__2479 (
            .O(N__13723),
            .I(N__13716));
    CascadeMux I__2478 (
            .O(N__13722),
            .I(N__13713));
    LocalMux I__2477 (
            .O(N__13719),
            .I(N__13709));
    LocalMux I__2476 (
            .O(N__13716),
            .I(N__13706));
    InMux I__2475 (
            .O(N__13713),
            .I(N__13703));
    InMux I__2474 (
            .O(N__13712),
            .I(N__13700));
    Span4Mux_v I__2473 (
            .O(N__13709),
            .I(N__13697));
    Span4Mux_v I__2472 (
            .O(N__13706),
            .I(N__13692));
    LocalMux I__2471 (
            .O(N__13703),
            .I(N__13692));
    LocalMux I__2470 (
            .O(N__13700),
            .I(data_in_7_7));
    Odrv4 I__2469 (
            .O(N__13697),
            .I(data_in_7_7));
    Odrv4 I__2468 (
            .O(N__13692),
            .I(data_in_7_7));
    InMux I__2467 (
            .O(N__13685),
            .I(N__13682));
    LocalMux I__2466 (
            .O(N__13682),
            .I(N__13678));
    InMux I__2465 (
            .O(N__13681),
            .I(N__13675));
    Span4Mux_h I__2464 (
            .O(N__13678),
            .I(N__13670));
    LocalMux I__2463 (
            .O(N__13675),
            .I(N__13667));
    InMux I__2462 (
            .O(N__13674),
            .I(N__13664));
    InMux I__2461 (
            .O(N__13673),
            .I(N__13661));
    Odrv4 I__2460 (
            .O(N__13670),
            .I(data_in_6_7));
    Odrv4 I__2459 (
            .O(N__13667),
            .I(data_in_6_7));
    LocalMux I__2458 (
            .O(N__13664),
            .I(data_in_6_7));
    LocalMux I__2457 (
            .O(N__13661),
            .I(data_in_6_7));
    CascadeMux I__2456 (
            .O(N__13652),
            .I(N__13649));
    InMux I__2455 (
            .O(N__13649),
            .I(N__13646));
    LocalMux I__2454 (
            .O(N__13646),
            .I(N__13640));
    InMux I__2453 (
            .O(N__13645),
            .I(N__13637));
    InMux I__2452 (
            .O(N__13644),
            .I(N__13631));
    InMux I__2451 (
            .O(N__13643),
            .I(N__13631));
    Span4Mux_h I__2450 (
            .O(N__13640),
            .I(N__13628));
    LocalMux I__2449 (
            .O(N__13637),
            .I(N__13625));
    InMux I__2448 (
            .O(N__13636),
            .I(N__13622));
    LocalMux I__2447 (
            .O(N__13631),
            .I(\c0.data_in_field_35 ));
    Odrv4 I__2446 (
            .O(N__13628),
            .I(\c0.data_in_field_35 ));
    Odrv4 I__2445 (
            .O(N__13625),
            .I(\c0.data_in_field_35 ));
    LocalMux I__2444 (
            .O(N__13622),
            .I(\c0.data_in_field_35 ));
    InMux I__2443 (
            .O(N__13613),
            .I(N__13609));
    CascadeMux I__2442 (
            .O(N__13612),
            .I(N__13605));
    LocalMux I__2441 (
            .O(N__13609),
            .I(N__13602));
    InMux I__2440 (
            .O(N__13608),
            .I(N__13599));
    InMux I__2439 (
            .O(N__13605),
            .I(N__13594));
    Span4Mux_v I__2438 (
            .O(N__13602),
            .I(N__13591));
    LocalMux I__2437 (
            .O(N__13599),
            .I(N__13588));
    InMux I__2436 (
            .O(N__13598),
            .I(N__13585));
    InMux I__2435 (
            .O(N__13597),
            .I(N__13582));
    LocalMux I__2434 (
            .O(N__13594),
            .I(\c0.data_in_field_36 ));
    Odrv4 I__2433 (
            .O(N__13591),
            .I(\c0.data_in_field_36 ));
    Odrv4 I__2432 (
            .O(N__13588),
            .I(\c0.data_in_field_36 ));
    LocalMux I__2431 (
            .O(N__13585),
            .I(\c0.data_in_field_36 ));
    LocalMux I__2430 (
            .O(N__13582),
            .I(\c0.data_in_field_36 ));
    InMux I__2429 (
            .O(N__13571),
            .I(N__13568));
    LocalMux I__2428 (
            .O(N__13568),
            .I(\c0.n11 ));
    CascadeMux I__2427 (
            .O(N__13565),
            .I(N__13562));
    InMux I__2426 (
            .O(N__13562),
            .I(N__13559));
    LocalMux I__2425 (
            .O(N__13559),
            .I(N__13555));
    InMux I__2424 (
            .O(N__13558),
            .I(N__13550));
    Span4Mux_h I__2423 (
            .O(N__13555),
            .I(N__13547));
    InMux I__2422 (
            .O(N__13554),
            .I(N__13542));
    InMux I__2421 (
            .O(N__13553),
            .I(N__13542));
    LocalMux I__2420 (
            .O(N__13550),
            .I(\c0.data_in_field_43 ));
    Odrv4 I__2419 (
            .O(N__13547),
            .I(\c0.data_in_field_43 ));
    LocalMux I__2418 (
            .O(N__13542),
            .I(\c0.data_in_field_43 ));
    InMux I__2417 (
            .O(N__13535),
            .I(N__13532));
    LocalMux I__2416 (
            .O(N__13532),
            .I(N__13527));
    InMux I__2415 (
            .O(N__13531),
            .I(N__13522));
    InMux I__2414 (
            .O(N__13530),
            .I(N__13519));
    Span4Mux_h I__2413 (
            .O(N__13527),
            .I(N__13516));
    InMux I__2412 (
            .O(N__13526),
            .I(N__13513));
    InMux I__2411 (
            .O(N__13525),
            .I(N__13510));
    LocalMux I__2410 (
            .O(N__13522),
            .I(\c0.data_in_field_26 ));
    LocalMux I__2409 (
            .O(N__13519),
            .I(\c0.data_in_field_26 ));
    Odrv4 I__2408 (
            .O(N__13516),
            .I(\c0.data_in_field_26 ));
    LocalMux I__2407 (
            .O(N__13513),
            .I(\c0.data_in_field_26 ));
    LocalMux I__2406 (
            .O(N__13510),
            .I(\c0.data_in_field_26 ));
    CascadeMux I__2405 (
            .O(N__13499),
            .I(\c0.n4415_cascade_ ));
    InMux I__2404 (
            .O(N__13496),
            .I(N__13492));
    InMux I__2403 (
            .O(N__13495),
            .I(N__13489));
    LocalMux I__2402 (
            .O(N__13492),
            .I(N__13486));
    LocalMux I__2401 (
            .O(N__13489),
            .I(N__13482));
    Span4Mux_v I__2400 (
            .O(N__13486),
            .I(N__13477));
    InMux I__2399 (
            .O(N__13485),
            .I(N__13474));
    Span4Mux_s3_h I__2398 (
            .O(N__13482),
            .I(N__13471));
    InMux I__2397 (
            .O(N__13481),
            .I(N__13466));
    InMux I__2396 (
            .O(N__13480),
            .I(N__13466));
    Odrv4 I__2395 (
            .O(N__13477),
            .I(\c0.data_in_field_9 ));
    LocalMux I__2394 (
            .O(N__13474),
            .I(\c0.data_in_field_9 ));
    Odrv4 I__2393 (
            .O(N__13471),
            .I(\c0.data_in_field_9 ));
    LocalMux I__2392 (
            .O(N__13466),
            .I(\c0.data_in_field_9 ));
    InMux I__2391 (
            .O(N__13457),
            .I(N__13454));
    LocalMux I__2390 (
            .O(N__13454),
            .I(N__13451));
    Odrv4 I__2389 (
            .O(N__13451),
            .I(\c0.n23 ));
    InMux I__2388 (
            .O(N__13448),
            .I(N__13444));
    CascadeMux I__2387 (
            .O(N__13447),
            .I(N__13440));
    LocalMux I__2386 (
            .O(N__13444),
            .I(N__13437));
    InMux I__2385 (
            .O(N__13443),
            .I(N__13434));
    InMux I__2384 (
            .O(N__13440),
            .I(N__13429));
    Span4Mux_v I__2383 (
            .O(N__13437),
            .I(N__13426));
    LocalMux I__2382 (
            .O(N__13434),
            .I(N__13423));
    InMux I__2381 (
            .O(N__13433),
            .I(N__13420));
    InMux I__2380 (
            .O(N__13432),
            .I(N__13417));
    LocalMux I__2379 (
            .O(N__13429),
            .I(\c0.data_in_field_30 ));
    Odrv4 I__2378 (
            .O(N__13426),
            .I(\c0.data_in_field_30 ));
    Odrv4 I__2377 (
            .O(N__13423),
            .I(\c0.data_in_field_30 ));
    LocalMux I__2376 (
            .O(N__13420),
            .I(\c0.data_in_field_30 ));
    LocalMux I__2375 (
            .O(N__13417),
            .I(\c0.data_in_field_30 ));
    InMux I__2374 (
            .O(N__13406),
            .I(N__13403));
    LocalMux I__2373 (
            .O(N__13403),
            .I(N__13400));
    Span4Mux_h I__2372 (
            .O(N__13400),
            .I(N__13397));
    Odrv4 I__2371 (
            .O(N__13397),
            .I(\c0.n4927 ));
    InMux I__2370 (
            .O(N__13394),
            .I(N__13390));
    InMux I__2369 (
            .O(N__13393),
            .I(N__13387));
    LocalMux I__2368 (
            .O(N__13390),
            .I(\c0.n1267 ));
    LocalMux I__2367 (
            .O(N__13387),
            .I(\c0.n1267 ));
    InMux I__2366 (
            .O(N__13382),
            .I(N__13379));
    LocalMux I__2365 (
            .O(N__13379),
            .I(\c0.n4421 ));
    InMux I__2364 (
            .O(N__13376),
            .I(N__13373));
    LocalMux I__2363 (
            .O(N__13373),
            .I(N__13370));
    Span4Mux_s3_h I__2362 (
            .O(N__13370),
            .I(N__13363));
    InMux I__2361 (
            .O(N__13369),
            .I(N__13360));
    InMux I__2360 (
            .O(N__13368),
            .I(N__13357));
    InMux I__2359 (
            .O(N__13367),
            .I(N__13352));
    InMux I__2358 (
            .O(N__13366),
            .I(N__13352));
    Odrv4 I__2357 (
            .O(N__13363),
            .I(\c0.data_in_field_23 ));
    LocalMux I__2356 (
            .O(N__13360),
            .I(\c0.data_in_field_23 ));
    LocalMux I__2355 (
            .O(N__13357),
            .I(\c0.data_in_field_23 ));
    LocalMux I__2354 (
            .O(N__13352),
            .I(\c0.data_in_field_23 ));
    InMux I__2353 (
            .O(N__13343),
            .I(N__13338));
    CascadeMux I__2352 (
            .O(N__13342),
            .I(N__13335));
    InMux I__2351 (
            .O(N__13341),
            .I(N__13332));
    LocalMux I__2350 (
            .O(N__13338),
            .I(N__13329));
    InMux I__2349 (
            .O(N__13335),
            .I(N__13324));
    LocalMux I__2348 (
            .O(N__13332),
            .I(N__13321));
    Span4Mux_h I__2347 (
            .O(N__13329),
            .I(N__13318));
    InMux I__2346 (
            .O(N__13328),
            .I(N__13313));
    InMux I__2345 (
            .O(N__13327),
            .I(N__13313));
    LocalMux I__2344 (
            .O(N__13324),
            .I(\c0.data_in_field_37 ));
    Odrv12 I__2343 (
            .O(N__13321),
            .I(\c0.data_in_field_37 ));
    Odrv4 I__2342 (
            .O(N__13318),
            .I(\c0.data_in_field_37 ));
    LocalMux I__2341 (
            .O(N__13313),
            .I(\c0.data_in_field_37 ));
    InMux I__2340 (
            .O(N__13304),
            .I(N__13301));
    LocalMux I__2339 (
            .O(N__13301),
            .I(\c0.n8_adj_883 ));
    CascadeMux I__2338 (
            .O(N__13298),
            .I(N__13294));
    InMux I__2337 (
            .O(N__13297),
            .I(N__13290));
    InMux I__2336 (
            .O(N__13294),
            .I(N__13285));
    InMux I__2335 (
            .O(N__13293),
            .I(N__13285));
    LocalMux I__2334 (
            .O(N__13290),
            .I(N__13280));
    LocalMux I__2333 (
            .O(N__13285),
            .I(N__13277));
    InMux I__2332 (
            .O(N__13284),
            .I(N__13272));
    InMux I__2331 (
            .O(N__13283),
            .I(N__13272));
    Odrv4 I__2330 (
            .O(N__13280),
            .I(\c0.data_in_field_25 ));
    Odrv4 I__2329 (
            .O(N__13277),
            .I(\c0.data_in_field_25 ));
    LocalMux I__2328 (
            .O(N__13272),
            .I(\c0.data_in_field_25 ));
    CascadeMux I__2327 (
            .O(N__13265),
            .I(N__13260));
    InMux I__2326 (
            .O(N__13264),
            .I(N__13257));
    InMux I__2325 (
            .O(N__13263),
            .I(N__13254));
    InMux I__2324 (
            .O(N__13260),
            .I(N__13251));
    LocalMux I__2323 (
            .O(N__13257),
            .I(N__13242));
    LocalMux I__2322 (
            .O(N__13254),
            .I(N__13242));
    LocalMux I__2321 (
            .O(N__13251),
            .I(N__13242));
    InMux I__2320 (
            .O(N__13250),
            .I(N__13237));
    InMux I__2319 (
            .O(N__13249),
            .I(N__13237));
    Odrv4 I__2318 (
            .O(N__13242),
            .I(\c0.n1290 ));
    LocalMux I__2317 (
            .O(N__13237),
            .I(\c0.n1290 ));
    InMux I__2316 (
            .O(N__13232),
            .I(N__13229));
    LocalMux I__2315 (
            .O(N__13229),
            .I(N__13226));
    Odrv4 I__2314 (
            .O(N__13226),
            .I(\c0.n4441 ));
    InMux I__2313 (
            .O(N__13223),
            .I(N__13218));
    InMux I__2312 (
            .O(N__13222),
            .I(N__13215));
    InMux I__2311 (
            .O(N__13221),
            .I(N__13211));
    LocalMux I__2310 (
            .O(N__13218),
            .I(N__13208));
    LocalMux I__2309 (
            .O(N__13215),
            .I(N__13205));
    InMux I__2308 (
            .O(N__13214),
            .I(N__13202));
    LocalMux I__2307 (
            .O(N__13211),
            .I(\c0.data_in_field_28 ));
    Odrv4 I__2306 (
            .O(N__13208),
            .I(\c0.data_in_field_28 ));
    Odrv4 I__2305 (
            .O(N__13205),
            .I(\c0.data_in_field_28 ));
    LocalMux I__2304 (
            .O(N__13202),
            .I(\c0.data_in_field_28 ));
    InMux I__2303 (
            .O(N__13193),
            .I(N__13190));
    LocalMux I__2302 (
            .O(N__13190),
            .I(N__13186));
    InMux I__2301 (
            .O(N__13189),
            .I(N__13179));
    Span4Mux_v I__2300 (
            .O(N__13186),
            .I(N__13176));
    InMux I__2299 (
            .O(N__13185),
            .I(N__13173));
    InMux I__2298 (
            .O(N__13184),
            .I(N__13170));
    InMux I__2297 (
            .O(N__13183),
            .I(N__13167));
    InMux I__2296 (
            .O(N__13182),
            .I(N__13164));
    LocalMux I__2295 (
            .O(N__13179),
            .I(\c0.data_in_field_42 ));
    Odrv4 I__2294 (
            .O(N__13176),
            .I(\c0.data_in_field_42 ));
    LocalMux I__2293 (
            .O(N__13173),
            .I(\c0.data_in_field_42 ));
    LocalMux I__2292 (
            .O(N__13170),
            .I(\c0.data_in_field_42 ));
    LocalMux I__2291 (
            .O(N__13167),
            .I(\c0.data_in_field_42 ));
    LocalMux I__2290 (
            .O(N__13164),
            .I(\c0.data_in_field_42 ));
    InMux I__2289 (
            .O(N__13151),
            .I(N__13148));
    LocalMux I__2288 (
            .O(N__13148),
            .I(N__13142));
    InMux I__2287 (
            .O(N__13147),
            .I(N__13139));
    InMux I__2286 (
            .O(N__13146),
            .I(N__13134));
    InMux I__2285 (
            .O(N__13145),
            .I(N__13134));
    Span4Mux_h I__2284 (
            .O(N__13142),
            .I(N__13131));
    LocalMux I__2283 (
            .O(N__13139),
            .I(N__13128));
    LocalMux I__2282 (
            .O(N__13134),
            .I(\c0.data_in_field_13 ));
    Odrv4 I__2281 (
            .O(N__13131),
            .I(\c0.data_in_field_13 ));
    Odrv12 I__2280 (
            .O(N__13128),
            .I(\c0.data_in_field_13 ));
    InMux I__2279 (
            .O(N__13121),
            .I(N__13117));
    InMux I__2278 (
            .O(N__13120),
            .I(N__13114));
    LocalMux I__2277 (
            .O(N__13117),
            .I(\c0.n4414 ));
    LocalMux I__2276 (
            .O(N__13114),
            .I(\c0.n4414 ));
    CascadeMux I__2275 (
            .O(N__13109),
            .I(\c0.n30_adj_892_cascade_ ));
    InMux I__2274 (
            .O(N__13106),
            .I(N__13103));
    LocalMux I__2273 (
            .O(N__13103),
            .I(\c0.n25_adj_893 ));
    CascadeMux I__2272 (
            .O(N__13100),
            .I(N__13095));
    CascadeMux I__2271 (
            .O(N__13099),
            .I(N__13092));
    InMux I__2270 (
            .O(N__13098),
            .I(N__13086));
    InMux I__2269 (
            .O(N__13095),
            .I(N__13086));
    InMux I__2268 (
            .O(N__13092),
            .I(N__13081));
    InMux I__2267 (
            .O(N__13091),
            .I(N__13081));
    LocalMux I__2266 (
            .O(N__13086),
            .I(\c0.n2637 ));
    LocalMux I__2265 (
            .O(N__13081),
            .I(\c0.n2637 ));
    InMux I__2264 (
            .O(N__13076),
            .I(N__13072));
    InMux I__2263 (
            .O(N__13075),
            .I(N__13069));
    LocalMux I__2262 (
            .O(N__13072),
            .I(N__13065));
    LocalMux I__2261 (
            .O(N__13069),
            .I(N__13062));
    InMux I__2260 (
            .O(N__13068),
            .I(N__13059));
    Span4Mux_h I__2259 (
            .O(N__13065),
            .I(N__13056));
    Span4Mux_h I__2258 (
            .O(N__13062),
            .I(N__13053));
    LocalMux I__2257 (
            .O(N__13059),
            .I(\c0.n1261 ));
    Odrv4 I__2256 (
            .O(N__13056),
            .I(\c0.n1261 ));
    Odrv4 I__2255 (
            .O(N__13053),
            .I(\c0.n1261 ));
    CascadeMux I__2254 (
            .O(N__13046),
            .I(N__13041));
    InMux I__2253 (
            .O(N__13045),
            .I(N__13038));
    InMux I__2252 (
            .O(N__13044),
            .I(N__13035));
    InMux I__2251 (
            .O(N__13041),
            .I(N__13032));
    LocalMux I__2250 (
            .O(N__13038),
            .I(N__13028));
    LocalMux I__2249 (
            .O(N__13035),
            .I(N__13023));
    LocalMux I__2248 (
            .O(N__13032),
            .I(N__13023));
    InMux I__2247 (
            .O(N__13031),
            .I(N__13019));
    Span4Mux_h I__2246 (
            .O(N__13028),
            .I(N__13014));
    Span4Mux_h I__2245 (
            .O(N__13023),
            .I(N__13014));
    InMux I__2244 (
            .O(N__13022),
            .I(N__13011));
    LocalMux I__2243 (
            .O(N__13019),
            .I(\c0.data_in_field_45 ));
    Odrv4 I__2242 (
            .O(N__13014),
            .I(\c0.data_in_field_45 ));
    LocalMux I__2241 (
            .O(N__13011),
            .I(\c0.data_in_field_45 ));
    InMux I__2240 (
            .O(N__13004),
            .I(N__13001));
    LocalMux I__2239 (
            .O(N__13001),
            .I(N__12998));
    Odrv4 I__2238 (
            .O(N__12998),
            .I(\c0.n14 ));
    InMux I__2237 (
            .O(N__12995),
            .I(N__12992));
    LocalMux I__2236 (
            .O(N__12992),
            .I(N__12989));
    Span4Mux_h I__2235 (
            .O(N__12989),
            .I(N__12986));
    Odrv4 I__2234 (
            .O(N__12986),
            .I(\c0.n12_adj_873 ));
    CascadeMux I__2233 (
            .O(N__12983),
            .I(\c0.n16_cascade_ ));
    InMux I__2232 (
            .O(N__12980),
            .I(N__12977));
    LocalMux I__2231 (
            .O(N__12977),
            .I(N__12974));
    Span4Mux_h I__2230 (
            .O(N__12974),
            .I(N__12971));
    Span4Mux_v I__2229 (
            .O(N__12971),
            .I(N__12968));
    Odrv4 I__2228 (
            .O(N__12968),
            .I(\c0.n15 ));
    InMux I__2227 (
            .O(N__12965),
            .I(N__12962));
    LocalMux I__2226 (
            .O(N__12962),
            .I(\c0.n24 ));
    InMux I__2225 (
            .O(N__12959),
            .I(N__12956));
    LocalMux I__2224 (
            .O(N__12956),
            .I(\c0.n4388 ));
    CascadeMux I__2223 (
            .O(N__12953),
            .I(N__12950));
    InMux I__2222 (
            .O(N__12950),
            .I(N__12947));
    LocalMux I__2221 (
            .O(N__12947),
            .I(N__12944));
    Span4Mux_h I__2220 (
            .O(N__12944),
            .I(N__12941));
    Odrv4 I__2219 (
            .O(N__12941),
            .I(\c0.n4445 ));
    InMux I__2218 (
            .O(N__12938),
            .I(N__12935));
    LocalMux I__2217 (
            .O(N__12935),
            .I(\c0.n26_adj_890 ));
    InMux I__2216 (
            .O(N__12932),
            .I(N__12929));
    LocalMux I__2215 (
            .O(N__12929),
            .I(N__12925));
    InMux I__2214 (
            .O(N__12928),
            .I(N__12922));
    Span4Mux_h I__2213 (
            .O(N__12925),
            .I(N__12919));
    LocalMux I__2212 (
            .O(N__12922),
            .I(\c0.data_in_frame_6_2 ));
    Odrv4 I__2211 (
            .O(N__12919),
            .I(\c0.data_in_frame_6_2 ));
    InMux I__2210 (
            .O(N__12914),
            .I(N__12911));
    LocalMux I__2209 (
            .O(N__12911),
            .I(N__12908));
    Span4Mux_h I__2208 (
            .O(N__12908),
            .I(N__12905));
    Span4Mux_v I__2207 (
            .O(N__12905),
            .I(N__12902));
    Odrv4 I__2206 (
            .O(N__12902),
            .I(\c0.n1280 ));
    InMux I__2205 (
            .O(N__12899),
            .I(N__12896));
    LocalMux I__2204 (
            .O(N__12896),
            .I(N__12892));
    InMux I__2203 (
            .O(N__12895),
            .I(N__12889));
    Span4Mux_v I__2202 (
            .O(N__12892),
            .I(N__12886));
    LocalMux I__2201 (
            .O(N__12889),
            .I(N__12883));
    Odrv4 I__2200 (
            .O(N__12886),
            .I(\c0.n4390 ));
    Odrv4 I__2199 (
            .O(N__12883),
            .I(\c0.n4390 ));
    CascadeMux I__2198 (
            .O(N__12878),
            .I(N__12873));
    CascadeMux I__2197 (
            .O(N__12877),
            .I(N__12870));
    InMux I__2196 (
            .O(N__12876),
            .I(N__12867));
    InMux I__2195 (
            .O(N__12873),
            .I(N__12863));
    InMux I__2194 (
            .O(N__12870),
            .I(N__12860));
    LocalMux I__2193 (
            .O(N__12867),
            .I(N__12857));
    InMux I__2192 (
            .O(N__12866),
            .I(N__12854));
    LocalMux I__2191 (
            .O(N__12863),
            .I(N__12851));
    LocalMux I__2190 (
            .O(N__12860),
            .I(\c0.data_in_field_47 ));
    Odrv4 I__2189 (
            .O(N__12857),
            .I(\c0.data_in_field_47 ));
    LocalMux I__2188 (
            .O(N__12854),
            .I(\c0.data_in_field_47 ));
    Odrv4 I__2187 (
            .O(N__12851),
            .I(\c0.data_in_field_47 ));
    InMux I__2186 (
            .O(N__12842),
            .I(N__12839));
    LocalMux I__2185 (
            .O(N__12839),
            .I(\c0.n4391 ));
    InMux I__2184 (
            .O(N__12836),
            .I(N__12831));
    InMux I__2183 (
            .O(N__12835),
            .I(N__12828));
    CascadeMux I__2182 (
            .O(N__12834),
            .I(N__12825));
    LocalMux I__2181 (
            .O(N__12831),
            .I(N__12822));
    LocalMux I__2180 (
            .O(N__12828),
            .I(N__12819));
    InMux I__2179 (
            .O(N__12825),
            .I(N__12814));
    Span4Mux_v I__2178 (
            .O(N__12822),
            .I(N__12809));
    Span4Mux_h I__2177 (
            .O(N__12819),
            .I(N__12809));
    InMux I__2176 (
            .O(N__12818),
            .I(N__12806));
    InMux I__2175 (
            .O(N__12817),
            .I(N__12803));
    LocalMux I__2174 (
            .O(N__12814),
            .I(\c0.data_in_field_1 ));
    Odrv4 I__2173 (
            .O(N__12809),
            .I(\c0.data_in_field_1 ));
    LocalMux I__2172 (
            .O(N__12806),
            .I(\c0.data_in_field_1 ));
    LocalMux I__2171 (
            .O(N__12803),
            .I(\c0.data_in_field_1 ));
    CascadeMux I__2170 (
            .O(N__12794),
            .I(N__12791));
    InMux I__2169 (
            .O(N__12791),
            .I(N__12787));
    InMux I__2168 (
            .O(N__12790),
            .I(N__12783));
    LocalMux I__2167 (
            .O(N__12787),
            .I(N__12780));
    InMux I__2166 (
            .O(N__12786),
            .I(N__12776));
    LocalMux I__2165 (
            .O(N__12783),
            .I(N__12773));
    Span12Mux_v I__2164 (
            .O(N__12780),
            .I(N__12770));
    InMux I__2163 (
            .O(N__12779),
            .I(N__12767));
    LocalMux I__2162 (
            .O(N__12776),
            .I(\c0.data_in_field_14 ));
    Odrv12 I__2161 (
            .O(N__12773),
            .I(\c0.data_in_field_14 ));
    Odrv12 I__2160 (
            .O(N__12770),
            .I(\c0.data_in_field_14 ));
    LocalMux I__2159 (
            .O(N__12767),
            .I(\c0.data_in_field_14 ));
    InMux I__2158 (
            .O(N__12758),
            .I(N__12755));
    LocalMux I__2157 (
            .O(N__12755),
            .I(\c0.n4474 ));
    InMux I__2156 (
            .O(N__12752),
            .I(N__12749));
    LocalMux I__2155 (
            .O(N__12749),
            .I(\c0.n12_adj_887 ));
    InMux I__2154 (
            .O(N__12746),
            .I(\c0.n3922 ));
    SRMux I__2153 (
            .O(N__12743),
            .I(N__12740));
    LocalMux I__2152 (
            .O(N__12740),
            .I(N__12737));
    Odrv4 I__2151 (
            .O(N__12737),
            .I(\c0.n1675 ));
    CEMux I__2150 (
            .O(N__12734),
            .I(N__12731));
    LocalMux I__2149 (
            .O(N__12731),
            .I(N__12728));
    Odrv12 I__2148 (
            .O(N__12728),
            .I(\c0.n688 ));
    InMux I__2147 (
            .O(N__12725),
            .I(N__12720));
    InMux I__2146 (
            .O(N__12724),
            .I(N__12715));
    InMux I__2145 (
            .O(N__12723),
            .I(N__12715));
    LocalMux I__2144 (
            .O(N__12720),
            .I(tx2_active));
    LocalMux I__2143 (
            .O(N__12715),
            .I(tx2_active));
    InMux I__2142 (
            .O(N__12710),
            .I(N__12707));
    LocalMux I__2141 (
            .O(N__12707),
            .I(\c0.n2643 ));
    CascadeMux I__2140 (
            .O(N__12704),
            .I(\c0.n2643_cascade_ ));
    CascadeMux I__2139 (
            .O(N__12701),
            .I(N__12698));
    InMux I__2138 (
            .O(N__12698),
            .I(N__12695));
    LocalMux I__2137 (
            .O(N__12695),
            .I(N__12689));
    CascadeMux I__2136 (
            .O(N__12694),
            .I(N__12685));
    InMux I__2135 (
            .O(N__12693),
            .I(N__12680));
    InMux I__2134 (
            .O(N__12692),
            .I(N__12680));
    Span4Mux_h I__2133 (
            .O(N__12689),
            .I(N__12677));
    InMux I__2132 (
            .O(N__12688),
            .I(N__12672));
    InMux I__2131 (
            .O(N__12685),
            .I(N__12672));
    LocalMux I__2130 (
            .O(N__12680),
            .I(\c0.tx2_transmit ));
    Odrv4 I__2129 (
            .O(N__12677),
            .I(\c0.tx2_transmit ));
    LocalMux I__2128 (
            .O(N__12672),
            .I(\c0.tx2_transmit ));
    InMux I__2127 (
            .O(N__12665),
            .I(N__12662));
    LocalMux I__2126 (
            .O(N__12662),
            .I(\c0.n21 ));
    CascadeMux I__2125 (
            .O(N__12659),
            .I(N__12656));
    InMux I__2124 (
            .O(N__12656),
            .I(N__12653));
    LocalMux I__2123 (
            .O(N__12653),
            .I(\c0.n22_adj_881 ));
    CascadeMux I__2122 (
            .O(N__12650),
            .I(N__12645));
    CascadeMux I__2121 (
            .O(N__12649),
            .I(N__12641));
    InMux I__2120 (
            .O(N__12648),
            .I(N__12631));
    InMux I__2119 (
            .O(N__12645),
            .I(N__12631));
    InMux I__2118 (
            .O(N__12644),
            .I(N__12631));
    InMux I__2117 (
            .O(N__12641),
            .I(N__12628));
    InMux I__2116 (
            .O(N__12640),
            .I(N__12625));
    InMux I__2115 (
            .O(N__12639),
            .I(N__12620));
    CascadeMux I__2114 (
            .O(N__12638),
            .I(N__12616));
    LocalMux I__2113 (
            .O(N__12631),
            .I(N__12609));
    LocalMux I__2112 (
            .O(N__12628),
            .I(N__12609));
    LocalMux I__2111 (
            .O(N__12625),
            .I(N__12609));
    InMux I__2110 (
            .O(N__12624),
            .I(N__12604));
    InMux I__2109 (
            .O(N__12623),
            .I(N__12604));
    LocalMux I__2108 (
            .O(N__12620),
            .I(N__12601));
    InMux I__2107 (
            .O(N__12619),
            .I(N__12595));
    InMux I__2106 (
            .O(N__12616),
            .I(N__12595));
    Sp12to4 I__2105 (
            .O(N__12609),
            .I(N__12592));
    LocalMux I__2104 (
            .O(N__12604),
            .I(N__12587));
    Span12Mux_s2_v I__2103 (
            .O(N__12601),
            .I(N__12587));
    InMux I__2102 (
            .O(N__12600),
            .I(N__12584));
    LocalMux I__2101 (
            .O(N__12595),
            .I(N__12579));
    Span12Mux_v I__2100 (
            .O(N__12592),
            .I(N__12579));
    Odrv12 I__2099 (
            .O(N__12587),
            .I(r_SM_Main_0_adj_954));
    LocalMux I__2098 (
            .O(N__12584),
            .I(r_SM_Main_0_adj_954));
    Odrv12 I__2097 (
            .O(N__12579),
            .I(r_SM_Main_0_adj_954));
    CascadeMux I__2096 (
            .O(N__12572),
            .I(N__12566));
    InMux I__2095 (
            .O(N__12571),
            .I(N__12562));
    CascadeMux I__2094 (
            .O(N__12570),
            .I(N__12555));
    InMux I__2093 (
            .O(N__12569),
            .I(N__12550));
    InMux I__2092 (
            .O(N__12566),
            .I(N__12547));
    CascadeMux I__2091 (
            .O(N__12565),
            .I(N__12544));
    LocalMux I__2090 (
            .O(N__12562),
            .I(N__12541));
    InMux I__2089 (
            .O(N__12561),
            .I(N__12534));
    InMux I__2088 (
            .O(N__12560),
            .I(N__12534));
    InMux I__2087 (
            .O(N__12559),
            .I(N__12534));
    InMux I__2086 (
            .O(N__12558),
            .I(N__12529));
    InMux I__2085 (
            .O(N__12555),
            .I(N__12529));
    CascadeMux I__2084 (
            .O(N__12554),
            .I(N__12525));
    CascadeMux I__2083 (
            .O(N__12553),
            .I(N__12521));
    LocalMux I__2082 (
            .O(N__12550),
            .I(N__12518));
    LocalMux I__2081 (
            .O(N__12547),
            .I(N__12515));
    InMux I__2080 (
            .O(N__12544),
            .I(N__12512));
    Span12Mux_s5_v I__2079 (
            .O(N__12541),
            .I(N__12509));
    LocalMux I__2078 (
            .O(N__12534),
            .I(N__12504));
    LocalMux I__2077 (
            .O(N__12529),
            .I(N__12504));
    InMux I__2076 (
            .O(N__12528),
            .I(N__12501));
    InMux I__2075 (
            .O(N__12525),
            .I(N__12494));
    InMux I__2074 (
            .O(N__12524),
            .I(N__12494));
    InMux I__2073 (
            .O(N__12521),
            .I(N__12494));
    Span4Mux_v I__2072 (
            .O(N__12518),
            .I(N__12489));
    Span4Mux_v I__2071 (
            .O(N__12515),
            .I(N__12489));
    LocalMux I__2070 (
            .O(N__12512),
            .I(r_SM_Main_1_adj_953));
    Odrv12 I__2069 (
            .O(N__12509),
            .I(r_SM_Main_1_adj_953));
    Odrv4 I__2068 (
            .O(N__12504),
            .I(r_SM_Main_1_adj_953));
    LocalMux I__2067 (
            .O(N__12501),
            .I(r_SM_Main_1_adj_953));
    LocalMux I__2066 (
            .O(N__12494),
            .I(r_SM_Main_1_adj_953));
    Odrv4 I__2065 (
            .O(N__12489),
            .I(r_SM_Main_1_adj_953));
    InMux I__2064 (
            .O(N__12476),
            .I(N__12473));
    LocalMux I__2063 (
            .O(N__12473),
            .I(N__12470));
    Span4Mux_v I__2062 (
            .O(N__12470),
            .I(N__12467));
    Odrv4 I__2061 (
            .O(N__12467),
            .I(n4780));
    InMux I__2060 (
            .O(N__12464),
            .I(N__12450));
    InMux I__2059 (
            .O(N__12463),
            .I(N__12450));
    CascadeMux I__2058 (
            .O(N__12462),
            .I(N__12445));
    CascadeMux I__2057 (
            .O(N__12461),
            .I(N__12442));
    CascadeMux I__2056 (
            .O(N__12460),
            .I(N__12439));
    CascadeMux I__2055 (
            .O(N__12459),
            .I(N__12436));
    CascadeMux I__2054 (
            .O(N__12458),
            .I(N__12433));
    CascadeMux I__2053 (
            .O(N__12457),
            .I(N__12430));
    CascadeMux I__2052 (
            .O(N__12456),
            .I(N__12427));
    CascadeMux I__2051 (
            .O(N__12455),
            .I(N__12424));
    LocalMux I__2050 (
            .O(N__12450),
            .I(N__12421));
    InMux I__2049 (
            .O(N__12449),
            .I(N__12418));
    CascadeMux I__2048 (
            .O(N__12448),
            .I(N__12415));
    InMux I__2047 (
            .O(N__12445),
            .I(N__12398));
    InMux I__2046 (
            .O(N__12442),
            .I(N__12398));
    InMux I__2045 (
            .O(N__12439),
            .I(N__12398));
    InMux I__2044 (
            .O(N__12436),
            .I(N__12398));
    InMux I__2043 (
            .O(N__12433),
            .I(N__12389));
    InMux I__2042 (
            .O(N__12430),
            .I(N__12389));
    InMux I__2041 (
            .O(N__12427),
            .I(N__12389));
    InMux I__2040 (
            .O(N__12424),
            .I(N__12389));
    Sp12to4 I__2039 (
            .O(N__12421),
            .I(N__12384));
    LocalMux I__2038 (
            .O(N__12418),
            .I(N__12384));
    InMux I__2037 (
            .O(N__12415),
            .I(N__12381));
    InMux I__2036 (
            .O(N__12414),
            .I(N__12378));
    InMux I__2035 (
            .O(N__12413),
            .I(N__12371));
    InMux I__2034 (
            .O(N__12412),
            .I(N__12371));
    InMux I__2033 (
            .O(N__12411),
            .I(N__12371));
    InMux I__2032 (
            .O(N__12410),
            .I(N__12368));
    InMux I__2031 (
            .O(N__12409),
            .I(N__12361));
    InMux I__2030 (
            .O(N__12408),
            .I(N__12361));
    InMux I__2029 (
            .O(N__12407),
            .I(N__12361));
    LocalMux I__2028 (
            .O(N__12398),
            .I(N__12356));
    LocalMux I__2027 (
            .O(N__12389),
            .I(N__12356));
    Odrv12 I__2026 (
            .O(N__12384),
            .I(r_SM_Main_2_adj_952));
    LocalMux I__2025 (
            .O(N__12381),
            .I(r_SM_Main_2_adj_952));
    LocalMux I__2024 (
            .O(N__12378),
            .I(r_SM_Main_2_adj_952));
    LocalMux I__2023 (
            .O(N__12371),
            .I(r_SM_Main_2_adj_952));
    LocalMux I__2022 (
            .O(N__12368),
            .I(r_SM_Main_2_adj_952));
    LocalMux I__2021 (
            .O(N__12361),
            .I(r_SM_Main_2_adj_952));
    Odrv4 I__2020 (
            .O(N__12356),
            .I(r_SM_Main_2_adj_952));
    CascadeMux I__2019 (
            .O(N__12341),
            .I(n3_cascade_));
    InMux I__2018 (
            .O(N__12338),
            .I(N__12335));
    LocalMux I__2017 (
            .O(N__12335),
            .I(N__12331));
    InMux I__2016 (
            .O(N__12334),
            .I(N__12328));
    Odrv12 I__2015 (
            .O(N__12331),
            .I(rx_data_6));
    LocalMux I__2014 (
            .O(N__12328),
            .I(rx_data_6));
    InMux I__2013 (
            .O(N__12323),
            .I(N__12320));
    LocalMux I__2012 (
            .O(N__12320),
            .I(\c0.rx.n4876 ));
    IoInMux I__2011 (
            .O(N__12317),
            .I(N__12314));
    LocalMux I__2010 (
            .O(N__12314),
            .I(tx_enable));
    CascadeMux I__2009 (
            .O(N__12311),
            .I(N__12305));
    CascadeMux I__2008 (
            .O(N__12310),
            .I(N__12302));
    InMux I__2007 (
            .O(N__12309),
            .I(N__12299));
    InMux I__2006 (
            .O(N__12308),
            .I(N__12296));
    InMux I__2005 (
            .O(N__12305),
            .I(N__12291));
    InMux I__2004 (
            .O(N__12302),
            .I(N__12291));
    LocalMux I__2003 (
            .O(N__12299),
            .I(data_in_7_5));
    LocalMux I__2002 (
            .O(N__12296),
            .I(data_in_7_5));
    LocalMux I__2001 (
            .O(N__12291),
            .I(data_in_7_5));
    InMux I__2000 (
            .O(N__12284),
            .I(N__12280));
    InMux I__1999 (
            .O(N__12283),
            .I(N__12277));
    LocalMux I__1998 (
            .O(N__12280),
            .I(N__12274));
    LocalMux I__1997 (
            .O(N__12277),
            .I(N__12269));
    Span4Mux_s3_h I__1996 (
            .O(N__12274),
            .I(N__12266));
    InMux I__1995 (
            .O(N__12273),
            .I(N__12263));
    InMux I__1994 (
            .O(N__12272),
            .I(N__12260));
    Span4Mux_v I__1993 (
            .O(N__12269),
            .I(N__12257));
    Odrv4 I__1992 (
            .O(N__12266),
            .I(data_in_6_5));
    LocalMux I__1991 (
            .O(N__12263),
            .I(data_in_6_5));
    LocalMux I__1990 (
            .O(N__12260),
            .I(data_in_6_5));
    Odrv4 I__1989 (
            .O(N__12257),
            .I(data_in_6_5));
    InMux I__1988 (
            .O(N__12248),
            .I(N__12245));
    LocalMux I__1987 (
            .O(N__12245),
            .I(n4519));
    InMux I__1986 (
            .O(N__12242),
            .I(N__12239));
    LocalMux I__1985 (
            .O(N__12239),
            .I(n4520));
    InMux I__1984 (
            .O(N__12236),
            .I(N__12233));
    LocalMux I__1983 (
            .O(N__12233),
            .I(N__12230));
    Span4Mux_v I__1982 (
            .O(N__12230),
            .I(N__12226));
    InMux I__1981 (
            .O(N__12229),
            .I(N__12223));
    Odrv4 I__1980 (
            .O(N__12226),
            .I(blink_counter_25));
    LocalMux I__1979 (
            .O(N__12223),
            .I(blink_counter_25));
    IoInMux I__1978 (
            .O(N__12218),
            .I(N__12215));
    LocalMux I__1977 (
            .O(N__12215),
            .I(N__12212));
    Span12Mux_s9_v I__1976 (
            .O(N__12212),
            .I(N__12209));
    Odrv12 I__1975 (
            .O(N__12209),
            .I(LED_c));
    InMux I__1974 (
            .O(N__12206),
            .I(\c0.n3921 ));
    InMux I__1973 (
            .O(N__12203),
            .I(N__12199));
    InMux I__1972 (
            .O(N__12202),
            .I(N__12196));
    LocalMux I__1971 (
            .O(N__12199),
            .I(\c0.data_in_frame_6_1 ));
    LocalMux I__1970 (
            .O(N__12196),
            .I(\c0.data_in_frame_6_1 ));
    InMux I__1969 (
            .O(N__12191),
            .I(N__12187));
    CascadeMux I__1968 (
            .O(N__12190),
            .I(N__12184));
    LocalMux I__1967 (
            .O(N__12187),
            .I(N__12181));
    InMux I__1966 (
            .O(N__12184),
            .I(N__12177));
    Span4Mux_v I__1965 (
            .O(N__12181),
            .I(N__12174));
    InMux I__1964 (
            .O(N__12180),
            .I(N__12171));
    LocalMux I__1963 (
            .O(N__12177),
            .I(data_in_5_4));
    Odrv4 I__1962 (
            .O(N__12174),
            .I(data_in_5_4));
    LocalMux I__1961 (
            .O(N__12171),
            .I(data_in_5_4));
    InMux I__1960 (
            .O(N__12164),
            .I(N__12160));
    InMux I__1959 (
            .O(N__12163),
            .I(N__12156));
    LocalMux I__1958 (
            .O(N__12160),
            .I(N__12153));
    InMux I__1957 (
            .O(N__12159),
            .I(N__12150));
    LocalMux I__1956 (
            .O(N__12156),
            .I(\c0.data_in_field_44 ));
    Odrv12 I__1955 (
            .O(N__12153),
            .I(\c0.data_in_field_44 ));
    LocalMux I__1954 (
            .O(N__12150),
            .I(\c0.data_in_field_44 ));
    CascadeMux I__1953 (
            .O(N__12143),
            .I(N__12140));
    InMux I__1952 (
            .O(N__12140),
            .I(N__12134));
    InMux I__1951 (
            .O(N__12139),
            .I(N__12131));
    InMux I__1950 (
            .O(N__12138),
            .I(N__12128));
    InMux I__1949 (
            .O(N__12137),
            .I(N__12125));
    LocalMux I__1948 (
            .O(N__12134),
            .I(N__12122));
    LocalMux I__1947 (
            .O(N__12131),
            .I(data_in_3_4));
    LocalMux I__1946 (
            .O(N__12128),
            .I(data_in_3_4));
    LocalMux I__1945 (
            .O(N__12125),
            .I(data_in_3_4));
    Odrv12 I__1944 (
            .O(N__12122),
            .I(data_in_3_4));
    InMux I__1943 (
            .O(N__12113),
            .I(N__12109));
    InMux I__1942 (
            .O(N__12112),
            .I(N__12106));
    LocalMux I__1941 (
            .O(N__12109),
            .I(N__12101));
    LocalMux I__1940 (
            .O(N__12106),
            .I(N__12098));
    InMux I__1939 (
            .O(N__12105),
            .I(N__12095));
    InMux I__1938 (
            .O(N__12104),
            .I(N__12092));
    Span4Mux_s3_h I__1937 (
            .O(N__12101),
            .I(N__12089));
    Span4Mux_s1_h I__1936 (
            .O(N__12098),
            .I(N__12084));
    LocalMux I__1935 (
            .O(N__12095),
            .I(N__12084));
    LocalMux I__1934 (
            .O(N__12092),
            .I(data_in_2_4));
    Odrv4 I__1933 (
            .O(N__12089),
            .I(data_in_2_4));
    Odrv4 I__1932 (
            .O(N__12084),
            .I(data_in_2_4));
    CascadeMux I__1931 (
            .O(N__12077),
            .I(N__12074));
    InMux I__1930 (
            .O(N__12074),
            .I(N__12068));
    InMux I__1929 (
            .O(N__12073),
            .I(N__12068));
    LocalMux I__1928 (
            .O(N__12068),
            .I(rx_data_5));
    InMux I__1927 (
            .O(N__12065),
            .I(N__12061));
    CascadeMux I__1926 (
            .O(N__12064),
            .I(N__12058));
    LocalMux I__1925 (
            .O(N__12061),
            .I(N__12055));
    InMux I__1924 (
            .O(N__12058),
            .I(N__12052));
    Odrv12 I__1923 (
            .O(N__12055),
            .I(rx_data_7));
    LocalMux I__1922 (
            .O(N__12052),
            .I(rx_data_7));
    CascadeMux I__1921 (
            .O(N__12047),
            .I(N__12043));
    InMux I__1920 (
            .O(N__12046),
            .I(N__12039));
    InMux I__1919 (
            .O(N__12043),
            .I(N__12034));
    InMux I__1918 (
            .O(N__12042),
            .I(N__12031));
    LocalMux I__1917 (
            .O(N__12039),
            .I(N__12028));
    InMux I__1916 (
            .O(N__12038),
            .I(N__12023));
    InMux I__1915 (
            .O(N__12037),
            .I(N__12023));
    LocalMux I__1914 (
            .O(N__12034),
            .I(N__12020));
    LocalMux I__1913 (
            .O(N__12031),
            .I(N__12017));
    Odrv4 I__1912 (
            .O(N__12028),
            .I(\c0.data_in_field_39 ));
    LocalMux I__1911 (
            .O(N__12023),
            .I(\c0.data_in_field_39 ));
    Odrv4 I__1910 (
            .O(N__12020),
            .I(\c0.data_in_field_39 ));
    Odrv4 I__1909 (
            .O(N__12017),
            .I(\c0.data_in_field_39 ));
    InMux I__1908 (
            .O(N__12008),
            .I(N__12004));
    InMux I__1907 (
            .O(N__12007),
            .I(N__11999));
    LocalMux I__1906 (
            .O(N__12004),
            .I(N__11996));
    InMux I__1905 (
            .O(N__12003),
            .I(N__11991));
    InMux I__1904 (
            .O(N__12002),
            .I(N__11991));
    LocalMux I__1903 (
            .O(N__11999),
            .I(\c0.data_in_field_38 ));
    Odrv4 I__1902 (
            .O(N__11996),
            .I(\c0.data_in_field_38 ));
    LocalMux I__1901 (
            .O(N__11991),
            .I(\c0.data_in_field_38 ));
    InMux I__1900 (
            .O(N__11984),
            .I(N__11980));
    InMux I__1899 (
            .O(N__11983),
            .I(N__11975));
    LocalMux I__1898 (
            .O(N__11980),
            .I(N__11972));
    InMux I__1897 (
            .O(N__11979),
            .I(N__11969));
    InMux I__1896 (
            .O(N__11978),
            .I(N__11966));
    LocalMux I__1895 (
            .O(N__11975),
            .I(N__11963));
    Span4Mux_s3_h I__1894 (
            .O(N__11972),
            .I(N__11960));
    LocalMux I__1893 (
            .O(N__11969),
            .I(N__11957));
    LocalMux I__1892 (
            .O(N__11966),
            .I(data_in_6_4));
    Odrv4 I__1891 (
            .O(N__11963),
            .I(data_in_6_4));
    Odrv4 I__1890 (
            .O(N__11960),
            .I(data_in_6_4));
    Odrv12 I__1889 (
            .O(N__11957),
            .I(data_in_6_4));
    InMux I__1888 (
            .O(N__11948),
            .I(N__11945));
    LocalMux I__1887 (
            .O(N__11945),
            .I(N__11940));
    InMux I__1886 (
            .O(N__11944),
            .I(N__11935));
    InMux I__1885 (
            .O(N__11943),
            .I(N__11935));
    Span4Mux_s3_h I__1884 (
            .O(N__11940),
            .I(N__11932));
    LocalMux I__1883 (
            .O(N__11935),
            .I(data_in_4_4));
    Odrv4 I__1882 (
            .O(N__11932),
            .I(data_in_4_4));
    InMux I__1881 (
            .O(N__11927),
            .I(N__11924));
    LocalMux I__1880 (
            .O(N__11924),
            .I(\c0.n8_adj_872 ));
    InMux I__1879 (
            .O(N__11921),
            .I(N__11918));
    LocalMux I__1878 (
            .O(N__11918),
            .I(N__11914));
    CascadeMux I__1877 (
            .O(N__11917),
            .I(N__11910));
    Span4Mux_h I__1876 (
            .O(N__11914),
            .I(N__11907));
    InMux I__1875 (
            .O(N__11913),
            .I(N__11902));
    InMux I__1874 (
            .O(N__11910),
            .I(N__11902));
    Odrv4 I__1873 (
            .O(N__11907),
            .I(data_in_0_2));
    LocalMux I__1872 (
            .O(N__11902),
            .I(data_in_0_2));
    InMux I__1871 (
            .O(N__11897),
            .I(N__11893));
    InMux I__1870 (
            .O(N__11896),
            .I(N__11888));
    LocalMux I__1869 (
            .O(N__11893),
            .I(N__11885));
    InMux I__1868 (
            .O(N__11892),
            .I(N__11882));
    InMux I__1867 (
            .O(N__11891),
            .I(N__11879));
    LocalMux I__1866 (
            .O(N__11888),
            .I(\c0.data_in_field_2 ));
    Odrv12 I__1865 (
            .O(N__11885),
            .I(\c0.data_in_field_2 ));
    LocalMux I__1864 (
            .O(N__11882),
            .I(\c0.data_in_field_2 ));
    LocalMux I__1863 (
            .O(N__11879),
            .I(\c0.data_in_field_2 ));
    CascadeMux I__1862 (
            .O(N__11870),
            .I(N__11867));
    InMux I__1861 (
            .O(N__11867),
            .I(N__11861));
    InMux I__1860 (
            .O(N__11866),
            .I(N__11861));
    LocalMux I__1859 (
            .O(N__11861),
            .I(\c0.data_in_frame_7_1 ));
    InMux I__1858 (
            .O(N__11858),
            .I(N__11855));
    LocalMux I__1857 (
            .O(N__11855),
            .I(N__11852));
    Span4Mux_s3_h I__1856 (
            .O(N__11852),
            .I(N__11849));
    Span4Mux_v I__1855 (
            .O(N__11849),
            .I(N__11846));
    Odrv4 I__1854 (
            .O(N__11846),
            .I(\c0.n4607 ));
    InMux I__1853 (
            .O(N__11843),
            .I(N__11840));
    LocalMux I__1852 (
            .O(N__11840),
            .I(N__11835));
    InMux I__1851 (
            .O(N__11839),
            .I(N__11829));
    InMux I__1850 (
            .O(N__11838),
            .I(N__11829));
    Span4Mux_v I__1849 (
            .O(N__11835),
            .I(N__11826));
    InMux I__1848 (
            .O(N__11834),
            .I(N__11823));
    LocalMux I__1847 (
            .O(N__11829),
            .I(N__11820));
    Odrv4 I__1846 (
            .O(N__11826),
            .I(data_in_3_6));
    LocalMux I__1845 (
            .O(N__11823),
            .I(data_in_3_6));
    Odrv12 I__1844 (
            .O(N__11820),
            .I(data_in_3_6));
    CascadeMux I__1843 (
            .O(N__11813),
            .I(N__11810));
    InMux I__1842 (
            .O(N__11810),
            .I(N__11807));
    LocalMux I__1841 (
            .O(N__11807),
            .I(N__11802));
    InMux I__1840 (
            .O(N__11806),
            .I(N__11798));
    InMux I__1839 (
            .O(N__11805),
            .I(N__11795));
    Span4Mux_h I__1838 (
            .O(N__11802),
            .I(N__11792));
    InMux I__1837 (
            .O(N__11801),
            .I(N__11789));
    LocalMux I__1836 (
            .O(N__11798),
            .I(data_in_1_1));
    LocalMux I__1835 (
            .O(N__11795),
            .I(data_in_1_1));
    Odrv4 I__1834 (
            .O(N__11792),
            .I(data_in_1_1));
    LocalMux I__1833 (
            .O(N__11789),
            .I(data_in_1_1));
    CascadeMux I__1832 (
            .O(N__11780),
            .I(\c0.n8_adj_871_cascade_ ));
    InMux I__1831 (
            .O(N__11777),
            .I(N__11774));
    LocalMux I__1830 (
            .O(N__11774),
            .I(\c0.n12 ));
    InMux I__1829 (
            .O(N__11771),
            .I(N__11768));
    LocalMux I__1828 (
            .O(N__11768),
            .I(\c0.n1418 ));
    InMux I__1827 (
            .O(N__11765),
            .I(N__11762));
    LocalMux I__1826 (
            .O(N__11762),
            .I(N__11758));
    InMux I__1825 (
            .O(N__11761),
            .I(N__11752));
    Span4Mux_v I__1824 (
            .O(N__11758),
            .I(N__11749));
    InMux I__1823 (
            .O(N__11757),
            .I(N__11746));
    InMux I__1822 (
            .O(N__11756),
            .I(N__11743));
    InMux I__1821 (
            .O(N__11755),
            .I(N__11740));
    LocalMux I__1820 (
            .O(N__11752),
            .I(\c0.data_in_field_4 ));
    Odrv4 I__1819 (
            .O(N__11749),
            .I(\c0.data_in_field_4 ));
    LocalMux I__1818 (
            .O(N__11746),
            .I(\c0.data_in_field_4 ));
    LocalMux I__1817 (
            .O(N__11743),
            .I(\c0.data_in_field_4 ));
    LocalMux I__1816 (
            .O(N__11740),
            .I(\c0.data_in_field_4 ));
    CascadeMux I__1815 (
            .O(N__11729),
            .I(\c0.n1418_cascade_ ));
    CascadeMux I__1814 (
            .O(N__11726),
            .I(\c0.n4474_cascade_ ));
    InMux I__1813 (
            .O(N__11723),
            .I(N__11720));
    LocalMux I__1812 (
            .O(N__11720),
            .I(N__11717));
    Span4Mux_h I__1811 (
            .O(N__11717),
            .I(N__11712));
    InMux I__1810 (
            .O(N__11716),
            .I(N__11707));
    InMux I__1809 (
            .O(N__11715),
            .I(N__11707));
    Odrv4 I__1808 (
            .O(N__11712),
            .I(data_in_4_6));
    LocalMux I__1807 (
            .O(N__11707),
            .I(data_in_4_6));
    InMux I__1806 (
            .O(N__11702),
            .I(N__11699));
    LocalMux I__1805 (
            .O(N__11699),
            .I(N__11696));
    Odrv12 I__1804 (
            .O(N__11696),
            .I(\c0.n4396 ));
    InMux I__1803 (
            .O(N__11693),
            .I(N__11689));
    InMux I__1802 (
            .O(N__11692),
            .I(N__11686));
    LocalMux I__1801 (
            .O(N__11689),
            .I(N__11681));
    LocalMux I__1800 (
            .O(N__11686),
            .I(N__11678));
    InMux I__1799 (
            .O(N__11685),
            .I(N__11673));
    InMux I__1798 (
            .O(N__11684),
            .I(N__11673));
    Odrv4 I__1797 (
            .O(N__11681),
            .I(\c0.data_in_field_21 ));
    Odrv4 I__1796 (
            .O(N__11678),
            .I(\c0.data_in_field_21 ));
    LocalMux I__1795 (
            .O(N__11673),
            .I(\c0.data_in_field_21 ));
    CascadeMux I__1794 (
            .O(N__11666),
            .I(\c0.n4396_cascade_ ));
    CascadeMux I__1793 (
            .O(N__11663),
            .I(N__11658));
    InMux I__1792 (
            .O(N__11662),
            .I(N__11655));
    InMux I__1791 (
            .O(N__11661),
            .I(N__11649));
    InMux I__1790 (
            .O(N__11658),
            .I(N__11649));
    LocalMux I__1789 (
            .O(N__11655),
            .I(N__11646));
    InMux I__1788 (
            .O(N__11654),
            .I(N__11643));
    LocalMux I__1787 (
            .O(N__11649),
            .I(\c0.data_in_field_7 ));
    Odrv4 I__1786 (
            .O(N__11646),
            .I(\c0.data_in_field_7 ));
    LocalMux I__1785 (
            .O(N__11643),
            .I(\c0.data_in_field_7 ));
    InMux I__1784 (
            .O(N__11636),
            .I(N__11632));
    InMux I__1783 (
            .O(N__11635),
            .I(N__11628));
    LocalMux I__1782 (
            .O(N__11632),
            .I(N__11625));
    InMux I__1781 (
            .O(N__11631),
            .I(N__11621));
    LocalMux I__1780 (
            .O(N__11628),
            .I(N__11618));
    Span4Mux_h I__1779 (
            .O(N__11625),
            .I(N__11615));
    InMux I__1778 (
            .O(N__11624),
            .I(N__11612));
    LocalMux I__1777 (
            .O(N__11621),
            .I(\c0.data_in_field_0 ));
    Odrv4 I__1776 (
            .O(N__11618),
            .I(\c0.data_in_field_0 ));
    Odrv4 I__1775 (
            .O(N__11615),
            .I(\c0.data_in_field_0 ));
    LocalMux I__1774 (
            .O(N__11612),
            .I(\c0.data_in_field_0 ));
    InMux I__1773 (
            .O(N__11603),
            .I(N__11597));
    InMux I__1772 (
            .O(N__11602),
            .I(N__11597));
    LocalMux I__1771 (
            .O(N__11597),
            .I(N__11593));
    InMux I__1770 (
            .O(N__11596),
            .I(N__11589));
    Span4Mux_v I__1769 (
            .O(N__11593),
            .I(N__11586));
    InMux I__1768 (
            .O(N__11592),
            .I(N__11583));
    LocalMux I__1767 (
            .O(N__11589),
            .I(\c0.data_in_field_8 ));
    Odrv4 I__1766 (
            .O(N__11586),
            .I(\c0.data_in_field_8 ));
    LocalMux I__1765 (
            .O(N__11583),
            .I(\c0.data_in_field_8 ));
    InMux I__1764 (
            .O(N__11576),
            .I(N__11573));
    LocalMux I__1763 (
            .O(N__11573),
            .I(N__11570));
    Span4Mux_v I__1762 (
            .O(N__11570),
            .I(N__11567));
    Odrv4 I__1761 (
            .O(N__11567),
            .I(\c0.n4570 ));
    InMux I__1760 (
            .O(N__11564),
            .I(N__11561));
    LocalMux I__1759 (
            .O(N__11561),
            .I(\c0.n17 ));
    InMux I__1758 (
            .O(N__11558),
            .I(N__11555));
    LocalMux I__1757 (
            .O(N__11555),
            .I(\c0.n4430 ));
    CascadeMux I__1756 (
            .O(N__11552),
            .I(N__11549));
    InMux I__1755 (
            .O(N__11549),
            .I(N__11546));
    LocalMux I__1754 (
            .O(N__11546),
            .I(\c0.n15_adj_885 ));
    InMux I__1753 (
            .O(N__11543),
            .I(N__11540));
    LocalMux I__1752 (
            .O(N__11540),
            .I(\c0.n16_adj_884 ));
    CascadeMux I__1751 (
            .O(N__11537),
            .I(\c0.n17_adj_889_cascade_ ));
    CascadeMux I__1750 (
            .O(N__11534),
            .I(\c0.n4387_cascade_ ));
    InMux I__1749 (
            .O(N__11531),
            .I(N__11527));
    CascadeMux I__1748 (
            .O(N__11530),
            .I(N__11524));
    LocalMux I__1747 (
            .O(N__11527),
            .I(N__11521));
    InMux I__1746 (
            .O(N__11524),
            .I(N__11518));
    Span4Mux_s1_v I__1745 (
            .O(N__11521),
            .I(N__11515));
    LocalMux I__1744 (
            .O(N__11518),
            .I(N__11511));
    Span4Mux_v I__1743 (
            .O(N__11515),
            .I(N__11508));
    InMux I__1742 (
            .O(N__11514),
            .I(N__11505));
    Odrv12 I__1741 (
            .O(N__11511),
            .I(data_in_4_7));
    Odrv4 I__1740 (
            .O(N__11508),
            .I(data_in_4_7));
    LocalMux I__1739 (
            .O(N__11505),
            .I(data_in_4_7));
    InMux I__1738 (
            .O(N__11498),
            .I(N__11494));
    InMux I__1737 (
            .O(N__11497),
            .I(N__11491));
    LocalMux I__1736 (
            .O(N__11494),
            .I(N__11488));
    LocalMux I__1735 (
            .O(N__11491),
            .I(N__11482));
    Span4Mux_s3_h I__1734 (
            .O(N__11488),
            .I(N__11482));
    InMux I__1733 (
            .O(N__11487),
            .I(N__11479));
    Odrv4 I__1732 (
            .O(N__11482),
            .I(data_in_5_7));
    LocalMux I__1731 (
            .O(N__11479),
            .I(data_in_5_7));
    InMux I__1730 (
            .O(N__11474),
            .I(N__11471));
    LocalMux I__1729 (
            .O(N__11471),
            .I(N__11466));
    InMux I__1728 (
            .O(N__11470),
            .I(N__11461));
    InMux I__1727 (
            .O(N__11469),
            .I(N__11461));
    Span4Mux_s3_h I__1726 (
            .O(N__11466),
            .I(N__11458));
    LocalMux I__1725 (
            .O(N__11461),
            .I(\c0.n1296 ));
    Odrv4 I__1724 (
            .O(N__11458),
            .I(\c0.n1296 ));
    InMux I__1723 (
            .O(N__11453),
            .I(N__11450));
    LocalMux I__1722 (
            .O(N__11450),
            .I(\c0.n11_adj_888 ));
    CascadeMux I__1721 (
            .O(N__11447),
            .I(N__11444));
    InMux I__1720 (
            .O(N__11444),
            .I(N__11441));
    LocalMux I__1719 (
            .O(N__11441),
            .I(N__11436));
    CascadeMux I__1718 (
            .O(N__11440),
            .I(N__11432));
    InMux I__1717 (
            .O(N__11439),
            .I(N__11429));
    Span4Mux_h I__1716 (
            .O(N__11436),
            .I(N__11426));
    InMux I__1715 (
            .O(N__11435),
            .I(N__11421));
    InMux I__1714 (
            .O(N__11432),
            .I(N__11421));
    LocalMux I__1713 (
            .O(N__11429),
            .I(data_in_2_7));
    Odrv4 I__1712 (
            .O(N__11426),
            .I(data_in_2_7));
    LocalMux I__1711 (
            .O(N__11421),
            .I(data_in_2_7));
    InMux I__1710 (
            .O(N__11414),
            .I(N__11404));
    InMux I__1709 (
            .O(N__11413),
            .I(N__11404));
    InMux I__1708 (
            .O(N__11412),
            .I(N__11404));
    InMux I__1707 (
            .O(N__11411),
            .I(N__11400));
    LocalMux I__1706 (
            .O(N__11404),
            .I(N__11397));
    InMux I__1705 (
            .O(N__11403),
            .I(N__11394));
    LocalMux I__1704 (
            .O(N__11400),
            .I(r_SM_Main_2_N_759_1));
    Odrv12 I__1703 (
            .O(N__11397),
            .I(r_SM_Main_2_N_759_1));
    LocalMux I__1702 (
            .O(N__11394),
            .I(r_SM_Main_2_N_759_1));
    CascadeMux I__1701 (
            .O(N__11387),
            .I(n4366_cascade_));
    InMux I__1700 (
            .O(N__11384),
            .I(N__11380));
    InMux I__1699 (
            .O(N__11383),
            .I(N__11377));
    LocalMux I__1698 (
            .O(N__11380),
            .I(N__11374));
    LocalMux I__1697 (
            .O(N__11377),
            .I(N__11370));
    Span4Mux_v I__1696 (
            .O(N__11374),
            .I(N__11367));
    InMux I__1695 (
            .O(N__11373),
            .I(N__11364));
    Odrv4 I__1694 (
            .O(N__11370),
            .I(data_in_4_2));
    Odrv4 I__1693 (
            .O(N__11367),
            .I(data_in_4_2));
    LocalMux I__1692 (
            .O(N__11364),
            .I(data_in_4_2));
    InMux I__1691 (
            .O(N__11357),
            .I(N__11352));
    InMux I__1690 (
            .O(N__11356),
            .I(N__11349));
    CascadeMux I__1689 (
            .O(N__11355),
            .I(N__11346));
    LocalMux I__1688 (
            .O(N__11352),
            .I(N__11343));
    LocalMux I__1687 (
            .O(N__11349),
            .I(N__11340));
    InMux I__1686 (
            .O(N__11346),
            .I(N__11335));
    Span4Mux_v I__1685 (
            .O(N__11343),
            .I(N__11332));
    Span4Mux_v I__1684 (
            .O(N__11340),
            .I(N__11329));
    InMux I__1683 (
            .O(N__11339),
            .I(N__11326));
    InMux I__1682 (
            .O(N__11338),
            .I(N__11323));
    LocalMux I__1681 (
            .O(N__11335),
            .I(\c0.data_in_field_11 ));
    Odrv4 I__1680 (
            .O(N__11332),
            .I(\c0.data_in_field_11 ));
    Odrv4 I__1679 (
            .O(N__11329),
            .I(\c0.data_in_field_11 ));
    LocalMux I__1678 (
            .O(N__11326),
            .I(\c0.data_in_field_11 ));
    LocalMux I__1677 (
            .O(N__11323),
            .I(\c0.data_in_field_11 ));
    CascadeMux I__1676 (
            .O(N__11312),
            .I(\c0.n8_adj_879_cascade_ ));
    CascadeMux I__1675 (
            .O(N__11309),
            .I(\c0.n4451_cascade_ ));
    InMux I__1674 (
            .O(N__11306),
            .I(N__11303));
    LocalMux I__1673 (
            .O(N__11303),
            .I(N__11300));
    Odrv4 I__1672 (
            .O(N__11300),
            .I(\c0.n8_adj_880 ));
    InMux I__1671 (
            .O(N__11297),
            .I(N__11294));
    LocalMux I__1670 (
            .O(N__11294),
            .I(N__11291));
    Odrv12 I__1669 (
            .O(N__11291),
            .I(\c0.n10_adj_876 ));
    InMux I__1668 (
            .O(N__11288),
            .I(N__11285));
    LocalMux I__1667 (
            .O(N__11285),
            .I(\c0.n4469 ));
    CascadeMux I__1666 (
            .O(N__11282),
            .I(\c0.n1357_cascade_ ));
    InMux I__1665 (
            .O(N__11279),
            .I(N__11276));
    LocalMux I__1664 (
            .O(N__11276),
            .I(N__11273));
    Span4Mux_h I__1663 (
            .O(N__11273),
            .I(N__11269));
    InMux I__1662 (
            .O(N__11272),
            .I(N__11266));
    Odrv4 I__1661 (
            .O(N__11269),
            .I(\c0.n4399 ));
    LocalMux I__1660 (
            .O(N__11266),
            .I(\c0.n4399 ));
    InMux I__1659 (
            .O(N__11261),
            .I(N__11258));
    LocalMux I__1658 (
            .O(N__11258),
            .I(\c0.n4819 ));
    CascadeMux I__1657 (
            .O(N__11255),
            .I(\c0.n4549_cascade_ ));
    InMux I__1656 (
            .O(N__11252),
            .I(N__11249));
    LocalMux I__1655 (
            .O(N__11249),
            .I(N__11243));
    InMux I__1654 (
            .O(N__11248),
            .I(N__11236));
    InMux I__1653 (
            .O(N__11247),
            .I(N__11236));
    InMux I__1652 (
            .O(N__11246),
            .I(N__11236));
    Span4Mux_v I__1651 (
            .O(N__11243),
            .I(N__11231));
    LocalMux I__1650 (
            .O(N__11236),
            .I(N__11231));
    Span4Mux_v I__1649 (
            .O(N__11231),
            .I(N__11224));
    InMux I__1648 (
            .O(N__11230),
            .I(N__11219));
    InMux I__1647 (
            .O(N__11229),
            .I(N__11219));
    InMux I__1646 (
            .O(N__11228),
            .I(N__11216));
    InMux I__1645 (
            .O(N__11227),
            .I(N__11213));
    Odrv4 I__1644 (
            .O(N__11224),
            .I(n1030));
    LocalMux I__1643 (
            .O(N__11219),
            .I(n1030));
    LocalMux I__1642 (
            .O(N__11216),
            .I(n1030));
    LocalMux I__1641 (
            .O(N__11213),
            .I(n1030));
    CascadeMux I__1640 (
            .O(N__11204),
            .I(tx2_data_4_keep_cascade_));
    InMux I__1639 (
            .O(N__11201),
            .I(N__11197));
    InMux I__1638 (
            .O(N__11200),
            .I(N__11194));
    LocalMux I__1637 (
            .O(N__11197),
            .I(r_Tx_Data_4_adj_960));
    LocalMux I__1636 (
            .O(N__11194),
            .I(r_Tx_Data_4_adj_960));
    InMux I__1635 (
            .O(N__11189),
            .I(N__11186));
    LocalMux I__1634 (
            .O(N__11186),
            .I(\c0.n4597 ));
    InMux I__1633 (
            .O(N__11183),
            .I(N__11179));
    CascadeMux I__1632 (
            .O(N__11182),
            .I(N__11176));
    LocalMux I__1631 (
            .O(N__11179),
            .I(N__11173));
    InMux I__1630 (
            .O(N__11176),
            .I(N__11169));
    Span4Mux_h I__1629 (
            .O(N__11173),
            .I(N__11166));
    InMux I__1628 (
            .O(N__11172),
            .I(N__11163));
    LocalMux I__1627 (
            .O(N__11169),
            .I(\c0.data_in_field_20 ));
    Odrv4 I__1626 (
            .O(N__11166),
            .I(\c0.data_in_field_20 ));
    LocalMux I__1625 (
            .O(N__11163),
            .I(\c0.data_in_field_20 ));
    InMux I__1624 (
            .O(N__11156),
            .I(N__11153));
    LocalMux I__1623 (
            .O(N__11153),
            .I(\c0.n4550 ));
    InMux I__1622 (
            .O(N__11150),
            .I(N__11147));
    LocalMux I__1621 (
            .O(N__11147),
            .I(\c0.tx2.n23 ));
    CascadeMux I__1620 (
            .O(N__11144),
            .I(n865_cascade_));
    InMux I__1619 (
            .O(N__11141),
            .I(N__11138));
    LocalMux I__1618 (
            .O(N__11138),
            .I(\c0.n4543 ));
    InMux I__1617 (
            .O(N__11135),
            .I(N__11129));
    InMux I__1616 (
            .O(N__11134),
            .I(N__11129));
    LocalMux I__1615 (
            .O(N__11129),
            .I(N__11126));
    Span4Mux_h I__1614 (
            .O(N__11126),
            .I(N__11122));
    InMux I__1613 (
            .O(N__11125),
            .I(N__11119));
    Odrv4 I__1612 (
            .O(N__11122),
            .I(blink_counter_22));
    LocalMux I__1611 (
            .O(N__11119),
            .I(blink_counter_22));
    InMux I__1610 (
            .O(N__11114),
            .I(N__11108));
    InMux I__1609 (
            .O(N__11113),
            .I(N__11108));
    LocalMux I__1608 (
            .O(N__11108),
            .I(N__11105));
    Span4Mux_v I__1607 (
            .O(N__11105),
            .I(N__11101));
    InMux I__1606 (
            .O(N__11104),
            .I(N__11098));
    Odrv4 I__1605 (
            .O(N__11101),
            .I(blink_counter_24));
    LocalMux I__1604 (
            .O(N__11098),
            .I(blink_counter_24));
    CascadeMux I__1603 (
            .O(N__11093),
            .I(N__11090));
    InMux I__1602 (
            .O(N__11090),
            .I(N__11084));
    InMux I__1601 (
            .O(N__11089),
            .I(N__11084));
    LocalMux I__1600 (
            .O(N__11084),
            .I(N__11081));
    Span4Mux_h I__1599 (
            .O(N__11081),
            .I(N__11077));
    InMux I__1598 (
            .O(N__11080),
            .I(N__11074));
    Odrv4 I__1597 (
            .O(N__11077),
            .I(blink_counter_21));
    LocalMux I__1596 (
            .O(N__11074),
            .I(blink_counter_21));
    CascadeMux I__1595 (
            .O(N__11069),
            .I(N__11065));
    InMux I__1594 (
            .O(N__11068),
            .I(N__11060));
    InMux I__1593 (
            .O(N__11065),
            .I(N__11060));
    LocalMux I__1592 (
            .O(N__11060),
            .I(N__11057));
    Span4Mux_h I__1591 (
            .O(N__11057),
            .I(N__11053));
    InMux I__1590 (
            .O(N__11056),
            .I(N__11050));
    Odrv4 I__1589 (
            .O(N__11053),
            .I(blink_counter_23));
    LocalMux I__1588 (
            .O(N__11050),
            .I(blink_counter_23));
    InMux I__1587 (
            .O(N__11045),
            .I(N__11042));
    LocalMux I__1586 (
            .O(N__11042),
            .I(N__11039));
    Span4Mux_h I__1585 (
            .O(N__11039),
            .I(N__11036));
    Span4Mux_v I__1584 (
            .O(N__11036),
            .I(N__11033));
    Odrv4 I__1583 (
            .O(N__11033),
            .I(\c0.n4580 ));
    InMux I__1582 (
            .O(N__11030),
            .I(N__11027));
    LocalMux I__1581 (
            .O(N__11027),
            .I(N__11024));
    Span4Mux_v I__1580 (
            .O(N__11024),
            .I(N__11021));
    Odrv4 I__1579 (
            .O(N__11021),
            .I(\c0.n4571 ));
    CascadeMux I__1578 (
            .O(N__11018),
            .I(\c0.n4855_cascade_ ));
    CascadeMux I__1577 (
            .O(N__11015),
            .I(tx2_data_0_keep_cascade_));
    InMux I__1576 (
            .O(N__11012),
            .I(N__11008));
    InMux I__1575 (
            .O(N__11011),
            .I(N__11005));
    LocalMux I__1574 (
            .O(N__11008),
            .I(r_Tx_Data_0_adj_964));
    LocalMux I__1573 (
            .O(N__11005),
            .I(r_Tx_Data_0_adj_964));
    InMux I__1572 (
            .O(N__11000),
            .I(N__10996));
    CascadeMux I__1571 (
            .O(N__10999),
            .I(N__10993));
    LocalMux I__1570 (
            .O(N__10996),
            .I(N__10990));
    InMux I__1569 (
            .O(N__10993),
            .I(N__10984));
    Span4Mux_v I__1568 (
            .O(N__10990),
            .I(N__10981));
    InMux I__1567 (
            .O(N__10989),
            .I(N__10976));
    InMux I__1566 (
            .O(N__10988),
            .I(N__10976));
    InMux I__1565 (
            .O(N__10987),
            .I(N__10973));
    LocalMux I__1564 (
            .O(N__10984),
            .I(\c0.data_in_field_32 ));
    Odrv4 I__1563 (
            .O(N__10981),
            .I(\c0.data_in_field_32 ));
    LocalMux I__1562 (
            .O(N__10976),
            .I(\c0.data_in_field_32 ));
    LocalMux I__1561 (
            .O(N__10973),
            .I(\c0.data_in_field_32 ));
    InMux I__1560 (
            .O(N__10964),
            .I(N__10961));
    LocalMux I__1559 (
            .O(N__10961),
            .I(\c0.n4579 ));
    InMux I__1558 (
            .O(N__10958),
            .I(N__10955));
    LocalMux I__1557 (
            .O(N__10955),
            .I(n1707));
    InMux I__1556 (
            .O(N__10952),
            .I(N__10949));
    LocalMux I__1555 (
            .O(N__10949),
            .I(n1768));
    InMux I__1554 (
            .O(N__10946),
            .I(N__10942));
    InMux I__1553 (
            .O(N__10945),
            .I(N__10939));
    LocalMux I__1552 (
            .O(N__10942),
            .I(\c0.tx2.r_Clock_Count_0 ));
    LocalMux I__1551 (
            .O(N__10939),
            .I(\c0.tx2.r_Clock_Count_0 ));
    InMux I__1550 (
            .O(N__10934),
            .I(N__10929));
    InMux I__1549 (
            .O(N__10933),
            .I(N__10926));
    InMux I__1548 (
            .O(N__10932),
            .I(N__10923));
    LocalMux I__1547 (
            .O(N__10929),
            .I(\c0.tx2.r_Clock_Count_2 ));
    LocalMux I__1546 (
            .O(N__10926),
            .I(\c0.tx2.r_Clock_Count_2 ));
    LocalMux I__1545 (
            .O(N__10923),
            .I(\c0.tx2.r_Clock_Count_2 ));
    InMux I__1544 (
            .O(N__10916),
            .I(N__10911));
    InMux I__1543 (
            .O(N__10915),
            .I(N__10908));
    InMux I__1542 (
            .O(N__10914),
            .I(N__10905));
    LocalMux I__1541 (
            .O(N__10911),
            .I(\c0.tx2.r_Clock_Count_5 ));
    LocalMux I__1540 (
            .O(N__10908),
            .I(\c0.tx2.r_Clock_Count_5 ));
    LocalMux I__1539 (
            .O(N__10905),
            .I(\c0.tx2.r_Clock_Count_5 ));
    CascadeMux I__1538 (
            .O(N__10898),
            .I(N__10893));
    InMux I__1537 (
            .O(N__10897),
            .I(N__10890));
    InMux I__1536 (
            .O(N__10896),
            .I(N__10887));
    InMux I__1535 (
            .O(N__10893),
            .I(N__10884));
    LocalMux I__1534 (
            .O(N__10890),
            .I(\c0.tx2.r_Clock_Count_1 ));
    LocalMux I__1533 (
            .O(N__10887),
            .I(\c0.tx2.r_Clock_Count_1 ));
    LocalMux I__1532 (
            .O(N__10884),
            .I(\c0.tx2.r_Clock_Count_1 ));
    InMux I__1531 (
            .O(N__10877),
            .I(N__10872));
    InMux I__1530 (
            .O(N__10876),
            .I(N__10869));
    InMux I__1529 (
            .O(N__10875),
            .I(N__10866));
    LocalMux I__1528 (
            .O(N__10872),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__1527 (
            .O(N__10869),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__1526 (
            .O(N__10866),
            .I(\c0.tx2.r_Clock_Count_3 ));
    CascadeMux I__1525 (
            .O(N__10859),
            .I(\c0.tx2.n5_cascade_ ));
    InMux I__1524 (
            .O(N__10856),
            .I(N__10853));
    LocalMux I__1523 (
            .O(N__10853),
            .I(n1701));
    InMux I__1522 (
            .O(N__10850),
            .I(N__10845));
    InMux I__1521 (
            .O(N__10849),
            .I(N__10842));
    InMux I__1520 (
            .O(N__10848),
            .I(N__10839));
    LocalMux I__1519 (
            .O(N__10845),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__1518 (
            .O(N__10842),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__1517 (
            .O(N__10839),
            .I(\c0.tx2.r_Clock_Count_4 ));
    CascadeMux I__1516 (
            .O(N__10832),
            .I(N__10829));
    InMux I__1515 (
            .O(N__10829),
            .I(N__10826));
    LocalMux I__1514 (
            .O(N__10826),
            .I(n1692));
    InMux I__1513 (
            .O(N__10823),
            .I(N__10818));
    InMux I__1512 (
            .O(N__10822),
            .I(N__10815));
    InMux I__1511 (
            .O(N__10821),
            .I(N__10812));
    LocalMux I__1510 (
            .O(N__10818),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1509 (
            .O(N__10815),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1508 (
            .O(N__10812),
            .I(\c0.tx2.r_Clock_Count_7 ));
    CascadeMux I__1507 (
            .O(N__10805),
            .I(r_SM_Main_2_N_759_1_cascade_));
    InMux I__1506 (
            .O(N__10802),
            .I(N__10794));
    InMux I__1505 (
            .O(N__10801),
            .I(N__10791));
    InMux I__1504 (
            .O(N__10800),
            .I(N__10788));
    InMux I__1503 (
            .O(N__10799),
            .I(N__10785));
    InMux I__1502 (
            .O(N__10798),
            .I(N__10780));
    InMux I__1501 (
            .O(N__10797),
            .I(N__10780));
    LocalMux I__1500 (
            .O(N__10794),
            .I(\c0.tx2.r_Clock_Count_8 ));
    LocalMux I__1499 (
            .O(N__10791),
            .I(\c0.tx2.r_Clock_Count_8 ));
    LocalMux I__1498 (
            .O(N__10788),
            .I(\c0.tx2.r_Clock_Count_8 ));
    LocalMux I__1497 (
            .O(N__10785),
            .I(\c0.tx2.r_Clock_Count_8 ));
    LocalMux I__1496 (
            .O(N__10780),
            .I(\c0.tx2.r_Clock_Count_8 ));
    InMux I__1495 (
            .O(N__10769),
            .I(N__10763));
    InMux I__1494 (
            .O(N__10768),
            .I(N__10760));
    InMux I__1493 (
            .O(N__10767),
            .I(N__10755));
    InMux I__1492 (
            .O(N__10766),
            .I(N__10755));
    LocalMux I__1491 (
            .O(N__10763),
            .I(\c0.tx2.n2902 ));
    LocalMux I__1490 (
            .O(N__10760),
            .I(\c0.tx2.n2902 ));
    LocalMux I__1489 (
            .O(N__10755),
            .I(\c0.tx2.n2902 ));
    InMux I__1488 (
            .O(N__10748),
            .I(N__10745));
    LocalMux I__1487 (
            .O(N__10745),
            .I(n4_adj_965));
    InMux I__1486 (
            .O(N__10742),
            .I(\c0.tx2.n3892 ));
    InMux I__1485 (
            .O(N__10739),
            .I(\c0.tx2.n3893 ));
    InMux I__1484 (
            .O(N__10736),
            .I(\c0.tx2.n3894 ));
    InMux I__1483 (
            .O(N__10733),
            .I(N__10730));
    LocalMux I__1482 (
            .O(N__10730),
            .I(n1698));
    InMux I__1481 (
            .O(N__10727),
            .I(\c0.tx2.n3895 ));
    InMux I__1480 (
            .O(N__10724),
            .I(\c0.tx2.n3896 ));
    InMux I__1479 (
            .O(N__10721),
            .I(\c0.tx2.n3897 ));
    InMux I__1478 (
            .O(N__10718),
            .I(bfn_4_22_0_));
    InMux I__1477 (
            .O(N__10715),
            .I(N__10712));
    LocalMux I__1476 (
            .O(N__10712),
            .I(n1689));
    InMux I__1475 (
            .O(N__10709),
            .I(N__10706));
    LocalMux I__1474 (
            .O(N__10706),
            .I(N__10703));
    Odrv4 I__1473 (
            .O(N__10703),
            .I(n1704));
    CascadeMux I__1472 (
            .O(N__10700),
            .I(N__10696));
    InMux I__1471 (
            .O(N__10699),
            .I(N__10693));
    InMux I__1470 (
            .O(N__10696),
            .I(N__10690));
    LocalMux I__1469 (
            .O(N__10693),
            .I(rx_data_3));
    LocalMux I__1468 (
            .O(N__10690),
            .I(rx_data_3));
    InMux I__1467 (
            .O(N__10685),
            .I(N__10681));
    InMux I__1466 (
            .O(N__10684),
            .I(N__10677));
    LocalMux I__1465 (
            .O(N__10681),
            .I(N__10674));
    InMux I__1464 (
            .O(N__10680),
            .I(N__10671));
    LocalMux I__1463 (
            .O(N__10677),
            .I(data_in_0_1));
    Odrv4 I__1462 (
            .O(N__10674),
            .I(data_in_0_1));
    LocalMux I__1461 (
            .O(N__10671),
            .I(data_in_0_1));
    CascadeMux I__1460 (
            .O(N__10664),
            .I(N__10661));
    InMux I__1459 (
            .O(N__10661),
            .I(N__10658));
    LocalMux I__1458 (
            .O(N__10658),
            .I(N__10655));
    Span4Mux_s2_h I__1457 (
            .O(N__10655),
            .I(N__10650));
    InMux I__1456 (
            .O(N__10654),
            .I(N__10645));
    InMux I__1455 (
            .O(N__10653),
            .I(N__10645));
    Odrv4 I__1454 (
            .O(N__10650),
            .I(data_in_5_5));
    LocalMux I__1453 (
            .O(N__10645),
            .I(data_in_5_5));
    InMux I__1452 (
            .O(N__10640),
            .I(N__10637));
    LocalMux I__1451 (
            .O(N__10637),
            .I(N__10633));
    InMux I__1450 (
            .O(N__10636),
            .I(N__10630));
    Span4Mux_v I__1449 (
            .O(N__10633),
            .I(N__10625));
    LocalMux I__1448 (
            .O(N__10630),
            .I(N__10625));
    Span4Mux_v I__1447 (
            .O(N__10625),
            .I(N__10622));
    Span4Mux_s1_h I__1446 (
            .O(N__10622),
            .I(N__10618));
    InMux I__1445 (
            .O(N__10621),
            .I(N__10615));
    Odrv4 I__1444 (
            .O(N__10618),
            .I(data_in_4_5));
    LocalMux I__1443 (
            .O(N__10615),
            .I(data_in_4_5));
    CascadeMux I__1442 (
            .O(N__10610),
            .I(\c0.rx.n4873_cascade_ ));
    InMux I__1441 (
            .O(N__10607),
            .I(N__10604));
    LocalMux I__1440 (
            .O(N__10604),
            .I(N__10599));
    InMux I__1439 (
            .O(N__10603),
            .I(N__10595));
    InMux I__1438 (
            .O(N__10602),
            .I(N__10592));
    Span4Mux_s3_h I__1437 (
            .O(N__10599),
            .I(N__10589));
    InMux I__1436 (
            .O(N__10598),
            .I(N__10586));
    LocalMux I__1435 (
            .O(N__10595),
            .I(data_in_3_7));
    LocalMux I__1434 (
            .O(N__10592),
            .I(data_in_3_7));
    Odrv4 I__1433 (
            .O(N__10589),
            .I(data_in_3_7));
    LocalMux I__1432 (
            .O(N__10586),
            .I(data_in_3_7));
    InMux I__1431 (
            .O(N__10577),
            .I(N__10574));
    LocalMux I__1430 (
            .O(N__10574),
            .I(N__10569));
    InMux I__1429 (
            .O(N__10573),
            .I(N__10566));
    InMux I__1428 (
            .O(N__10572),
            .I(N__10563));
    Odrv4 I__1427 (
            .O(N__10569),
            .I(data_in_4_1));
    LocalMux I__1426 (
            .O(N__10566),
            .I(data_in_4_1));
    LocalMux I__1425 (
            .O(N__10563),
            .I(data_in_4_1));
    InMux I__1424 (
            .O(N__10556),
            .I(N__10553));
    LocalMux I__1423 (
            .O(N__10553),
            .I(N__10549));
    InMux I__1422 (
            .O(N__10552),
            .I(N__10546));
    Span4Mux_v I__1421 (
            .O(N__10549),
            .I(N__10542));
    LocalMux I__1420 (
            .O(N__10546),
            .I(N__10539));
    InMux I__1419 (
            .O(N__10545),
            .I(N__10535));
    Span4Mux_s0_h I__1418 (
            .O(N__10542),
            .I(N__10532));
    Span4Mux_v I__1417 (
            .O(N__10539),
            .I(N__10529));
    InMux I__1416 (
            .O(N__10538),
            .I(N__10526));
    LocalMux I__1415 (
            .O(N__10535),
            .I(data_in_3_1));
    Odrv4 I__1414 (
            .O(N__10532),
            .I(data_in_3_1));
    Odrv4 I__1413 (
            .O(N__10529),
            .I(data_in_3_1));
    LocalMux I__1412 (
            .O(N__10526),
            .I(data_in_3_1));
    InMux I__1411 (
            .O(N__10517),
            .I(bfn_4_21_0_));
    InMux I__1410 (
            .O(N__10514),
            .I(N__10511));
    LocalMux I__1409 (
            .O(N__10511),
            .I(n1710));
    InMux I__1408 (
            .O(N__10508),
            .I(\c0.tx2.n3891 ));
    InMux I__1407 (
            .O(N__10505),
            .I(N__10500));
    InMux I__1406 (
            .O(N__10504),
            .I(N__10496));
    InMux I__1405 (
            .O(N__10503),
            .I(N__10493));
    LocalMux I__1404 (
            .O(N__10500),
            .I(N__10490));
    InMux I__1403 (
            .O(N__10499),
            .I(N__10487));
    LocalMux I__1402 (
            .O(N__10496),
            .I(data_in_2_1));
    LocalMux I__1401 (
            .O(N__10493),
            .I(data_in_2_1));
    Odrv4 I__1400 (
            .O(N__10490),
            .I(data_in_2_1));
    LocalMux I__1399 (
            .O(N__10487),
            .I(data_in_2_1));
    InMux I__1398 (
            .O(N__10478),
            .I(N__10475));
    LocalMux I__1397 (
            .O(N__10475),
            .I(N__10471));
    InMux I__1396 (
            .O(N__10474),
            .I(N__10467));
    Span4Mux_v I__1395 (
            .O(N__10471),
            .I(N__10464));
    InMux I__1394 (
            .O(N__10470),
            .I(N__10461));
    LocalMux I__1393 (
            .O(N__10467),
            .I(\c0.data_in_field_17 ));
    Odrv4 I__1392 (
            .O(N__10464),
            .I(\c0.data_in_field_17 ));
    LocalMux I__1391 (
            .O(N__10461),
            .I(\c0.data_in_field_17 ));
    InMux I__1390 (
            .O(N__10454),
            .I(N__10451));
    LocalMux I__1389 (
            .O(N__10451),
            .I(N__10447));
    InMux I__1388 (
            .O(N__10450),
            .I(N__10442));
    Span4Mux_h I__1387 (
            .O(N__10447),
            .I(N__10439));
    InMux I__1386 (
            .O(N__10446),
            .I(N__10436));
    InMux I__1385 (
            .O(N__10445),
            .I(N__10433));
    LocalMux I__1384 (
            .O(N__10442),
            .I(\c0.data_in_field_15 ));
    Odrv4 I__1383 (
            .O(N__10439),
            .I(\c0.data_in_field_15 ));
    LocalMux I__1382 (
            .O(N__10436),
            .I(\c0.data_in_field_15 ));
    LocalMux I__1381 (
            .O(N__10433),
            .I(\c0.data_in_field_15 ));
    CascadeMux I__1380 (
            .O(N__10424),
            .I(N__10419));
    InMux I__1379 (
            .O(N__10423),
            .I(N__10416));
    CascadeMux I__1378 (
            .O(N__10422),
            .I(N__10413));
    InMux I__1377 (
            .O(N__10419),
            .I(N__10410));
    LocalMux I__1376 (
            .O(N__10416),
            .I(N__10407));
    InMux I__1375 (
            .O(N__10413),
            .I(N__10404));
    LocalMux I__1374 (
            .O(N__10410),
            .I(\c0.data_in_field_27 ));
    Odrv4 I__1373 (
            .O(N__10407),
            .I(\c0.data_in_field_27 ));
    LocalMux I__1372 (
            .O(N__10404),
            .I(\c0.data_in_field_27 ));
    CascadeMux I__1371 (
            .O(N__10397),
            .I(N__10394));
    InMux I__1370 (
            .O(N__10394),
            .I(N__10391));
    LocalMux I__1369 (
            .O(N__10391),
            .I(N__10388));
    Span4Mux_s3_h I__1368 (
            .O(N__10388),
            .I(N__10385));
    Odrv4 I__1367 (
            .O(N__10385),
            .I(\c0.n4547 ));
    InMux I__1366 (
            .O(N__10382),
            .I(N__10379));
    LocalMux I__1365 (
            .O(N__10379),
            .I(N__10376));
    Span4Mux_h I__1364 (
            .O(N__10376),
            .I(N__10371));
    InMux I__1363 (
            .O(N__10375),
            .I(N__10368));
    InMux I__1362 (
            .O(N__10374),
            .I(N__10365));
    Odrv4 I__1361 (
            .O(N__10371),
            .I(data_in_0_3));
    LocalMux I__1360 (
            .O(N__10368),
            .I(data_in_0_3));
    LocalMux I__1359 (
            .O(N__10365),
            .I(data_in_0_3));
    InMux I__1358 (
            .O(N__10358),
            .I(N__10354));
    InMux I__1357 (
            .O(N__10357),
            .I(N__10351));
    LocalMux I__1356 (
            .O(N__10354),
            .I(N__10346));
    LocalMux I__1355 (
            .O(N__10351),
            .I(N__10346));
    Odrv4 I__1354 (
            .O(N__10346),
            .I(\c0.data_in_frame_7_5 ));
    InMux I__1353 (
            .O(N__10343),
            .I(N__10338));
    InMux I__1352 (
            .O(N__10342),
            .I(N__10335));
    InMux I__1351 (
            .O(N__10341),
            .I(N__10332));
    LocalMux I__1350 (
            .O(N__10338),
            .I(N__10323));
    LocalMux I__1349 (
            .O(N__10335),
            .I(N__10323));
    LocalMux I__1348 (
            .O(N__10332),
            .I(N__10323));
    InMux I__1347 (
            .O(N__10331),
            .I(N__10318));
    InMux I__1346 (
            .O(N__10330),
            .I(N__10318));
    Odrv12 I__1345 (
            .O(N__10323),
            .I(\c0.data_in_field_34 ));
    LocalMux I__1344 (
            .O(N__10318),
            .I(\c0.data_in_field_34 ));
    InMux I__1343 (
            .O(N__10313),
            .I(N__10310));
    LocalMux I__1342 (
            .O(N__10310),
            .I(N__10306));
    InMux I__1341 (
            .O(N__10309),
            .I(N__10303));
    Span4Mux_v I__1340 (
            .O(N__10306),
            .I(N__10296));
    LocalMux I__1339 (
            .O(N__10303),
            .I(N__10296));
    InMux I__1338 (
            .O(N__10302),
            .I(N__10290));
    InMux I__1337 (
            .O(N__10301),
            .I(N__10290));
    Span4Mux_v I__1336 (
            .O(N__10296),
            .I(N__10287));
    InMux I__1335 (
            .O(N__10295),
            .I(N__10284));
    LocalMux I__1334 (
            .O(N__10290),
            .I(\c0.data_in_field_3 ));
    Odrv4 I__1333 (
            .O(N__10287),
            .I(\c0.data_in_field_3 ));
    LocalMux I__1332 (
            .O(N__10284),
            .I(\c0.data_in_field_3 ));
    CascadeMux I__1331 (
            .O(N__10277),
            .I(N__10272));
    InMux I__1330 (
            .O(N__10276),
            .I(N__10267));
    InMux I__1329 (
            .O(N__10275),
            .I(N__10267));
    InMux I__1328 (
            .O(N__10272),
            .I(N__10263));
    LocalMux I__1327 (
            .O(N__10267),
            .I(N__10260));
    InMux I__1326 (
            .O(N__10266),
            .I(N__10257));
    LocalMux I__1325 (
            .O(N__10263),
            .I(\c0.data_in_field_19 ));
    Odrv12 I__1324 (
            .O(N__10260),
            .I(\c0.data_in_field_19 ));
    LocalMux I__1323 (
            .O(N__10257),
            .I(\c0.data_in_field_19 ));
    InMux I__1322 (
            .O(N__10250),
            .I(N__10247));
    LocalMux I__1321 (
            .O(N__10247),
            .I(N__10244));
    Odrv12 I__1320 (
            .O(N__10244),
            .I(\c0.n10 ));
    CascadeMux I__1319 (
            .O(N__10241),
            .I(N__10237));
    InMux I__1318 (
            .O(N__10240),
            .I(N__10234));
    InMux I__1317 (
            .O(N__10237),
            .I(N__10229));
    LocalMux I__1316 (
            .O(N__10234),
            .I(N__10226));
    InMux I__1315 (
            .O(N__10233),
            .I(N__10223));
    InMux I__1314 (
            .O(N__10232),
            .I(N__10220));
    LocalMux I__1313 (
            .O(N__10229),
            .I(\c0.data_in_field_29 ));
    Odrv12 I__1312 (
            .O(N__10226),
            .I(\c0.data_in_field_29 ));
    LocalMux I__1311 (
            .O(N__10223),
            .I(\c0.data_in_field_29 ));
    LocalMux I__1310 (
            .O(N__10220),
            .I(\c0.data_in_field_29 ));
    InMux I__1309 (
            .O(N__10211),
            .I(N__10208));
    LocalMux I__1308 (
            .O(N__10208),
            .I(\c0.n4411 ));
    CascadeMux I__1307 (
            .O(N__10205),
            .I(\c0.n4411_cascade_ ));
    CascadeMux I__1306 (
            .O(N__10202),
            .I(N__10199));
    InMux I__1305 (
            .O(N__10199),
            .I(N__10193));
    InMux I__1304 (
            .O(N__10198),
            .I(N__10193));
    LocalMux I__1303 (
            .O(N__10193),
            .I(\c0.data_in_frame_6_5 ));
    InMux I__1302 (
            .O(N__10190),
            .I(N__10187));
    LocalMux I__1301 (
            .O(N__10187),
            .I(N__10184));
    Span4Mux_s3_h I__1300 (
            .O(N__10184),
            .I(N__10181));
    Odrv4 I__1299 (
            .O(N__10181),
            .I(\c0.n4595 ));
    CascadeMux I__1298 (
            .O(N__10178),
            .I(\c0.n1340_cascade_ ));
    InMux I__1297 (
            .O(N__10175),
            .I(N__10170));
    InMux I__1296 (
            .O(N__10174),
            .I(N__10167));
    InMux I__1295 (
            .O(N__10173),
            .I(N__10164));
    LocalMux I__1294 (
            .O(N__10170),
            .I(N__10160));
    LocalMux I__1293 (
            .O(N__10167),
            .I(N__10155));
    LocalMux I__1292 (
            .O(N__10164),
            .I(N__10155));
    InMux I__1291 (
            .O(N__10163),
            .I(N__10151));
    Span4Mux_v I__1290 (
            .O(N__10160),
            .I(N__10148));
    Span4Mux_v I__1289 (
            .O(N__10155),
            .I(N__10145));
    InMux I__1288 (
            .O(N__10154),
            .I(N__10142));
    LocalMux I__1287 (
            .O(N__10151),
            .I(\c0.data_in_field_16 ));
    Odrv4 I__1286 (
            .O(N__10148),
            .I(\c0.data_in_field_16 ));
    Odrv4 I__1285 (
            .O(N__10145),
            .I(\c0.data_in_field_16 ));
    LocalMux I__1284 (
            .O(N__10142),
            .I(\c0.data_in_field_16 ));
    CascadeMux I__1283 (
            .O(N__10133),
            .I(N__10127));
    InMux I__1282 (
            .O(N__10132),
            .I(N__10124));
    InMux I__1281 (
            .O(N__10131),
            .I(N__10121));
    CascadeMux I__1280 (
            .O(N__10130),
            .I(N__10116));
    InMux I__1279 (
            .O(N__10127),
            .I(N__10113));
    LocalMux I__1278 (
            .O(N__10124),
            .I(N__10108));
    LocalMux I__1277 (
            .O(N__10121),
            .I(N__10108));
    InMux I__1276 (
            .O(N__10120),
            .I(N__10105));
    InMux I__1275 (
            .O(N__10119),
            .I(N__10100));
    InMux I__1274 (
            .O(N__10116),
            .I(N__10100));
    LocalMux I__1273 (
            .O(N__10113),
            .I(\c0.data_in_field_33 ));
    Odrv4 I__1272 (
            .O(N__10108),
            .I(\c0.data_in_field_33 ));
    LocalMux I__1271 (
            .O(N__10105),
            .I(\c0.data_in_field_33 ));
    LocalMux I__1270 (
            .O(N__10100),
            .I(\c0.data_in_field_33 ));
    InMux I__1269 (
            .O(N__10091),
            .I(N__10088));
    LocalMux I__1268 (
            .O(N__10088),
            .I(N__10082));
    InMux I__1267 (
            .O(N__10087),
            .I(N__10079));
    InMux I__1266 (
            .O(N__10086),
            .I(N__10076));
    InMux I__1265 (
            .O(N__10085),
            .I(N__10073));
    Span4Mux_h I__1264 (
            .O(N__10082),
            .I(N__10066));
    LocalMux I__1263 (
            .O(N__10079),
            .I(N__10066));
    LocalMux I__1262 (
            .O(N__10076),
            .I(N__10066));
    LocalMux I__1261 (
            .O(N__10073),
            .I(data_in_2_2));
    Odrv4 I__1260 (
            .O(N__10066),
            .I(data_in_2_2));
    InMux I__1259 (
            .O(N__10061),
            .I(N__10057));
    InMux I__1258 (
            .O(N__10060),
            .I(N__10054));
    LocalMux I__1257 (
            .O(N__10057),
            .I(N__10049));
    LocalMux I__1256 (
            .O(N__10054),
            .I(N__10046));
    InMux I__1255 (
            .O(N__10053),
            .I(N__10041));
    InMux I__1254 (
            .O(N__10052),
            .I(N__10041));
    Odrv12 I__1253 (
            .O(N__10049),
            .I(\c0.data_in_field_18 ));
    Odrv4 I__1252 (
            .O(N__10046),
            .I(\c0.data_in_field_18 ));
    LocalMux I__1251 (
            .O(N__10041),
            .I(\c0.data_in_field_18 ));
    CascadeMux I__1250 (
            .O(N__10034),
            .I(\c0.n4429_cascade_ ));
    InMux I__1249 (
            .O(N__10031),
            .I(N__10028));
    LocalMux I__1248 (
            .O(N__10028),
            .I(\c0.n4429 ));
    CascadeMux I__1247 (
            .O(N__10025),
            .I(N__10022));
    InMux I__1246 (
            .O(N__10022),
            .I(N__10015));
    InMux I__1245 (
            .O(N__10021),
            .I(N__10012));
    InMux I__1244 (
            .O(N__10020),
            .I(N__10009));
    InMux I__1243 (
            .O(N__10019),
            .I(N__10006));
    InMux I__1242 (
            .O(N__10018),
            .I(N__10003));
    LocalMux I__1241 (
            .O(N__10015),
            .I(\c0.data_in_field_46 ));
    LocalMux I__1240 (
            .O(N__10012),
            .I(\c0.data_in_field_46 ));
    LocalMux I__1239 (
            .O(N__10009),
            .I(\c0.data_in_field_46 ));
    LocalMux I__1238 (
            .O(N__10006),
            .I(\c0.data_in_field_46 ));
    LocalMux I__1237 (
            .O(N__10003),
            .I(\c0.data_in_field_46 ));
    CascadeMux I__1236 (
            .O(N__9992),
            .I(N__9989));
    InMux I__1235 (
            .O(N__9989),
            .I(N__9986));
    LocalMux I__1234 (
            .O(N__9986),
            .I(N__9983));
    Odrv4 I__1233 (
            .O(N__9983),
            .I(\c0.n6_adj_877 ));
    InMux I__1232 (
            .O(N__9980),
            .I(N__9974));
    InMux I__1231 (
            .O(N__9979),
            .I(N__9971));
    InMux I__1230 (
            .O(N__9978),
            .I(N__9968));
    InMux I__1229 (
            .O(N__9977),
            .I(N__9965));
    LocalMux I__1228 (
            .O(N__9974),
            .I(\c0.data_in_field_5 ));
    LocalMux I__1227 (
            .O(N__9971),
            .I(\c0.data_in_field_5 ));
    LocalMux I__1226 (
            .O(N__9968),
            .I(\c0.data_in_field_5 ));
    LocalMux I__1225 (
            .O(N__9965),
            .I(\c0.data_in_field_5 ));
    InMux I__1224 (
            .O(N__9956),
            .I(N__9953));
    LocalMux I__1223 (
            .O(N__9953),
            .I(\c0.n4450 ));
    InMux I__1222 (
            .O(N__9950),
            .I(N__9947));
    LocalMux I__1221 (
            .O(N__9947),
            .I(N__9944));
    Span4Mux_v I__1220 (
            .O(N__9944),
            .I(N__9939));
    InMux I__1219 (
            .O(N__9943),
            .I(N__9934));
    InMux I__1218 (
            .O(N__9942),
            .I(N__9934));
    Odrv4 I__1217 (
            .O(N__9939),
            .I(data_in_0_4));
    LocalMux I__1216 (
            .O(N__9934),
            .I(data_in_0_4));
    InMux I__1215 (
            .O(N__9929),
            .I(N__9925));
    InMux I__1214 (
            .O(N__9928),
            .I(N__9922));
    LocalMux I__1213 (
            .O(N__9925),
            .I(N__9914));
    LocalMux I__1212 (
            .O(N__9922),
            .I(N__9914));
    InMux I__1211 (
            .O(N__9921),
            .I(N__9909));
    InMux I__1210 (
            .O(N__9920),
            .I(N__9909));
    InMux I__1209 (
            .O(N__9919),
            .I(N__9906));
    Odrv4 I__1208 (
            .O(N__9914),
            .I(\c0.data_in_field_31 ));
    LocalMux I__1207 (
            .O(N__9909),
            .I(\c0.data_in_field_31 ));
    LocalMux I__1206 (
            .O(N__9906),
            .I(\c0.data_in_field_31 ));
    CascadeMux I__1205 (
            .O(N__9899),
            .I(\c0.n1261_cascade_ ));
    InMux I__1204 (
            .O(N__9896),
            .I(N__9891));
    InMux I__1203 (
            .O(N__9895),
            .I(N__9888));
    InMux I__1202 (
            .O(N__9894),
            .I(N__9884));
    LocalMux I__1201 (
            .O(N__9891),
            .I(N__9881));
    LocalMux I__1200 (
            .O(N__9888),
            .I(N__9878));
    InMux I__1199 (
            .O(N__9887),
            .I(N__9875));
    LocalMux I__1198 (
            .O(N__9884),
            .I(\c0.data_in_field_6 ));
    Odrv12 I__1197 (
            .O(N__9881),
            .I(\c0.data_in_field_6 ));
    Odrv4 I__1196 (
            .O(N__9878),
            .I(\c0.data_in_field_6 ));
    LocalMux I__1195 (
            .O(N__9875),
            .I(\c0.data_in_field_6 ));
    InMux I__1194 (
            .O(N__9866),
            .I(N__9862));
    InMux I__1193 (
            .O(N__9865),
            .I(N__9859));
    LocalMux I__1192 (
            .O(N__9862),
            .I(\c0.n1284 ));
    LocalMux I__1191 (
            .O(N__9859),
            .I(\c0.n1284 ));
    CascadeMux I__1190 (
            .O(N__9854),
            .I(\c0.n4408_cascade_ ));
    InMux I__1189 (
            .O(N__9851),
            .I(N__9847));
    InMux I__1188 (
            .O(N__9850),
            .I(N__9844));
    LocalMux I__1187 (
            .O(N__9847),
            .I(\c0.n4468 ));
    LocalMux I__1186 (
            .O(N__9844),
            .I(\c0.n4468 ));
    InMux I__1185 (
            .O(N__9839),
            .I(N__9836));
    LocalMux I__1184 (
            .O(N__9836),
            .I(N__9833));
    Span4Mux_h I__1183 (
            .O(N__9833),
            .I(N__9830));
    Span4Mux_v I__1182 (
            .O(N__9830),
            .I(N__9824));
    InMux I__1181 (
            .O(N__9829),
            .I(N__9819));
    InMux I__1180 (
            .O(N__9828),
            .I(N__9819));
    InMux I__1179 (
            .O(N__9827),
            .I(N__9816));
    Odrv4 I__1178 (
            .O(N__9824),
            .I(data_in_2_3));
    LocalMux I__1177 (
            .O(N__9819),
            .I(data_in_2_3));
    LocalMux I__1176 (
            .O(N__9816),
            .I(data_in_2_3));
    CascadeMux I__1175 (
            .O(N__9809),
            .I(N__9805));
    InMux I__1174 (
            .O(N__9808),
            .I(N__9802));
    InMux I__1173 (
            .O(N__9805),
            .I(N__9797));
    LocalMux I__1172 (
            .O(N__9802),
            .I(N__9794));
    InMux I__1171 (
            .O(N__9801),
            .I(N__9789));
    InMux I__1170 (
            .O(N__9800),
            .I(N__9789));
    LocalMux I__1169 (
            .O(N__9797),
            .I(N__9786));
    Span4Mux_h I__1168 (
            .O(N__9794),
            .I(N__9783));
    LocalMux I__1167 (
            .O(N__9789),
            .I(data_in_3_2));
    Odrv4 I__1166 (
            .O(N__9786),
            .I(data_in_3_2));
    Odrv4 I__1165 (
            .O(N__9783),
            .I(data_in_3_2));
    InMux I__1164 (
            .O(N__9776),
            .I(N__9773));
    LocalMux I__1163 (
            .O(N__9773),
            .I(N__9768));
    InMux I__1162 (
            .O(N__9772),
            .I(N__9765));
    CascadeMux I__1161 (
            .O(N__9771),
            .I(N__9761));
    Span4Mux_h I__1160 (
            .O(N__9768),
            .I(N__9756));
    LocalMux I__1159 (
            .O(N__9765),
            .I(N__9756));
    InMux I__1158 (
            .O(N__9764),
            .I(N__9751));
    InMux I__1157 (
            .O(N__9761),
            .I(N__9751));
    Odrv4 I__1156 (
            .O(N__9756),
            .I(data_in_2_5));
    LocalMux I__1155 (
            .O(N__9751),
            .I(data_in_2_5));
    CascadeMux I__1154 (
            .O(N__9746),
            .I(\c0.n1271_cascade_ ));
    InMux I__1153 (
            .O(N__9743),
            .I(N__9738));
    InMux I__1152 (
            .O(N__9742),
            .I(N__9733));
    InMux I__1151 (
            .O(N__9741),
            .I(N__9733));
    LocalMux I__1150 (
            .O(N__9738),
            .I(\c0.data_in_field_22 ));
    LocalMux I__1149 (
            .O(N__9733),
            .I(\c0.data_in_field_22 ));
    InMux I__1148 (
            .O(N__9728),
            .I(N__9725));
    LocalMux I__1147 (
            .O(N__9725),
            .I(N__9722));
    Span4Mux_v I__1146 (
            .O(N__9722),
            .I(N__9719));
    Odrv4 I__1145 (
            .O(N__9719),
            .I(\c0.n4556 ));
    CascadeMux I__1144 (
            .O(N__9716),
            .I(\c0.n10_adj_874_cascade_ ));
    InMux I__1143 (
            .O(N__9713),
            .I(N__9710));
    LocalMux I__1142 (
            .O(N__9710),
            .I(N__9707));
    Odrv4 I__1141 (
            .O(N__9707),
            .I(\c0.n4567 ));
    InMux I__1140 (
            .O(N__9704),
            .I(N__9701));
    LocalMux I__1139 (
            .O(N__9701),
            .I(N__9698));
    Span4Mux_v I__1138 (
            .O(N__9698),
            .I(N__9693));
    CascadeMux I__1137 (
            .O(N__9697),
            .I(N__9690));
    InMux I__1136 (
            .O(N__9696),
            .I(N__9687));
    Span4Mux_h I__1135 (
            .O(N__9693),
            .I(N__9684));
    InMux I__1134 (
            .O(N__9690),
            .I(N__9681));
    LocalMux I__1133 (
            .O(N__9687),
            .I(data_in_0_7));
    Odrv4 I__1132 (
            .O(N__9684),
            .I(data_in_0_7));
    LocalMux I__1131 (
            .O(N__9681),
            .I(data_in_0_7));
    InMux I__1130 (
            .O(N__9674),
            .I(N__9671));
    LocalMux I__1129 (
            .O(N__9671),
            .I(\c0.n4541 ));
    InMux I__1128 (
            .O(N__9668),
            .I(N__9665));
    LocalMux I__1127 (
            .O(N__9665),
            .I(N__9662));
    Odrv12 I__1126 (
            .O(N__9662),
            .I(\c0.n4544 ));
    CascadeMux I__1125 (
            .O(N__9659),
            .I(n4512_cascade_));
    InMux I__1124 (
            .O(N__9656),
            .I(N__9653));
    LocalMux I__1123 (
            .O(N__9653),
            .I(N__9650));
    Span4Mux_v I__1122 (
            .O(N__9650),
            .I(N__9647));
    Odrv4 I__1121 (
            .O(N__9647),
            .I(\c0.n4546 ));
    InMux I__1120 (
            .O(N__9644),
            .I(N__9641));
    LocalMux I__1119 (
            .O(N__9641),
            .I(\c0.n4603 ));
    CascadeMux I__1118 (
            .O(N__9638),
            .I(N__9634));
    InMux I__1117 (
            .O(N__9637),
            .I(N__9626));
    InMux I__1116 (
            .O(N__9634),
            .I(N__9626));
    InMux I__1115 (
            .O(N__9633),
            .I(N__9626));
    LocalMux I__1114 (
            .O(N__9626),
            .I(n1611));
    CascadeMux I__1113 (
            .O(N__9623),
            .I(n2326_cascade_));
    InMux I__1112 (
            .O(N__9620),
            .I(N__9617));
    LocalMux I__1111 (
            .O(N__9617),
            .I(n4514));
    InMux I__1110 (
            .O(N__9614),
            .I(N__9605));
    InMux I__1109 (
            .O(N__9613),
            .I(N__9605));
    InMux I__1108 (
            .O(N__9612),
            .I(N__9605));
    LocalMux I__1107 (
            .O(N__9605),
            .I(n4512));
    InMux I__1106 (
            .O(N__9602),
            .I(N__9599));
    LocalMux I__1105 (
            .O(N__9599),
            .I(N__9596));
    Span4Mux_v I__1104 (
            .O(N__9596),
            .I(N__9593));
    Odrv4 I__1103 (
            .O(N__9593),
            .I(n4523));
    CascadeMux I__1102 (
            .O(N__9590),
            .I(n4522_cascade_));
    InMux I__1101 (
            .O(N__9587),
            .I(N__9584));
    LocalMux I__1100 (
            .O(N__9584),
            .I(n4777));
    InMux I__1099 (
            .O(N__9581),
            .I(N__9576));
    InMux I__1098 (
            .O(N__9580),
            .I(N__9569));
    InMux I__1097 (
            .O(N__9579),
            .I(N__9569));
    LocalMux I__1096 (
            .O(N__9576),
            .I(N__9566));
    InMux I__1095 (
            .O(N__9575),
            .I(N__9563));
    InMux I__1094 (
            .O(N__9574),
            .I(N__9560));
    LocalMux I__1093 (
            .O(N__9569),
            .I(r_Bit_Index_1));
    Odrv4 I__1092 (
            .O(N__9566),
            .I(r_Bit_Index_1));
    LocalMux I__1091 (
            .O(N__9563),
            .I(r_Bit_Index_1));
    LocalMux I__1090 (
            .O(N__9560),
            .I(r_Bit_Index_1));
    CascadeMux I__1089 (
            .O(N__9551),
            .I(N__9545));
    InMux I__1088 (
            .O(N__9550),
            .I(N__9539));
    CascadeMux I__1087 (
            .O(N__9549),
            .I(N__9536));
    InMux I__1086 (
            .O(N__9548),
            .I(N__9533));
    InMux I__1085 (
            .O(N__9545),
            .I(N__9528));
    InMux I__1084 (
            .O(N__9544),
            .I(N__9528));
    InMux I__1083 (
            .O(N__9543),
            .I(N__9523));
    InMux I__1082 (
            .O(N__9542),
            .I(N__9523));
    LocalMux I__1081 (
            .O(N__9539),
            .I(N__9520));
    InMux I__1080 (
            .O(N__9536),
            .I(N__9517));
    LocalMux I__1079 (
            .O(N__9533),
            .I(r_Bit_Index_0_adj_956));
    LocalMux I__1078 (
            .O(N__9528),
            .I(r_Bit_Index_0_adj_956));
    LocalMux I__1077 (
            .O(N__9523),
            .I(r_Bit_Index_0_adj_956));
    Odrv4 I__1076 (
            .O(N__9520),
            .I(r_Bit_Index_0_adj_956));
    LocalMux I__1075 (
            .O(N__9517),
            .I(r_Bit_Index_0_adj_956));
    InMux I__1074 (
            .O(N__9506),
            .I(N__9502));
    InMux I__1073 (
            .O(N__9505),
            .I(N__9495));
    LocalMux I__1072 (
            .O(N__9502),
            .I(N__9492));
    InMux I__1071 (
            .O(N__9501),
            .I(N__9485));
    InMux I__1070 (
            .O(N__9500),
            .I(N__9485));
    InMux I__1069 (
            .O(N__9499),
            .I(N__9480));
    InMux I__1068 (
            .O(N__9498),
            .I(N__9480));
    LocalMux I__1067 (
            .O(N__9495),
            .I(N__9475));
    Span4Mux_s2_h I__1066 (
            .O(N__9492),
            .I(N__9475));
    InMux I__1065 (
            .O(N__9491),
            .I(N__9470));
    InMux I__1064 (
            .O(N__9490),
            .I(N__9470));
    LocalMux I__1063 (
            .O(N__9485),
            .I(r_Bit_Index_2_adj_955));
    LocalMux I__1062 (
            .O(N__9480),
            .I(r_Bit_Index_2_adj_955));
    Odrv4 I__1061 (
            .O(N__9475),
            .I(r_Bit_Index_2_adj_955));
    LocalMux I__1060 (
            .O(N__9470),
            .I(r_Bit_Index_2_adj_955));
    InMux I__1059 (
            .O(N__9461),
            .I(N__9458));
    LocalMux I__1058 (
            .O(N__9458),
            .I(N__9455));
    Odrv4 I__1057 (
            .O(N__9455),
            .I(n11_adj_941));
    CascadeMux I__1056 (
            .O(N__9452),
            .I(n4638_cascade_));
    InMux I__1055 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__1054 (
            .O(N__9446),
            .I(tx2_done));
    InMux I__1053 (
            .O(N__9443),
            .I(N__9440));
    LocalMux I__1052 (
            .O(N__9440),
            .I(\c0.n4598 ));
    InMux I__1051 (
            .O(N__9437),
            .I(N__9434));
    LocalMux I__1050 (
            .O(N__9434),
            .I(\c0.n4807 ));
    CascadeMux I__1049 (
            .O(N__9431),
            .I(tx2_data_2_keep_cascade_));
    InMux I__1048 (
            .O(N__9428),
            .I(N__9424));
    InMux I__1047 (
            .O(N__9427),
            .I(N__9421));
    LocalMux I__1046 (
            .O(N__9424),
            .I(r_Tx_Data_2_adj_962));
    LocalMux I__1045 (
            .O(N__9421),
            .I(r_Tx_Data_2_adj_962));
    InMux I__1044 (
            .O(N__9416),
            .I(N__9413));
    LocalMux I__1043 (
            .O(N__9413),
            .I(n9_adj_939));
    InMux I__1042 (
            .O(N__9410),
            .I(N__9405));
    InMux I__1041 (
            .O(N__9409),
            .I(N__9401));
    InMux I__1040 (
            .O(N__9408),
            .I(N__9398));
    LocalMux I__1039 (
            .O(N__9405),
            .I(N__9395));
    InMux I__1038 (
            .O(N__9404),
            .I(N__9392));
    LocalMux I__1037 (
            .O(N__9401),
            .I(data_in_2_0));
    LocalMux I__1036 (
            .O(N__9398),
            .I(data_in_2_0));
    Odrv4 I__1035 (
            .O(N__9395),
            .I(data_in_2_0));
    LocalMux I__1034 (
            .O(N__9392),
            .I(data_in_2_0));
    InMux I__1033 (
            .O(N__9383),
            .I(N__9380));
    LocalMux I__1032 (
            .O(N__9380),
            .I(N__9377));
    Odrv4 I__1031 (
            .O(N__9377),
            .I(\c0.n27 ));
    InMux I__1030 (
            .O(N__9374),
            .I(N__9371));
    LocalMux I__1029 (
            .O(N__9371),
            .I(\c0.rx.r_Rx_Data_R ));
    InMux I__1028 (
            .O(N__9368),
            .I(N__9363));
    InMux I__1027 (
            .O(N__9367),
            .I(N__9360));
    CascadeMux I__1026 (
            .O(N__9366),
            .I(N__9356));
    LocalMux I__1025 (
            .O(N__9363),
            .I(N__9353));
    LocalMux I__1024 (
            .O(N__9360),
            .I(N__9350));
    InMux I__1023 (
            .O(N__9359),
            .I(N__9345));
    InMux I__1022 (
            .O(N__9356),
            .I(N__9345));
    Odrv4 I__1021 (
            .O(N__9353),
            .I(data_in_1_4));
    Odrv4 I__1020 (
            .O(N__9350),
            .I(data_in_1_4));
    LocalMux I__1019 (
            .O(N__9345),
            .I(data_in_1_4));
    CascadeMux I__1018 (
            .O(N__9338),
            .I(N__9333));
    CascadeMux I__1017 (
            .O(N__9337),
            .I(N__9329));
    InMux I__1016 (
            .O(N__9336),
            .I(N__9326));
    InMux I__1015 (
            .O(N__9333),
            .I(N__9323));
    InMux I__1014 (
            .O(N__9332),
            .I(N__9320));
    InMux I__1013 (
            .O(N__9329),
            .I(N__9317));
    LocalMux I__1012 (
            .O(N__9326),
            .I(N__9310));
    LocalMux I__1011 (
            .O(N__9323),
            .I(N__9310));
    LocalMux I__1010 (
            .O(N__9320),
            .I(N__9310));
    LocalMux I__1009 (
            .O(N__9317),
            .I(data_in_1_7));
    Odrv4 I__1008 (
            .O(N__9310),
            .I(data_in_1_7));
    CascadeMux I__1007 (
            .O(N__9305),
            .I(N__9301));
    InMux I__1006 (
            .O(N__9304),
            .I(N__9298));
    InMux I__1005 (
            .O(N__9301),
            .I(N__9295));
    LocalMux I__1004 (
            .O(N__9298),
            .I(\c0.data_in_frame_7_0 ));
    LocalMux I__1003 (
            .O(N__9295),
            .I(\c0.data_in_frame_7_0 ));
    CascadeMux I__1002 (
            .O(N__9290),
            .I(N__9286));
    InMux I__1001 (
            .O(N__9289),
            .I(N__9283));
    InMux I__1000 (
            .O(N__9286),
            .I(N__9280));
    LocalMux I__999 (
            .O(N__9283),
            .I(N__9277));
    LocalMux I__998 (
            .O(N__9280),
            .I(N__9274));
    Span4Mux_h I__997 (
            .O(N__9277),
            .I(N__9269));
    Span4Mux_v I__996 (
            .O(N__9274),
            .I(N__9266));
    InMux I__995 (
            .O(N__9273),
            .I(N__9261));
    InMux I__994 (
            .O(N__9272),
            .I(N__9261));
    Odrv4 I__993 (
            .O(N__9269),
            .I(data_in_2_6));
    Odrv4 I__992 (
            .O(N__9266),
            .I(data_in_2_6));
    LocalMux I__991 (
            .O(N__9261),
            .I(data_in_2_6));
    InMux I__990 (
            .O(N__9254),
            .I(N__9251));
    LocalMux I__989 (
            .O(N__9251),
            .I(N__9247));
    CascadeMux I__988 (
            .O(N__9250),
            .I(N__9244));
    Span4Mux_v I__987 (
            .O(N__9247),
            .I(N__9241));
    InMux I__986 (
            .O(N__9244),
            .I(N__9238));
    Odrv4 I__985 (
            .O(N__9241),
            .I(rx_data_2));
    LocalMux I__984 (
            .O(N__9238),
            .I(rx_data_2));
    InMux I__983 (
            .O(N__9233),
            .I(N__9230));
    LocalMux I__982 (
            .O(N__9230),
            .I(PIN_2_c));
    InMux I__981 (
            .O(N__9227),
            .I(N__9223));
    CascadeMux I__980 (
            .O(N__9226),
            .I(N__9220));
    LocalMux I__979 (
            .O(N__9223),
            .I(N__9215));
    InMux I__978 (
            .O(N__9220),
            .I(N__9212));
    InMux I__977 (
            .O(N__9219),
            .I(N__9209));
    InMux I__976 (
            .O(N__9218),
            .I(N__9206));
    Odrv4 I__975 (
            .O(N__9215),
            .I(data_in_1_6));
    LocalMux I__974 (
            .O(N__9212),
            .I(data_in_1_6));
    LocalMux I__973 (
            .O(N__9209),
            .I(data_in_1_6));
    LocalMux I__972 (
            .O(N__9206),
            .I(data_in_1_6));
    InMux I__971 (
            .O(N__9197),
            .I(N__9194));
    LocalMux I__970 (
            .O(N__9194),
            .I(N__9191));
    Odrv4 I__969 (
            .O(N__9191),
            .I(\c0.n26_adj_869 ));
    CascadeMux I__968 (
            .O(N__9188),
            .I(N__9185));
    InMux I__967 (
            .O(N__9185),
            .I(N__9182));
    LocalMux I__966 (
            .O(N__9182),
            .I(N__9177));
    InMux I__965 (
            .O(N__9181),
            .I(N__9174));
    InMux I__964 (
            .O(N__9180),
            .I(N__9171));
    Span4Mux_v I__963 (
            .O(N__9177),
            .I(N__9168));
    LocalMux I__962 (
            .O(N__9174),
            .I(data_in_0_0));
    LocalMux I__961 (
            .O(N__9171),
            .I(data_in_0_0));
    Odrv4 I__960 (
            .O(N__9168),
            .I(data_in_0_0));
    InMux I__959 (
            .O(N__9161),
            .I(N__9158));
    LocalMux I__958 (
            .O(N__9158),
            .I(\c0.n30 ));
    CascadeMux I__957 (
            .O(N__9155),
            .I(\c0.n25_adj_870_cascade_ ));
    InMux I__956 (
            .O(N__9152),
            .I(N__9149));
    LocalMux I__955 (
            .O(N__9149),
            .I(\c0.n3933 ));
    CascadeMux I__954 (
            .O(N__9146),
            .I(\c0.n1197_cascade_ ));
    InMux I__953 (
            .O(N__9143),
            .I(N__9139));
    InMux I__952 (
            .O(N__9142),
            .I(N__9136));
    LocalMux I__951 (
            .O(N__9139),
            .I(\c0.data_in_frame_6_0 ));
    LocalMux I__950 (
            .O(N__9136),
            .I(\c0.data_in_frame_6_0 ));
    InMux I__949 (
            .O(N__9131),
            .I(N__9125));
    InMux I__948 (
            .O(N__9130),
            .I(N__9122));
    InMux I__947 (
            .O(N__9129),
            .I(N__9119));
    InMux I__946 (
            .O(N__9128),
            .I(N__9116));
    LocalMux I__945 (
            .O(N__9125),
            .I(data_in_3_5));
    LocalMux I__944 (
            .O(N__9122),
            .I(data_in_3_5));
    LocalMux I__943 (
            .O(N__9119),
            .I(data_in_3_5));
    LocalMux I__942 (
            .O(N__9116),
            .I(data_in_3_5));
    InMux I__941 (
            .O(N__9107),
            .I(N__9104));
    LocalMux I__940 (
            .O(N__9104),
            .I(N__9100));
    InMux I__939 (
            .O(N__9103),
            .I(N__9096));
    Span4Mux_v I__938 (
            .O(N__9100),
            .I(N__9093));
    InMux I__937 (
            .O(N__9099),
            .I(N__9090));
    LocalMux I__936 (
            .O(N__9096),
            .I(data_in_0_6));
    Odrv4 I__935 (
            .O(N__9093),
            .I(data_in_0_6));
    LocalMux I__934 (
            .O(N__9090),
            .I(data_in_0_6));
    InMux I__933 (
            .O(N__9083),
            .I(N__9079));
    InMux I__932 (
            .O(N__9082),
            .I(N__9074));
    LocalMux I__931 (
            .O(N__9079),
            .I(N__9071));
    InMux I__930 (
            .O(N__9078),
            .I(N__9066));
    InMux I__929 (
            .O(N__9077),
            .I(N__9066));
    LocalMux I__928 (
            .O(N__9074),
            .I(N__9063));
    Odrv4 I__927 (
            .O(N__9071),
            .I(data_in_1_3));
    LocalMux I__926 (
            .O(N__9066),
            .I(data_in_1_3));
    Odrv4 I__925 (
            .O(N__9063),
            .I(data_in_1_3));
    InMux I__924 (
            .O(N__9056),
            .I(N__9051));
    InMux I__923 (
            .O(N__9055),
            .I(N__9048));
    InMux I__922 (
            .O(N__9054),
            .I(N__9045));
    LocalMux I__921 (
            .O(N__9051),
            .I(data_in_5_6));
    LocalMux I__920 (
            .O(N__9048),
            .I(data_in_5_6));
    LocalMux I__919 (
            .O(N__9045),
            .I(data_in_5_6));
    InMux I__918 (
            .O(N__9038),
            .I(N__9035));
    LocalMux I__917 (
            .O(N__9035),
            .I(\c0.n4594 ));
    InMux I__916 (
            .O(N__9032),
            .I(N__9029));
    LocalMux I__915 (
            .O(N__9029),
            .I(\c0.n4825 ));
    InMux I__914 (
            .O(N__9026),
            .I(N__9023));
    LocalMux I__913 (
            .O(N__9023),
            .I(\c0.n4813 ));
    CascadeMux I__912 (
            .O(N__9020),
            .I(tx2_data_3_keep_cascade_));
    InMux I__911 (
            .O(N__9017),
            .I(N__9013));
    InMux I__910 (
            .O(N__9016),
            .I(N__9010));
    LocalMux I__909 (
            .O(N__9013),
            .I(N__9007));
    LocalMux I__908 (
            .O(N__9010),
            .I(r_Tx_Data_3_adj_961));
    Odrv4 I__907 (
            .O(N__9007),
            .I(r_Tx_Data_3_adj_961));
    InMux I__906 (
            .O(N__9002),
            .I(N__8999));
    LocalMux I__905 (
            .O(N__8999),
            .I(\c0.n4600 ));
    InMux I__904 (
            .O(N__8996),
            .I(N__8993));
    LocalMux I__903 (
            .O(N__8993),
            .I(N__8990));
    Odrv4 I__902 (
            .O(N__8990),
            .I(\c0.n4552 ));
    CascadeMux I__901 (
            .O(N__8987),
            .I(\c0.n4553_cascade_ ));
    InMux I__900 (
            .O(N__8984),
            .I(N__8981));
    LocalMux I__899 (
            .O(N__8981),
            .I(tx2_data_5_keep));
    CascadeMux I__898 (
            .O(N__8978),
            .I(N__8974));
    InMux I__897 (
            .O(N__8977),
            .I(N__8970));
    InMux I__896 (
            .O(N__8974),
            .I(N__8967));
    InMux I__895 (
            .O(N__8973),
            .I(N__8964));
    LocalMux I__894 (
            .O(N__8970),
            .I(data_in_0_5));
    LocalMux I__893 (
            .O(N__8967),
            .I(data_in_0_5));
    LocalMux I__892 (
            .O(N__8964),
            .I(data_in_0_5));
    CascadeMux I__891 (
            .O(N__8957),
            .I(N__8953));
    InMux I__890 (
            .O(N__8956),
            .I(N__8949));
    InMux I__889 (
            .O(N__8953),
            .I(N__8946));
    InMux I__888 (
            .O(N__8952),
            .I(N__8942));
    LocalMux I__887 (
            .O(N__8949),
            .I(N__8937));
    LocalMux I__886 (
            .O(N__8946),
            .I(N__8937));
    InMux I__885 (
            .O(N__8945),
            .I(N__8934));
    LocalMux I__884 (
            .O(N__8942),
            .I(data_in_1_0));
    Odrv4 I__883 (
            .O(N__8937),
            .I(data_in_1_0));
    LocalMux I__882 (
            .O(N__8934),
            .I(data_in_1_0));
    InMux I__881 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__880 (
            .O(N__8924),
            .I(tx2_data_7_keep));
    InMux I__879 (
            .O(N__8921),
            .I(N__8915));
    InMux I__878 (
            .O(N__8920),
            .I(N__8915));
    LocalMux I__877 (
            .O(N__8915),
            .I(r_Tx_Data_5_adj_959));
    InMux I__876 (
            .O(N__8912),
            .I(N__8909));
    LocalMux I__875 (
            .O(N__8909),
            .I(n4624));
    CascadeMux I__874 (
            .O(N__8906),
            .I(\c0.n4801_cascade_ ));
    CascadeMux I__873 (
            .O(N__8903),
            .I(tx2_data_1_keep_cascade_));
    InMux I__872 (
            .O(N__8900),
            .I(N__8894));
    InMux I__871 (
            .O(N__8899),
            .I(N__8894));
    LocalMux I__870 (
            .O(N__8894),
            .I(r_Tx_Data_1_adj_963));
    InMux I__869 (
            .O(N__8891),
            .I(N__8885));
    InMux I__868 (
            .O(N__8890),
            .I(N__8885));
    LocalMux I__867 (
            .O(N__8885),
            .I(r_Tx_Data_7_adj_957));
    InMux I__866 (
            .O(N__8882),
            .I(N__8879));
    LocalMux I__865 (
            .O(N__8879),
            .I(n4625));
    InMux I__864 (
            .O(N__8876),
            .I(N__8873));
    LocalMux I__863 (
            .O(N__8873),
            .I(\c0.n4540 ));
    InMux I__862 (
            .O(N__8870),
            .I(N__8867));
    LocalMux I__861 (
            .O(N__8867),
            .I(\c0.n4606 ));
    InMux I__860 (
            .O(N__8864),
            .I(N__8861));
    LocalMux I__859 (
            .O(N__8861),
            .I(N__8858));
    Span4Mux_v I__858 (
            .O(N__8858),
            .I(N__8854));
    InMux I__857 (
            .O(N__8857),
            .I(N__8851));
    Span4Mux_v I__856 (
            .O(N__8854),
            .I(N__8848));
    LocalMux I__855 (
            .O(N__8851),
            .I(\c0.data_in_frame_6_4 ));
    Odrv4 I__854 (
            .O(N__8848),
            .I(\c0.data_in_frame_6_4 ));
    InMux I__853 (
            .O(N__8843),
            .I(N__8840));
    LocalMux I__852 (
            .O(N__8840),
            .I(N__8836));
    InMux I__851 (
            .O(N__8839),
            .I(N__8833));
    Span4Mux_h I__850 (
            .O(N__8836),
            .I(N__8830));
    LocalMux I__849 (
            .O(N__8833),
            .I(\c0.data_in_frame_7_2 ));
    Odrv4 I__848 (
            .O(N__8830),
            .I(\c0.data_in_frame_7_2 ));
    CascadeMux I__847 (
            .O(N__8825),
            .I(\c0.n4604_cascade_ ));
    InMux I__846 (
            .O(N__8822),
            .I(N__8818));
    InMux I__845 (
            .O(N__8821),
            .I(N__8815));
    LocalMux I__844 (
            .O(N__8818),
            .I(\c0.data_in_frame_6_7 ));
    LocalMux I__843 (
            .O(N__8815),
            .I(\c0.data_in_frame_6_7 ));
    InMux I__842 (
            .O(N__8810),
            .I(N__8807));
    LocalMux I__841 (
            .O(N__8807),
            .I(N__8804));
    Odrv4 I__840 (
            .O(N__8804),
            .I(\c0.n4583 ));
    CascadeMux I__839 (
            .O(N__8801),
            .I(N__8798));
    InMux I__838 (
            .O(N__8798),
            .I(N__8792));
    InMux I__837 (
            .O(N__8797),
            .I(N__8792));
    LocalMux I__836 (
            .O(N__8792),
            .I(N__8789));
    Odrv4 I__835 (
            .O(N__8789),
            .I(\c0.data_in_frame_7_7 ));
    InMux I__834 (
            .O(N__8786),
            .I(N__8782));
    InMux I__833 (
            .O(N__8785),
            .I(N__8779));
    LocalMux I__832 (
            .O(N__8782),
            .I(\c0.data_in_frame_7_4 ));
    LocalMux I__831 (
            .O(N__8779),
            .I(\c0.data_in_frame_7_4 ));
    InMux I__830 (
            .O(N__8774),
            .I(N__8771));
    LocalMux I__829 (
            .O(N__8771),
            .I(\c0.n4555 ));
    InMux I__828 (
            .O(N__8768),
            .I(N__8762));
    InMux I__827 (
            .O(N__8767),
            .I(N__8762));
    LocalMux I__826 (
            .O(N__8762),
            .I(\c0.data_in_frame_6_3 ));
    CascadeMux I__825 (
            .O(N__8759),
            .I(N__8755));
    InMux I__824 (
            .O(N__8758),
            .I(N__8752));
    InMux I__823 (
            .O(N__8755),
            .I(N__8749));
    LocalMux I__822 (
            .O(N__8752),
            .I(N__8746));
    LocalMux I__821 (
            .O(N__8749),
            .I(\c0.data_in_frame_7_6 ));
    Odrv12 I__820 (
            .O(N__8746),
            .I(\c0.data_in_frame_7_6 ));
    InMux I__819 (
            .O(N__8741),
            .I(N__8738));
    LocalMux I__818 (
            .O(N__8738),
            .I(N__8735));
    Span4Mux_v I__817 (
            .O(N__8735),
            .I(N__8732));
    Odrv4 I__816 (
            .O(N__8732),
            .I(\c0.n4831 ));
    CascadeMux I__815 (
            .O(N__8729),
            .I(tx2_data_6_keep_cascade_));
    InMux I__814 (
            .O(N__8726),
            .I(N__8722));
    InMux I__813 (
            .O(N__8725),
            .I(N__8719));
    LocalMux I__812 (
            .O(N__8722),
            .I(r_Tx_Data_6_adj_958));
    LocalMux I__811 (
            .O(N__8719),
            .I(r_Tx_Data_6_adj_958));
    InMux I__810 (
            .O(N__8714),
            .I(N__8709));
    InMux I__809 (
            .O(N__8713),
            .I(N__8705));
    InMux I__808 (
            .O(N__8712),
            .I(N__8702));
    LocalMux I__807 (
            .O(N__8709),
            .I(N__8699));
    InMux I__806 (
            .O(N__8708),
            .I(N__8696));
    LocalMux I__805 (
            .O(N__8705),
            .I(data_in_1_5));
    LocalMux I__804 (
            .O(N__8702),
            .I(data_in_1_5));
    Odrv4 I__803 (
            .O(N__8699),
            .I(data_in_1_5));
    LocalMux I__802 (
            .O(N__8696),
            .I(data_in_1_5));
    InMux I__801 (
            .O(N__8687),
            .I(N__8684));
    LocalMux I__800 (
            .O(N__8684),
            .I(\c0.n28_adj_868 ));
    InMux I__799 (
            .O(N__8681),
            .I(N__8678));
    LocalMux I__798 (
            .O(N__8678),
            .I(\c0.n26 ));
    CascadeMux I__797 (
            .O(N__8675),
            .I(N__8672));
    InMux I__796 (
            .O(N__8672),
            .I(N__8666));
    InMux I__795 (
            .O(N__8671),
            .I(N__8666));
    LocalMux I__794 (
            .O(N__8666),
            .I(\c0.data_in_frame_7_3 ));
    InMux I__793 (
            .O(N__8663),
            .I(N__8660));
    LocalMux I__792 (
            .O(N__8660),
            .I(N__8657));
    Odrv4 I__791 (
            .O(N__8657),
            .I(\c0.n4601 ));
    InMux I__790 (
            .O(N__8654),
            .I(N__8648));
    InMux I__789 (
            .O(N__8653),
            .I(N__8648));
    LocalMux I__788 (
            .O(N__8648),
            .I(\c0.data_in_frame_6_6 ));
    InMux I__787 (
            .O(N__8645),
            .I(N__8642));
    LocalMux I__786 (
            .O(N__8642),
            .I(\c0.n4592 ));
    CascadeMux I__785 (
            .O(N__8639),
            .I(\c0.n25_cascade_ ));
    CascadeMux I__784 (
            .O(N__8636),
            .I(\c0.n4591_cascade_ ));
    CascadeMux I__783 (
            .O(N__8633),
            .I(\c0.n28_cascade_ ));
    InMux I__782 (
            .O(N__8630),
            .I(N__8627));
    LocalMux I__781 (
            .O(N__8627),
            .I(\c0.n22 ));
    CascadeMux I__780 (
            .O(N__8624),
            .I(\c0.n4849_cascade_ ));
    InMux I__779 (
            .O(N__8621),
            .I(N__8618));
    LocalMux I__778 (
            .O(N__8618),
            .I(\c0.n4568 ));
    InMux I__777 (
            .O(N__8615),
            .I(N__8612));
    LocalMux I__776 (
            .O(N__8612),
            .I(\c0.n4582 ));
    InMux I__775 (
            .O(N__8609),
            .I(N__8606));
    LocalMux I__774 (
            .O(N__8606),
            .I(n6));
    InMux I__773 (
            .O(N__8603),
            .I(n3870));
    InMux I__772 (
            .O(N__8600),
            .I(n3871));
    InMux I__771 (
            .O(N__8597),
            .I(n3872));
    InMux I__770 (
            .O(N__8594),
            .I(n3873));
    InMux I__769 (
            .O(N__8591),
            .I(bfn_1_25_0_));
    InMux I__768 (
            .O(N__8588),
            .I(n3875));
    InMux I__767 (
            .O(N__8585),
            .I(N__8582));
    LocalMux I__766 (
            .O(N__8582),
            .I(n14));
    InMux I__765 (
            .O(N__8579),
            .I(n3862));
    InMux I__764 (
            .O(N__8576),
            .I(N__8573));
    LocalMux I__763 (
            .O(N__8573),
            .I(n13));
    InMux I__762 (
            .O(N__8570),
            .I(n3863));
    InMux I__761 (
            .O(N__8567),
            .I(N__8564));
    LocalMux I__760 (
            .O(N__8564),
            .I(n12));
    InMux I__759 (
            .O(N__8561),
            .I(n3864));
    InMux I__758 (
            .O(N__8558),
            .I(N__8555));
    LocalMux I__757 (
            .O(N__8555),
            .I(n11));
    InMux I__756 (
            .O(N__8552),
            .I(n3865));
    InMux I__755 (
            .O(N__8549),
            .I(N__8546));
    LocalMux I__754 (
            .O(N__8546),
            .I(n10));
    InMux I__753 (
            .O(N__8543),
            .I(bfn_1_24_0_));
    InMux I__752 (
            .O(N__8540),
            .I(N__8537));
    LocalMux I__751 (
            .O(N__8537),
            .I(n9));
    InMux I__750 (
            .O(N__8534),
            .I(n3867));
    InMux I__749 (
            .O(N__8531),
            .I(N__8528));
    LocalMux I__748 (
            .O(N__8528),
            .I(n8));
    InMux I__747 (
            .O(N__8525),
            .I(n3868));
    InMux I__746 (
            .O(N__8522),
            .I(N__8519));
    LocalMux I__745 (
            .O(N__8519),
            .I(n7));
    InMux I__744 (
            .O(N__8516),
            .I(n3869));
    InMux I__743 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__742 (
            .O(N__8510),
            .I(n22));
    InMux I__741 (
            .O(N__8507),
            .I(n3854));
    InMux I__740 (
            .O(N__8504),
            .I(N__8501));
    LocalMux I__739 (
            .O(N__8501),
            .I(n21));
    InMux I__738 (
            .O(N__8498),
            .I(n3855));
    InMux I__737 (
            .O(N__8495),
            .I(N__8492));
    LocalMux I__736 (
            .O(N__8492),
            .I(n20));
    InMux I__735 (
            .O(N__8489),
            .I(n3856));
    InMux I__734 (
            .O(N__8486),
            .I(N__8483));
    LocalMux I__733 (
            .O(N__8483),
            .I(n19));
    InMux I__732 (
            .O(N__8480),
            .I(n3857));
    InMux I__731 (
            .O(N__8477),
            .I(N__8474));
    LocalMux I__730 (
            .O(N__8474),
            .I(n18));
    InMux I__729 (
            .O(N__8471),
            .I(bfn_1_23_0_));
    InMux I__728 (
            .O(N__8468),
            .I(N__8465));
    LocalMux I__727 (
            .O(N__8465),
            .I(n17));
    InMux I__726 (
            .O(N__8462),
            .I(n3859));
    InMux I__725 (
            .O(N__8459),
            .I(N__8456));
    LocalMux I__724 (
            .O(N__8456),
            .I(n16));
    InMux I__723 (
            .O(N__8453),
            .I(n3860));
    InMux I__722 (
            .O(N__8450),
            .I(N__8447));
    LocalMux I__721 (
            .O(N__8447),
            .I(n15));
    InMux I__720 (
            .O(N__8444),
            .I(n3861));
    IoInMux I__719 (
            .O(N__8441),
            .I(N__8438));
    LocalMux I__718 (
            .O(N__8438),
            .I(N__8435));
    IoSpan4Mux I__717 (
            .O(N__8435),
            .I(N__8432));
    IoSpan4Mux I__716 (
            .O(N__8432),
            .I(N__8429));
    IoSpan4Mux I__715 (
            .O(N__8429),
            .I(N__8426));
    Odrv4 I__714 (
            .O(N__8426),
            .I(CLK_pad_gb_input));
    InMux I__713 (
            .O(N__8423),
            .I(N__8420));
    LocalMux I__712 (
            .O(N__8420),
            .I(n26));
    InMux I__711 (
            .O(N__8417),
            .I(bfn_1_22_0_));
    InMux I__710 (
            .O(N__8414),
            .I(N__8411));
    LocalMux I__709 (
            .O(N__8411),
            .I(n25));
    InMux I__708 (
            .O(N__8408),
            .I(n3851));
    InMux I__707 (
            .O(N__8405),
            .I(N__8402));
    LocalMux I__706 (
            .O(N__8402),
            .I(n24));
    InMux I__705 (
            .O(N__8399),
            .I(n3852));
    InMux I__704 (
            .O(N__8396),
            .I(N__8393));
    LocalMux I__703 (
            .O(N__8393),
            .I(n23));
    InMux I__702 (
            .O(N__8390),
            .I(n3853));
    defparam IN_MUX_bfv_4_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_21_0_));
    defparam IN_MUX_bfv_4_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_22_0_ (
            .carryinitin(\c0.tx2.n3898 ),
            .carryinitout(bfn_4_22_0_));
    defparam IN_MUX_bfv_14_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_27_0_));
    defparam IN_MUX_bfv_14_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_28_0_ (
            .carryinitin(\c0.tx.n3883 ),
            .carryinitout(bfn_14_28_0_));
    defparam IN_MUX_bfv_5_32_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_32_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_32_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_6_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_25_0_));
    defparam IN_MUX_bfv_6_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_26_0_ (
            .carryinitin(\c0.n3913 ),
            .carryinitout(bfn_6_26_0_));
    defparam IN_MUX_bfv_5_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_24_0_));
    defparam IN_MUX_bfv_11_27_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_27_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(n3858),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(n3866),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(n3874),
            .carryinitout(bfn_1_25_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__8441),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam blink_counter_323__i0_LC_1_22_0.C_ON=1'b1;
    defparam blink_counter_323__i0_LC_1_22_0.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i0_LC_1_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i0_LC_1_22_0 (
            .in0(_gnd_net_),
            .in1(N__8423),
            .in2(_gnd_net_),
            .in3(N__8417),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(n3851),
            .clk(N__22866),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i1_LC_1_22_1.C_ON=1'b1;
    defparam blink_counter_323__i1_LC_1_22_1.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i1_LC_1_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i1_LC_1_22_1 (
            .in0(_gnd_net_),
            .in1(N__8414),
            .in2(_gnd_net_),
            .in3(N__8408),
            .lcout(n25),
            .ltout(),
            .carryin(n3851),
            .carryout(n3852),
            .clk(N__22866),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i2_LC_1_22_2.C_ON=1'b1;
    defparam blink_counter_323__i2_LC_1_22_2.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i2_LC_1_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i2_LC_1_22_2 (
            .in0(_gnd_net_),
            .in1(N__8405),
            .in2(_gnd_net_),
            .in3(N__8399),
            .lcout(n24),
            .ltout(),
            .carryin(n3852),
            .carryout(n3853),
            .clk(N__22866),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i3_LC_1_22_3.C_ON=1'b1;
    defparam blink_counter_323__i3_LC_1_22_3.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i3_LC_1_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i3_LC_1_22_3 (
            .in0(_gnd_net_),
            .in1(N__8396),
            .in2(_gnd_net_),
            .in3(N__8390),
            .lcout(n23),
            .ltout(),
            .carryin(n3853),
            .carryout(n3854),
            .clk(N__22866),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i4_LC_1_22_4.C_ON=1'b1;
    defparam blink_counter_323__i4_LC_1_22_4.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i4_LC_1_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i4_LC_1_22_4 (
            .in0(_gnd_net_),
            .in1(N__8513),
            .in2(_gnd_net_),
            .in3(N__8507),
            .lcout(n22),
            .ltout(),
            .carryin(n3854),
            .carryout(n3855),
            .clk(N__22866),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i5_LC_1_22_5.C_ON=1'b1;
    defparam blink_counter_323__i5_LC_1_22_5.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i5_LC_1_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i5_LC_1_22_5 (
            .in0(_gnd_net_),
            .in1(N__8504),
            .in2(_gnd_net_),
            .in3(N__8498),
            .lcout(n21),
            .ltout(),
            .carryin(n3855),
            .carryout(n3856),
            .clk(N__22866),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i6_LC_1_22_6.C_ON=1'b1;
    defparam blink_counter_323__i6_LC_1_22_6.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i6_LC_1_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i6_LC_1_22_6 (
            .in0(_gnd_net_),
            .in1(N__8495),
            .in2(_gnd_net_),
            .in3(N__8489),
            .lcout(n20),
            .ltout(),
            .carryin(n3856),
            .carryout(n3857),
            .clk(N__22866),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i7_LC_1_22_7.C_ON=1'b1;
    defparam blink_counter_323__i7_LC_1_22_7.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i7_LC_1_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i7_LC_1_22_7 (
            .in0(_gnd_net_),
            .in1(N__8486),
            .in2(_gnd_net_),
            .in3(N__8480),
            .lcout(n19),
            .ltout(),
            .carryin(n3857),
            .carryout(n3858),
            .clk(N__22866),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i8_LC_1_23_0.C_ON=1'b1;
    defparam blink_counter_323__i8_LC_1_23_0.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i8_LC_1_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i8_LC_1_23_0 (
            .in0(_gnd_net_),
            .in1(N__8477),
            .in2(_gnd_net_),
            .in3(N__8471),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(n3859),
            .clk(N__22867),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i9_LC_1_23_1.C_ON=1'b1;
    defparam blink_counter_323__i9_LC_1_23_1.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i9_LC_1_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i9_LC_1_23_1 (
            .in0(_gnd_net_),
            .in1(N__8468),
            .in2(_gnd_net_),
            .in3(N__8462),
            .lcout(n17),
            .ltout(),
            .carryin(n3859),
            .carryout(n3860),
            .clk(N__22867),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i10_LC_1_23_2.C_ON=1'b1;
    defparam blink_counter_323__i10_LC_1_23_2.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i10_LC_1_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i10_LC_1_23_2 (
            .in0(_gnd_net_),
            .in1(N__8459),
            .in2(_gnd_net_),
            .in3(N__8453),
            .lcout(n16),
            .ltout(),
            .carryin(n3860),
            .carryout(n3861),
            .clk(N__22867),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i11_LC_1_23_3.C_ON=1'b1;
    defparam blink_counter_323__i11_LC_1_23_3.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i11_LC_1_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i11_LC_1_23_3 (
            .in0(_gnd_net_),
            .in1(N__8450),
            .in2(_gnd_net_),
            .in3(N__8444),
            .lcout(n15),
            .ltout(),
            .carryin(n3861),
            .carryout(n3862),
            .clk(N__22867),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i12_LC_1_23_4.C_ON=1'b1;
    defparam blink_counter_323__i12_LC_1_23_4.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i12_LC_1_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i12_LC_1_23_4 (
            .in0(_gnd_net_),
            .in1(N__8585),
            .in2(_gnd_net_),
            .in3(N__8579),
            .lcout(n14),
            .ltout(),
            .carryin(n3862),
            .carryout(n3863),
            .clk(N__22867),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i13_LC_1_23_5.C_ON=1'b1;
    defparam blink_counter_323__i13_LC_1_23_5.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i13_LC_1_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i13_LC_1_23_5 (
            .in0(_gnd_net_),
            .in1(N__8576),
            .in2(_gnd_net_),
            .in3(N__8570),
            .lcout(n13),
            .ltout(),
            .carryin(n3863),
            .carryout(n3864),
            .clk(N__22867),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i14_LC_1_23_6.C_ON=1'b1;
    defparam blink_counter_323__i14_LC_1_23_6.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i14_LC_1_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i14_LC_1_23_6 (
            .in0(_gnd_net_),
            .in1(N__8567),
            .in2(_gnd_net_),
            .in3(N__8561),
            .lcout(n12),
            .ltout(),
            .carryin(n3864),
            .carryout(n3865),
            .clk(N__22867),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i15_LC_1_23_7.C_ON=1'b1;
    defparam blink_counter_323__i15_LC_1_23_7.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i15_LC_1_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i15_LC_1_23_7 (
            .in0(_gnd_net_),
            .in1(N__8558),
            .in2(_gnd_net_),
            .in3(N__8552),
            .lcout(n11),
            .ltout(),
            .carryin(n3865),
            .carryout(n3866),
            .clk(N__22867),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i16_LC_1_24_0.C_ON=1'b1;
    defparam blink_counter_323__i16_LC_1_24_0.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i16_LC_1_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i16_LC_1_24_0 (
            .in0(_gnd_net_),
            .in1(N__8549),
            .in2(_gnd_net_),
            .in3(N__8543),
            .lcout(n10),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(n3867),
            .clk(N__22868),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i17_LC_1_24_1.C_ON=1'b1;
    defparam blink_counter_323__i17_LC_1_24_1.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i17_LC_1_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i17_LC_1_24_1 (
            .in0(_gnd_net_),
            .in1(N__8540),
            .in2(_gnd_net_),
            .in3(N__8534),
            .lcout(n9),
            .ltout(),
            .carryin(n3867),
            .carryout(n3868),
            .clk(N__22868),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i18_LC_1_24_2.C_ON=1'b1;
    defparam blink_counter_323__i18_LC_1_24_2.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i18_LC_1_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i18_LC_1_24_2 (
            .in0(_gnd_net_),
            .in1(N__8531),
            .in2(_gnd_net_),
            .in3(N__8525),
            .lcout(n8),
            .ltout(),
            .carryin(n3868),
            .carryout(n3869),
            .clk(N__22868),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i19_LC_1_24_3.C_ON=1'b1;
    defparam blink_counter_323__i19_LC_1_24_3.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i19_LC_1_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i19_LC_1_24_3 (
            .in0(_gnd_net_),
            .in1(N__8522),
            .in2(_gnd_net_),
            .in3(N__8516),
            .lcout(n7),
            .ltout(),
            .carryin(n3869),
            .carryout(n3870),
            .clk(N__22868),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i20_LC_1_24_4.C_ON=1'b1;
    defparam blink_counter_323__i20_LC_1_24_4.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i20_LC_1_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i20_LC_1_24_4 (
            .in0(_gnd_net_),
            .in1(N__8609),
            .in2(_gnd_net_),
            .in3(N__8603),
            .lcout(n6),
            .ltout(),
            .carryin(n3870),
            .carryout(n3871),
            .clk(N__22868),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i21_LC_1_24_5.C_ON=1'b1;
    defparam blink_counter_323__i21_LC_1_24_5.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i21_LC_1_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i21_LC_1_24_5 (
            .in0(_gnd_net_),
            .in1(N__11080),
            .in2(_gnd_net_),
            .in3(N__8600),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n3871),
            .carryout(n3872),
            .clk(N__22868),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i22_LC_1_24_6.C_ON=1'b1;
    defparam blink_counter_323__i22_LC_1_24_6.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i22_LC_1_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i22_LC_1_24_6 (
            .in0(_gnd_net_),
            .in1(N__11125),
            .in2(_gnd_net_),
            .in3(N__8597),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n3872),
            .carryout(n3873),
            .clk(N__22868),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i23_LC_1_24_7.C_ON=1'b1;
    defparam blink_counter_323__i23_LC_1_24_7.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i23_LC_1_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i23_LC_1_24_7 (
            .in0(_gnd_net_),
            .in1(N__11056),
            .in2(_gnd_net_),
            .in3(N__8594),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n3873),
            .carryout(n3874),
            .clk(N__22868),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i24_LC_1_25_0.C_ON=1'b1;
    defparam blink_counter_323__i24_LC_1_25_0.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i24_LC_1_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i24_LC_1_25_0 (
            .in0(_gnd_net_),
            .in1(N__11104),
            .in2(_gnd_net_),
            .in3(N__8591),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_1_25_0_),
            .carryout(n3875),
            .clk(N__22871),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_323__i25_LC_1_25_1.C_ON=1'b0;
    defparam blink_counter_323__i25_LC_1_25_1.SEQ_MODE=4'b1000;
    defparam blink_counter_323__i25_LC_1_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_323__i25_LC_1_25_1 (
            .in0(_gnd_net_),
            .in1(N__12229),
            .in2(_gnd_net_),
            .in3(N__8588),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22871),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i55_LC_1_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i55_LC_1_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i55_LC_1_25_7 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i55_LC_1_25_7  (
            .in0(N__8822),
            .in1(N__15028),
            .in2(N__14589),
            .in3(N__13685),
            .lcout(\c0.data_in_frame_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22871),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i39_LC_1_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i39_LC_1_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i39_LC_1_26_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i39_LC_1_26_0  (
            .in0(N__17090),
            .in1(N__9055),
            .in2(_gnd_net_),
            .in3(N__11715),
            .lcout(data_in_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i31_LC_1_26_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i31_LC_1_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i31_LC_1_26_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i31_LC_1_26_1  (
            .in0(N__11716),
            .in1(N__17091),
            .in2(_gnd_net_),
            .in3(N__11834),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4483_LC_1_26_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4483_LC_1_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4483_LC_1_26_2 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_4483_LC_1_26_2  (
            .in0(N__8810),
            .in1(N__15638),
            .in2(N__15783),
            .in3(N__8615),
            .lcout(),
            .ltout(\c0.n4849_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4849_bdd_4_lut_LC_1_26_3 .C_ON=1'b0;
    defparam \c0.n4849_bdd_4_lut_LC_1_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.n4849_bdd_4_lut_LC_1_26_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n4849_bdd_4_lut_LC_1_26_3  (
            .in0(N__15761),
            .in1(N__9713),
            .in2(N__8624),
            .in3(N__8621),
            .lcout(tx2_data_7_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4213_3_lut_LC_1_26_5 .C_ON=1'b0;
    defparam \c0.i4213_3_lut_LC_1_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4213_3_lut_LC_1_26_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4213_3_lut_LC_1_26_5  (
            .in0(N__15517),
            .in1(N__9929),
            .in2(_gnd_net_),
            .in3(N__13376),
            .lcout(\c0.n4568 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4216_3_lut_LC_1_26_7 .C_ON=1'b0;
    defparam \c0.i4216_3_lut_LC_1_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4216_3_lut_LC_1_26_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4216_3_lut_LC_1_26_7  (
            .in0(N__15516),
            .in1(N__13763),
            .in2(_gnd_net_),
            .in3(N__10175),
            .lcout(\c0.n4571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i6_LC_1_27_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i6_LC_1_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i6_LC_1_27_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i6_LC_1_27_0  (
            .in0(N__8977),
            .in1(N__8714),
            .in2(_gnd_net_),
            .in3(N__17002),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22879),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i40_LC_1_27_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i40_LC_1_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i40_LC_1_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i40_LC_1_27_1  (
            .in0(N__17001),
            .in1(N__11514),
            .in2(_gnd_net_),
            .in3(N__11498),
            .lcout(data_in_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22879),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i27_LC_1_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i27_LC_1_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i27_LC_1_27_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i27_LC_1_27_3  (
            .in0(N__17000),
            .in1(N__11384),
            .in2(_gnd_net_),
            .in3(N__9801),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22879),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4227_3_lut_LC_1_27_4 .C_ON=1'b0;
    defparam \c0.i4227_3_lut_LC_1_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4227_3_lut_LC_1_27_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4227_3_lut_LC_1_27_4  (
            .in0(N__15560),
            .in1(N__12046),
            .in2(_gnd_net_),
            .in3(N__12876),
            .lcout(\c0.n4582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i19_LC_1_27_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i19_LC_1_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i19_LC_1_27_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i19_LC_1_27_5  (
            .in0(N__16999),
            .in1(N__9800),
            .in2(_gnd_net_),
            .in3(N__10085),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22879),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i58_LC_1_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i58_LC_1_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i58_LC_1_27_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i58_LC_1_27_6  (
            .in0(N__8839),
            .in1(N__15882),
            .in2(N__14715),
            .in3(N__14962),
            .lcout(\c0.data_in_frame_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22879),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i1_LC_1_28_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i1_LC_1_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i1_LC_1_28_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i1_LC_1_28_1  (
            .in0(N__17126),
            .in1(N__9180),
            .in2(_gnd_net_),
            .in3(N__8956),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22882),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4454_LC_1_28_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4454_LC_1_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4454_LC_1_28_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_4454_LC_1_28_2  (
            .in0(N__15646),
            .in1(N__8663),
            .in2(N__15788),
            .in3(N__9002),
            .lcout(\c0.n4813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i13_LC_1_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i13_LC_1_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i13_LC_1_28_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i13_LC_1_28_3  (
            .in0(N__8712),
            .in1(N__14961),
            .in2(N__14721),
            .in3(N__13146),
            .lcout(\c0.data_in_field_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22882),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4236_3_lut_LC_1_28_4 .C_ON=1'b0;
    defparam \c0.i4236_3_lut_LC_1_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4236_3_lut_LC_1_28_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4236_3_lut_LC_1_28_4  (
            .in0(N__15559),
            .in1(N__12008),
            .in2(_gnd_net_),
            .in3(N__10021),
            .lcout(),
            .ltout(\c0.n4591_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4478_LC_1_28_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4478_LC_1_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4478_LC_1_28_5 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_4478_LC_1_28_5  (
            .in0(N__15778),
            .in1(N__15647),
            .in2(N__8636),
            .in3(N__8645),
            .lcout(\c0.n4831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_LC_1_28_6 .C_ON=1'b0;
    defparam \c0.i6_2_lut_LC_1_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_LC_1_28_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i6_2_lut_LC_1_28_6  (
            .in0(_gnd_net_),
            .in1(N__8973),
            .in2(_gnd_net_),
            .in3(N__15078),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4197_3_lut_LC_1_28_7 .C_ON=1'b0;
    defparam \c0.i4197_3_lut_LC_1_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4197_3_lut_LC_1_28_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4197_3_lut_LC_1_28_7  (
            .in0(N__15558),
            .in1(N__9979),
            .in2(_gnd_net_),
            .in3(N__13145),
            .lcout(\c0.n4552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_1_29_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_1_29_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i12_4_lut_LC_1_29_0  (
            .in0(N__13784),
            .in1(N__9128),
            .in2(N__12143),
            .in3(N__9272),
            .lcout(),
            .ltout(\c0.n28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_1_29_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_1_29_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_LC_1_29_1  (
            .in0(N__10499),
            .in1(N__11838),
            .in2(N__8633),
            .in3(N__8630),
            .lcout(\c0.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i14_LC_1_29_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i14_LC_1_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i14_LC_1_29_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i14_LC_1_29_2  (
            .in0(N__8713),
            .in1(N__9772),
            .in2(_gnd_net_),
            .in3(N__17120),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22888),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i11_LC_1_29_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i11_LC_1_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i11_LC_1_29_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i11_LC_1_29_3  (
            .in0(N__17116),
            .in1(N__15071),
            .in2(_gnd_net_),
            .in3(N__10087),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22888),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i54_LC_1_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i54_LC_1_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i54_LC_1_29_4 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i54_LC_1_29_4  (
            .in0(N__8654),
            .in1(N__14946),
            .in2(N__14725),
            .in3(N__13939),
            .lcout(\c0.data_in_frame_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22888),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i23_LC_1_29_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i23_LC_1_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i23_LC_1_29_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i23_LC_1_29_5  (
            .in0(N__9273),
            .in1(_gnd_net_),
            .in2(N__17127),
            .in3(N__11839),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22888),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i41_LC_1_29_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i41_LC_1_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i41_LC_1_29_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i41_LC_1_29_6  (
            .in0(N__14707),
            .in1(N__14945),
            .in2(N__17468),
            .in3(N__13895),
            .lcout(\c0.data_in_field_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22888),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4237_3_lut_LC_1_29_7 .C_ON=1'b0;
    defparam \c0.i4237_3_lut_LC_1_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4237_3_lut_LC_1_29_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.i4237_3_lut_LC_1_29_7  (
            .in0(N__8758),
            .in1(N__8653),
            .in2(N__15546),
            .in3(_gnd_net_),
            .lcout(\c0.n4592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_1_30_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_1_30_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i9_4_lut_LC_1_30_0  (
            .in0(N__9082),
            .in1(N__10086),
            .in2(N__9366),
            .in3(N__8945),
            .lcout(),
            .ltout(\c0.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_1_30_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_1_30_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i15_4_lut_LC_1_30_1  (
            .in0(N__8687),
            .in1(N__8681),
            .in2(N__8639),
            .in3(N__9383),
            .lcout(\c0.n3933 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i9_LC_1_30_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i9_LC_1_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i9_LC_1_30_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i9_LC_1_30_2  (
            .in0(N__8952),
            .in1(N__16923),
            .in2(_gnd_net_),
            .in3(N__9410),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22893),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i30_LC_1_30_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i30_LC_1_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i30_LC_1_30_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i30_LC_1_30_3  (
            .in0(N__16920),
            .in1(N__10636),
            .in2(_gnd_net_),
            .in3(N__9129),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22893),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i18_LC_1_30_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i18_LC_1_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i18_LC_1_30_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i18_LC_1_30_4  (
            .in0(N__10556),
            .in1(N__16922),
            .in2(_gnd_net_),
            .in3(N__10503),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22893),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i13_LC_1_30_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i13_LC_1_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i13_LC_1_30_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i13_LC_1_30_5  (
            .in0(N__16919),
            .in1(N__12112),
            .in2(_gnd_net_),
            .in3(N__9359),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22893),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_291_LC_1_30_6 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_291_LC_1_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_291_LC_1_30_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i12_4_lut_adj_291_LC_1_30_6  (
            .in0(N__9332),
            .in1(N__9099),
            .in2(N__9697),
            .in3(N__8708),
            .lcout(\c0.n28_adj_868 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i7_LC_1_30_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i7_LC_1_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i7_LC_1_30_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_0___i7_LC_1_30_7  (
            .in0(N__16921),
            .in1(_gnd_net_),
            .in2(N__9226),
            .in3(N__9103),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22893),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_1_31_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_1_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_1_31_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10_4_lut_LC_1_31_0  (
            .in0(N__10374),
            .in1(N__9827),
            .in2(N__9771),
            .in3(N__9404),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i59_LC_1_31_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i59_LC_1_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i59_LC_1_31_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i59_LC_1_31_1  (
            .in0(N__14937),
            .in1(N__14716),
            .in2(N__8675),
            .in3(N__14118),
            .lcout(\c0.data_in_frame_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22899),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4225_3_lut_LC_1_31_2 .C_ON=1'b0;
    defparam \c0.i4225_3_lut_LC_1_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4225_3_lut_LC_1_31_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.i4225_3_lut_LC_1_31_2  (
            .in0(N__15547),
            .in1(_gnd_net_),
            .in2(N__9305),
            .in3(N__9142),
            .lcout(\c0.n4580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i63_LC_1_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i63_LC_1_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i63_LC_1_31_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i63_LC_1_31_3  (
            .in0(N__17020),
            .in1(N__12338),
            .in2(_gnd_net_),
            .in3(N__14084),
            .lcout(data_in_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22899),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i22_LC_1_31_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i22_LC_1_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i22_LC_1_31_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i22_LC_1_31_4  (
            .in0(N__9764),
            .in1(N__17021),
            .in2(_gnd_net_),
            .in3(N__9130),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22899),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4246_3_lut_LC_1_31_5 .C_ON=1'b0;
    defparam \c0.i4246_3_lut_LC_1_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4246_3_lut_LC_1_31_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4246_3_lut_LC_1_31_5  (
            .in0(N__8671),
            .in1(N__8767),
            .in2(_gnd_net_),
            .in3(N__15548),
            .lcout(\c0.n4601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i51_LC_1_31_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i51_LC_1_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i51_LC_1_31_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i51_LC_1_31_6  (
            .in0(N__8768),
            .in1(N__14939),
            .in2(N__14726),
            .in3(N__16595),
            .lcout(\c0.data_in_frame_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22899),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i62_LC_1_31_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i62_LC_1_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i62_LC_1_31_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i62_LC_1_31_7  (
            .in0(N__14938),
            .in1(N__14085),
            .in2(N__8759),
            .in3(N__14720),
            .lcout(\c0.data_in_frame_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22899),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i52_LC_1_32_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i52_LC_1_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i52_LC_1_32_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i52_LC_1_32_2  (
            .in0(N__8857),
            .in1(N__11984),
            .in2(N__14714),
            .in3(N__15046),
            .lcout(\c0.data_in_frame_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22907),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i12_LC_1_32_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i12_LC_1_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i12_LC_1_32_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i12_LC_1_32_3  (
            .in0(N__9829),
            .in1(N__17094),
            .in2(_gnd_net_),
            .in3(N__9077),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22907),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i20_LC_1_32_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i20_LC_1_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i20_LC_1_32_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i20_LC_1_32_4  (
            .in0(N__17093),
            .in1(N__14209),
            .in2(_gnd_net_),
            .in3(N__9828),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22907),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i4_LC_1_32_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i4_LC_1_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i4_LC_1_32_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i4_LC_1_32_5  (
            .in0(N__17095),
            .in1(N__10375),
            .in2(_gnd_net_),
            .in3(N__9078),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22907),
            .ce(),
            .sr(_gnd_net_));
    defparam i4168_3_lut_LC_2_22_1.C_ON=1'b0;
    defparam i4168_3_lut_LC_2_22_1.SEQ_MODE=4'b0000;
    defparam i4168_3_lut_LC_2_22_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 i4168_3_lut_LC_2_22_1 (
            .in0(N__8725),
            .in1(N__9427),
            .in2(_gnd_net_),
            .in3(N__9506),
            .lcout(n4523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_388_LC_2_22_3.C_ON=1'b0;
    defparam i1_2_lut_adj_388_LC_2_22_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_388_LC_2_22_3.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_388_LC_2_22_3 (
            .in0(_gnd_net_),
            .in1(N__12569),
            .in2(_gnd_net_),
            .in3(N__12640),
            .lcout(n11_adj_941),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4831_bdd_4_lut_LC_2_23_1 .C_ON=1'b0;
    defparam \c0.n4831_bdd_4_lut_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n4831_bdd_4_lut_LC_2_23_1 .LUT_INIT=16'b1111110000001010;
    LogicCell40 \c0.n4831_bdd_4_lut_LC_2_23_1  (
            .in0(N__8774),
            .in1(N__9728),
            .in2(N__15787),
            .in3(N__8741),
            .lcout(),
            .ltout(tx2_data_6_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i6_LC_2_23_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i6_LC_2_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i6_LC_2_23_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx2.r_Tx_Data_i6_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(N__11228),
            .in2(N__8729),
            .in3(N__8726),
            .lcout(r_Tx_Data_6_adj_958),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22869),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4243_3_lut_LC_2_23_5 .C_ON=1'b0;
    defparam \c0.i4243_3_lut_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4243_3_lut_LC_2_23_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4243_3_lut_LC_2_23_5  (
            .in0(N__8785),
            .in1(N__8864),
            .in2(_gnd_net_),
            .in3(N__15518),
            .lcout(\c0.n4598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4249_3_lut_LC_2_24_0 .C_ON=1'b0;
    defparam \c0.i4249_3_lut_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4249_3_lut_LC_2_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4249_3_lut_LC_2_24_0  (
            .in0(N__8843),
            .in1(N__12932),
            .in2(_gnd_net_),
            .in3(N__15467),
            .lcout(),
            .ltout(\c0.n4604_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4449_LC_2_24_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4449_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4449_LC_2_24_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_4449_LC_2_24_1  (
            .in0(N__15731),
            .in1(N__15635),
            .in2(N__8825),
            .in3(N__9644),
            .lcout(\c0.n4807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4228_3_lut_LC_2_24_2 .C_ON=1'b0;
    defparam \c0.i4228_3_lut_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4228_3_lut_LC_2_24_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.i4228_3_lut_LC_2_24_2  (
            .in0(N__8797),
            .in1(N__15466),
            .in2(_gnd_net_),
            .in3(N__8821),
            .lcout(\c0.n4583 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i63_LC_2_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i63_LC_2_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i63_LC_2_24_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i63_LC_2_24_4  (
            .in0(N__14963),
            .in1(N__14574),
            .in2(N__8801),
            .in3(N__13723),
            .lcout(\c0.data_in_frame_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22872),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i60_LC_2_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i60_LC_2_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i60_LC_2_24_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i60_LC_2_24_5  (
            .in0(N__8786),
            .in1(N__13835),
            .in2(N__14670),
            .in3(N__14964),
            .lcout(\c0.data_in_frame_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22872),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4200_3_lut_LC_2_24_6 .C_ON=1'b0;
    defparam \c0.i4200_3_lut_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4200_3_lut_LC_2_24_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4200_3_lut_LC_2_24_6  (
            .in0(N__15471),
            .in1(N__12790),
            .in2(_gnd_net_),
            .in3(N__9896),
            .lcout(\c0.n4555 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1384_2_lut_4_lut_LC_2_24_7 .C_ON=1'b0;
    defparam \c0.tx2.i1384_2_lut_4_lut_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1384_2_lut_4_lut_LC_2_24_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \c0.tx2.i1384_2_lut_4_lut_LC_2_24_7  (
            .in0(N__9550),
            .in1(N__9575),
            .in2(N__12572),
            .in3(N__9505),
            .lcout(n1611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_1__bdd_4_lut_LC_2_25_0.C_ON=1'b0;
    defparam r_Bit_Index_1__bdd_4_lut_LC_2_25_0.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_1__bdd_4_lut_LC_2_25_0.LUT_INIT=16'b1101101010001010;
    LogicCell40 r_Bit_Index_1__bdd_4_lut_LC_2_25_0 (
            .in0(N__9574),
            .in1(N__8882),
            .in2(N__9549),
            .in3(N__8912),
            .lcout(n4777),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i5_LC_2_25_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i5_LC_2_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i5_LC_2_25_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx2.r_Tx_Data_i5_LC_2_25_1  (
            .in0(N__11247),
            .in1(N__8984),
            .in2(_gnd_net_),
            .in3(N__8921),
            .lcout(r_Tx_Data_5_adj_959),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22876),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i7_LC_2_25_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i7_LC_2_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i7_LC_2_25_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx2.r_Tx_Data_i7_LC_2_25_2  (
            .in0(N__8891),
            .in1(N__11248),
            .in2(_gnd_net_),
            .in3(N__8927),
            .lcout(r_Tx_Data_7_adj_957),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22876),
            .ce(),
            .sr(_gnd_net_));
    defparam i4269_3_lut_LC_2_25_3.C_ON=1'b0;
    defparam i4269_3_lut_LC_2_25_3.SEQ_MODE=4'b0000;
    defparam i4269_3_lut_LC_2_25_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 i4269_3_lut_LC_2_25_3 (
            .in0(N__9490),
            .in1(N__8920),
            .in2(_gnd_net_),
            .in3(N__8899),
            .lcout(n4624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4444_LC_2_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4444_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4444_LC_2_25_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_4444_LC_2_25_4  (
            .in0(N__15639),
            .in1(N__8870),
            .in2(N__15784),
            .in3(N__11858),
            .lcout(),
            .ltout(\c0.n4801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4801_bdd_4_lut_LC_2_25_5 .C_ON=1'b0;
    defparam \c0.n4801_bdd_4_lut_LC_2_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.n4801_bdd_4_lut_LC_2_25_5 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n4801_bdd_4_lut_LC_2_25_5  (
            .in0(N__8876),
            .in1(N__15765),
            .in2(N__8906),
            .in3(N__9674),
            .lcout(),
            .ltout(tx2_data_1_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i1_LC_2_25_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i1_LC_2_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i1_LC_2_25_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.tx2.r_Tx_Data_i1_LC_2_25_6  (
            .in0(N__8900),
            .in1(_gnd_net_),
            .in2(N__8903),
            .in3(N__11246),
            .lcout(r_Tx_Data_1_adj_963),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22876),
            .ce(),
            .sr(_gnd_net_));
    defparam i4270_3_lut_LC_2_25_7.C_ON=1'b0;
    defparam i4270_3_lut_LC_2_25_7.SEQ_MODE=4'b0000;
    defparam i4270_3_lut_LC_2_25_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i4270_3_lut_LC_2_25_7 (
            .in0(N__9491),
            .in1(N__8890),
            .in2(_gnd_net_),
            .in3(N__9017),
            .lcout(n4625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4185_3_lut_LC_2_26_0 .C_ON=1'b0;
    defparam \c0.i4185_3_lut_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4185_3_lut_LC_2_26_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4185_3_lut_LC_2_26_0  (
            .in0(N__15512),
            .in1(N__12836),
            .in2(_gnd_net_),
            .in3(N__13496),
            .lcout(\c0.n4540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4251_3_lut_LC_2_26_1 .C_ON=1'b0;
    defparam \c0.i4251_3_lut_LC_2_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4251_3_lut_LC_2_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4251_3_lut_LC_2_26_1  (
            .in0(N__15525),
            .in1(N__13906),
            .in2(_gnd_net_),
            .in3(N__10132),
            .lcout(\c0.n4606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i22_LC_2_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i22_LC_2_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i22_LC_2_26_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i22_LC_2_26_2  (
            .in0(N__9742),
            .in1(N__14646),
            .in2(N__9290),
            .in3(N__15033),
            .lcout(\c0.data_in_field_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22880),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4239_3_lut_LC_2_26_3 .C_ON=1'b0;
    defparam \c0.i4239_3_lut_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4239_3_lut_LC_2_26_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.i4239_3_lut_LC_2_26_3  (
            .in0(N__13044),
            .in1(N__15511),
            .in2(_gnd_net_),
            .in3(N__13328),
            .lcout(\c0.n4594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4198_3_lut_LC_2_26_4 .C_ON=1'b0;
    defparam \c0.i4198_3_lut_LC_2_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4198_3_lut_LC_2_26_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.i4198_3_lut_LC_2_26_4  (
            .in0(N__11693),
            .in1(N__15526),
            .in2(_gnd_net_),
            .in3(N__10240),
            .lcout(),
            .ltout(\c0.n4553_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4825_bdd_4_lut_LC_2_26_5 .C_ON=1'b0;
    defparam \c0.n4825_bdd_4_lut_LC_2_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.n4825_bdd_4_lut_LC_2_26_5 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n4825_bdd_4_lut_LC_2_26_5  (
            .in0(N__15760),
            .in1(N__8996),
            .in2(N__8987),
            .in3(N__9032),
            .lcout(tx2_data_5_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_321_LC_2_26_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_321_LC_2_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_321_LC_2_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_321_LC_2_26_6  (
            .in0(N__10174),
            .in1(N__9928),
            .in2(N__15883),
            .in3(N__10019),
            .lcout(\c0.n10_adj_876 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_2_26_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_2_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_LC_2_26_7  (
            .in0(N__13597),
            .in1(N__9741),
            .in2(_gnd_net_),
            .in3(N__13327),
            .lcout(\c0.n1284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i5_LC_2_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i5_LC_2_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i5_LC_2_27_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i5_LC_2_27_0  (
            .in0(N__14958),
            .in1(N__14641),
            .in2(N__8978),
            .in3(N__9980),
            .lcout(\c0.data_in_field_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i59_LC_2_27_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i59_LC_2_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i59_LC_2_27_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i59_LC_2_27_1  (
            .in0(N__17129),
            .in1(N__9254),
            .in2(_gnd_net_),
            .in3(N__15878),
            .lcout(data_in_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i8_LC_2_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i8_LC_2_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i8_LC_2_27_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i8_LC_2_27_2  (
            .in0(N__14959),
            .in1(N__14644),
            .in2(N__8957),
            .in3(N__11596),
            .lcout(\c0.data_in_field_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i47_LC_2_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i47_LC_2_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i47_LC_2_27_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i47_LC_2_27_3  (
            .in0(N__17128),
            .in1(N__9054),
            .in2(_gnd_net_),
            .in3(N__13940),
            .lcout(data_in_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i46_LC_2_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i46_LC_2_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i46_LC_2_27_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i46_LC_2_27_4  (
            .in0(N__14957),
            .in1(N__9056),
            .in2(N__10025),
            .in3(N__14643),
            .lcout(\c0.data_in_field_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i36_LC_2_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i36_LC_2_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i36_LC_2_27_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i36_LC_2_27_5  (
            .in0(N__14645),
            .in1(N__14960),
            .in2(N__13612),
            .in3(N__11948),
            .lcout(\c0.data_in_field_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i37_LC_2_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i37_LC_2_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i37_LC_2_27_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i37_LC_2_27_6  (
            .in0(N__14956),
            .in1(N__10640),
            .in2(N__13342),
            .in3(N__14642),
            .lcout(\c0.data_in_field_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4464_LC_2_27_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4464_LC_2_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4464_LC_2_27_7 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_4464_LC_2_27_7  (
            .in0(N__10190),
            .in1(N__15640),
            .in2(N__15782),
            .in3(N__9038),
            .lcout(\c0.n4825 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4813_bdd_4_lut_LC_2_28_0 .C_ON=1'b0;
    defparam \c0.n4813_bdd_4_lut_LC_2_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.n4813_bdd_4_lut_LC_2_28_0 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \c0.n4813_bdd_4_lut_LC_2_28_0  (
            .in0(N__9656),
            .in1(N__15766),
            .in2(N__10397),
            .in3(N__9026),
            .lcout(),
            .ltout(tx2_data_3_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_28_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_28_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx2.r_Tx_Data_i3_LC_2_28_1  (
            .in0(_gnd_net_),
            .in1(N__11252),
            .in2(N__9020),
            .in3(N__9016),
            .lcout(r_Tx_Data_3_adj_961),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22889),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i20_LC_2_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i20_LC_2_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i20_LC_2_28_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i20_LC_2_28_2  (
            .in0(N__15021),
            .in1(N__12113),
            .in2(N__11182),
            .in3(N__14628),
            .lcout(\c0.data_in_field_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22889),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i35_LC_2_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i35_LC_2_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i35_LC_2_28_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i35_LC_2_28_3  (
            .in0(N__13644),
            .in1(N__14234),
            .in2(N__14702),
            .in3(N__15024),
            .lcout(\c0.data_in_field_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22889),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4245_3_lut_LC_2_28_4 .C_ON=1'b0;
    defparam \c0.i4245_3_lut_LC_2_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4245_3_lut_LC_2_28_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4245_3_lut_LC_2_28_4  (
            .in0(N__15520),
            .in1(N__13558),
            .in2(_gnd_net_),
            .in3(N__13643),
            .lcout(\c0.n4600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i6_LC_2_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i6_LC_2_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i6_LC_2_28_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i6_LC_2_28_5  (
            .in0(N__9107),
            .in1(N__15023),
            .in2(N__14703),
            .in3(N__9894),
            .lcout(\c0.data_in_field_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22889),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_296_LC_2_28_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_296_LC_2_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_296_LC_2_28_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_296_LC_2_28_6  (
            .in0(_gnd_net_),
            .in1(N__13886),
            .in2(_gnd_net_),
            .in3(N__11338),
            .lcout(\c0.n4450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i45_LC_2_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i45_LC_2_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i45_LC_2_28_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i45_LC_2_28_7  (
            .in0(N__14621),
            .in1(N__15022),
            .in2(N__10664),
            .in3(N__13031),
            .lcout(\c0.data_in_field_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22889),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_323_LC_2_29_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_323_LC_2_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_323_LC_2_29_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_323_LC_2_29_0  (
            .in0(_gnd_net_),
            .in1(N__14086),
            .in2(_gnd_net_),
            .in3(N__10988),
            .lcout(\c0.n6_adj_877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i33_LC_2_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i33_LC_2_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i33_LC_2_29_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i33_LC_2_29_1  (
            .in0(N__14629),
            .in1(N__14932),
            .in2(N__10133),
            .in3(N__10577),
            .lcout(\c0.data_in_field_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22894),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_38_2_lut_LC_2_29_2 .C_ON=1'b0;
    defparam \c0.i1_rep_38_2_lut_LC_2_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_38_2_lut_LC_2_29_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_rep_38_2_lut_LC_2_29_2  (
            .in0(_gnd_net_),
            .in1(N__10989),
            .in2(_gnd_net_),
            .in3(N__9920),
            .lcout(\c0.n4927 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i31_LC_2_29_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i31_LC_2_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i31_LC_2_29_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i31_LC_2_29_3  (
            .in0(N__9921),
            .in1(N__10607),
            .in2(N__14706),
            .in3(N__14933),
            .lcout(\c0.data_in_field_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22894),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i11_LC_2_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i11_LC_2_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i11_LC_2_29_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i11_LC_2_29_4  (
            .in0(N__14928),
            .in1(N__9083),
            .in2(N__11355),
            .in3(N__14639),
            .lcout(\c0.data_in_field_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22894),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i0_LC_2_29_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i0_LC_2_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i0_LC_2_29_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i0_LC_2_29_5  (
            .in0(N__9181),
            .in1(N__14930),
            .in2(N__14704),
            .in3(N__11631),
            .lcout(\c0.data_in_field_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22894),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i27_LC_2_29_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i27_LC_2_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i27_LC_2_29_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i27_LC_2_29_6  (
            .in0(N__14929),
            .in1(N__14210),
            .in2(N__10424),
            .in3(N__14640),
            .lcout(\c0.data_in_field_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22894),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i12_LC_2_29_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i12_LC_2_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i12_LC_2_29_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i12_LC_2_29_7  (
            .in0(N__9368),
            .in1(N__14931),
            .in2(N__14705),
            .in3(N__14012),
            .lcout(\c0.data_in_field_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22894),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_293_LC_2_30_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_293_LC_2_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_293_LC_2_30_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_293_LC_2_30_0  (
            .in0(N__12105),
            .in1(N__14202),
            .in2(N__9188),
            .in3(N__9808),
            .lcout(),
            .ltout(\c0.n25_adj_870_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_LC_2_30_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_LC_2_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_LC_2_30_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i1_4_lut_LC_2_30_1  (
            .in0(N__9161),
            .in1(N__9197),
            .in2(N__9155),
            .in3(N__9152),
            .lcout(\c0.n1197 ),
            .ltout(\c0.n1197_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i48_LC_2_30_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i48_LC_2_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i48_LC_2_30_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i48_LC_2_30_2  (
            .in0(N__14687),
            .in1(N__9143),
            .in2(N__9146),
            .in3(N__16088),
            .lcout(\c0.data_in_frame_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22900),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i8_LC_2_30_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i8_LC_2_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i8_LC_2_30_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i8_LC_2_30_3  (
            .in0(N__9336),
            .in1(N__9696),
            .in2(_gnd_net_),
            .in3(N__16918),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22900),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i15_LC_2_30_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i15_LC_2_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i15_LC_2_30_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i15_LC_2_30_4  (
            .in0(N__14686),
            .in1(N__14940),
            .in2(N__9338),
            .in3(N__10450),
            .lcout(\c0.data_in_field_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22900),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i14_LC_2_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i14_LC_2_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i14_LC_2_30_5 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i14_LC_2_30_5  (
            .in0(N__9227),
            .in1(N__12786),
            .in2(N__15025),
            .in3(N__14688),
            .lcout(\c0.data_in_field_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22900),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i25_LC_2_30_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i25_LC_2_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i25_LC_2_30_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i25_LC_2_30_6  (
            .in0(N__16917),
            .in1(N__14254),
            .in2(_gnd_net_),
            .in3(N__13785),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22900),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i29_LC_2_30_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i29_LC_2_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i29_LC_2_30_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i29_LC_2_30_7  (
            .in0(N__9131),
            .in1(N__14944),
            .in2(N__10241),
            .in3(N__14689),
            .lcout(\c0.data_in_field_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22900),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i60_LC_2_31_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i60_LC_2_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i60_LC_2_31_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i60_LC_2_31_0  (
            .in0(N__10699),
            .in1(_gnd_net_),
            .in2(N__17098),
            .in3(N__14114),
            .lcout(data_in_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i56_LC_2_31_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i56_LC_2_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i56_LC_2_31_1 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i56_LC_2_31_1  (
            .in0(N__15019),
            .in1(N__9304),
            .in2(N__16132),
            .in3(N__14693),
            .lcout(\c0.data_in_frame_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i10_LC_2_31_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i10_LC_2_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i10_LC_2_31_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i10_LC_2_31_2  (
            .in0(N__17064),
            .in1(N__10504),
            .in2(_gnd_net_),
            .in3(N__11806),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i24_LC_2_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i24_LC_2_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i24_LC_2_31_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i24_LC_2_31_3  (
            .in0(N__11439),
            .in1(N__17069),
            .in2(_gnd_net_),
            .in3(N__10602),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i16_LC_2_31_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i16_LC_2_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i16_LC_2_31_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i16_LC_2_31_4  (
            .in0(N__9408),
            .in1(N__15020),
            .in2(N__14722),
            .in3(N__10163),
            .lcout(\c0.data_in_field_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i34_LC_2_31_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i34_LC_2_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i34_LC_2_31_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i34_LC_2_31_5  (
            .in0(N__17019),
            .in1(N__10572),
            .in2(_gnd_net_),
            .in3(N__17458),
            .lcout(data_in_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i15_LC_2_31_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i15_LC_2_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i15_LC_2_31_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i15_LC_2_31_6  (
            .in0(N__17065),
            .in1(N__9219),
            .in2(_gnd_net_),
            .in3(N__9289),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_2_31_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_2_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_2_31_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_2_31_7  (
            .in0(N__14150),
            .in1(N__15143),
            .in2(N__9250),
            .in3(N__17683),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_R_49_LC_2_32_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_R_49_LC_2_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_R_49_LC_2_32_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_R_49_LC_2_32_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9233),
            .lcout(\c0.rx.r_Rx_Data_R ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22915),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_292_LC_2_32_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_292_LC_2_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_292_LC_2_32_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_292_LC_2_32_1  (
            .in0(N__10598),
            .in1(N__9218),
            .in2(N__11917),
            .in3(N__10538),
            .lcout(\c0.n26_adj_869 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i17_LC_2_32_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i17_LC_2_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i17_LC_2_32_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i17_LC_2_32_2  (
            .in0(N__17101),
            .in1(N__13792),
            .in2(_gnd_net_),
            .in3(N__9409),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22915),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_2_32_3 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_2_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_2_32_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i11_4_lut_LC_2_32_3  (
            .in0(N__11801),
            .in1(N__9942),
            .in2(N__11440),
            .in3(N__10680),
            .lcout(\c0.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_2_32_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_2_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_2_32_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_2_32_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9374),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22915),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i5_LC_2_32_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i5_LC_2_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i5_LC_2_32_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i5_LC_2_32_5  (
            .in0(N__17100),
            .in1(N__9367),
            .in2(_gnd_net_),
            .in3(N__9943),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22915),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i16_LC_2_32_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i16_LC_2_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i16_LC_2_32_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_in_0___i16_LC_2_32_6  (
            .in0(_gnd_net_),
            .in1(N__17099),
            .in2(N__9337),
            .in3(N__11435),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22915),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i3_LC_2_32_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i3_LC_2_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i3_LC_2_32_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i3_LC_2_32_7  (
            .in0(N__11913),
            .in1(N__17102),
            .in2(_gnd_net_),
            .in3(N__15079),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22915),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_4_lut_LC_3_22_0 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_4_lut_LC_3_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_4_lut_LC_3_22_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx2.i1_4_lut_4_lut_LC_3_22_0  (
            .in0(N__12410),
            .in1(N__10799),
            .in2(N__12649),
            .in3(N__10768),
            .lcout(n9_adj_939),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i5_LC_3_22_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i5_LC_3_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i5_LC_3_22_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i5_LC_3_22_1  (
            .in0(N__15223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10733),
            .lcout(\c0.tx2.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i8_LC_3_22_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i8_LC_3_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i8_LC_3_22_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i8_LC_3_22_3  (
            .in0(N__15224),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10715),
            .lcout(\c0.tx2.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i1_LC_3_22_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i1_LC_3_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i1_LC_3_22_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i1_LC_3_22_6  (
            .in0(_gnd_net_),
            .in1(N__10514),
            .in2(_gnd_net_),
            .in3(N__15222),
            .lcout(\c0.tx2.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4362_2_lut_3_lut_4_lut_LC_3_23_0 .C_ON=1'b0;
    defparam \c0.tx2.i4362_2_lut_3_lut_4_lut_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4362_2_lut_3_lut_4_lut_LC_3_23_0 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \c0.tx2.i4362_2_lut_3_lut_4_lut_LC_3_23_0  (
            .in0(N__12648),
            .in1(N__10802),
            .in2(N__12565),
            .in3(N__10769),
            .lcout(),
            .ltout(n4638_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Done_44_LC_3_23_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Done_44_LC_3_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Done_44_LC_3_23_1 .LUT_INIT=16'b1011101111111000;
    LogicCell40 \c0.tx2.r_Tx_Done_44_LC_3_23_1  (
            .in0(N__9449),
            .in1(N__9461),
            .in2(N__9452),
            .in3(N__12413),
            .lcout(tx2_done),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22873),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4459_LC_3_23_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4459_LC_3_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_4459_LC_3_23_2 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_4459_LC_3_23_2  (
            .in0(N__9443),
            .in1(N__15636),
            .in2(N__15785),
            .in3(N__11189),
            .lcout(\c0.n4819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_3_lut_4_lut_LC_3_23_3 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_3_lut_4_lut_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_3_lut_4_lut_LC_3_23_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx2.i2_2_lut_3_lut_4_lut_LC_3_23_3  (
            .in0(N__12528),
            .in1(N__12644),
            .in2(N__12701),
            .in3(N__12411),
            .lcout(n1030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4807_bdd_4_lut_LC_3_23_4 .C_ON=1'b0;
    defparam \c0.n4807_bdd_4_lut_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.n4807_bdd_4_lut_LC_3_23_4 .LUT_INIT=16'b1111110000001010;
    LogicCell40 \c0.n4807_bdd_4_lut_LC_3_23_4  (
            .in0(N__11141),
            .in1(N__9668),
            .in2(N__15786),
            .in3(N__9437),
            .lcout(),
            .ltout(tx2_data_2_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i2_LC_3_23_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i2_LC_3_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i2_LC_3_23_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx2.r_Tx_Data_i2_LC_3_23_5  (
            .in0(_gnd_net_),
            .in1(N__11227),
            .in2(N__9431),
            .in3(N__9428),
            .lcout(r_Tx_Data_2_adj_962),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22873),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_3_23_6.C_ON=1'b0;
    defparam i1_4_lut_LC_3_23_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_3_23_6.LUT_INIT=16'b1111111110101110;
    LogicCell40 i1_4_lut_LC_3_23_6 (
            .in0(N__12412),
            .in1(N__10748),
            .in2(N__12650),
            .in3(N__9416),
            .lcout(n6_adj_940),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i1_LC_3_24_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i1_LC_3_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i1_LC_3_24_0 .LUT_INIT=16'b1001110010001000;
    LogicCell40 \c0.tx2.r_Bit_Index_i1_LC_3_24_0  (
            .in0(N__9614),
            .in1(N__9580),
            .in2(N__9551),
            .in3(N__9637),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22877),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4157_4_lut_LC_3_24_1 .C_ON=1'b0;
    defparam \c0.tx2.i4157_4_lut_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4157_4_lut_LC_3_24_1 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \c0.tx2.i4157_4_lut_LC_3_24_1  (
            .in0(N__12414),
            .in1(N__11403),
            .in2(N__12570),
            .in3(N__12600),
            .lcout(n4512),
            .ltout(n4512_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4159_2_lut_LC_3_24_2.C_ON=1'b0;
    defparam i4159_2_lut_LC_3_24_2.SEQ_MODE=4'b0000;
    defparam i4159_2_lut_LC_3_24_2.LUT_INIT=16'b1111111111110000;
    LogicCell40 i4159_2_lut_LC_3_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9659),
            .in3(N__9633),
            .lcout(n4514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4191_3_lut_LC_3_24_3 .C_ON=1'b0;
    defparam \c0.i4191_3_lut_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4191_3_lut_LC_3_24_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4191_3_lut_LC_3_24_3  (
            .in0(N__15470),
            .in1(N__11357),
            .in2(_gnd_net_),
            .in3(N__10313),
            .lcout(\c0.n4546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4248_3_lut_LC_3_24_4 .C_ON=1'b0;
    defparam \c0.i4248_3_lut_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4248_3_lut_LC_3_24_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4248_3_lut_LC_3_24_4  (
            .in0(N__15519),
            .in1(N__13193),
            .in2(_gnd_net_),
            .in3(N__10343),
            .lcout(\c0.n4603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2099_4_lut_LC_3_24_5.C_ON=1'b0;
    defparam i2099_4_lut_LC_3_24_5.SEQ_MODE=4'b0000;
    defparam i2099_4_lut_LC_3_24_5.LUT_INIT=16'b1100110001100000;
    LogicCell40 i2099_4_lut_LC_3_24_5 (
            .in0(N__9579),
            .in1(N__9500),
            .in2(N__9638),
            .in3(N__9612),
            .lcout(),
            .ltout(n2326_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i2_LC_3_24_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i2_LC_3_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i2_LC_3_24_6 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i2_LC_3_24_6  (
            .in0(N__9501),
            .in1(N__9548),
            .in2(N__9623),
            .in3(N__9620),
            .lcout(r_Bit_Index_2_adj_955),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22877),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_24_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_24_7 .LUT_INIT=16'b1100110000100010;
    LogicCell40 \c0.tx2.r_Bit_Index_i0_LC_3_24_7  (
            .in0(N__12558),
            .in1(N__9544),
            .in2(_gnd_net_),
            .in3(N__9613),
            .lcout(r_Bit_Index_0_adj_956),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22877),
            .ce(),
            .sr(_gnd_net_));
    defparam i4167_3_lut_LC_3_25_1.C_ON=1'b0;
    defparam i4167_3_lut_LC_3_25_1.SEQ_MODE=4'b0000;
    defparam i4167_3_lut_LC_3_25_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 i4167_3_lut_LC_3_25_1 (
            .in0(N__11200),
            .in1(N__11011),
            .in2(_gnd_net_),
            .in3(N__9498),
            .lcout(),
            .ltout(n4522_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n4777_bdd_4_lut_LC_3_25_2.C_ON=1'b0;
    defparam n4777_bdd_4_lut_LC_3_25_2.SEQ_MODE=4'b0000;
    defparam n4777_bdd_4_lut_LC_3_25_2.LUT_INIT=16'b1110111001010000;
    LogicCell40 n4777_bdd_4_lut_LC_3_25_2 (
            .in0(N__9542),
            .in1(N__9602),
            .in2(N__9590),
            .in3(N__9587),
            .lcout(n4780),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_LC_3_25_3 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_LC_3_25_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx2.i2_3_lut_LC_3_25_3  (
            .in0(N__9581),
            .in1(N__9543),
            .in2(_gnd_net_),
            .in3(N__9499),
            .lcout(\c0.tx2.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_330_LC_3_25_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_330_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_330_LC_3_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_330_LC_3_25_5  (
            .in0(N__13495),
            .in1(N__13759),
            .in2(N__12047),
            .in3(N__9866),
            .lcout(\c0.n8_adj_880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4201_3_lut_LC_3_25_6 .C_ON=1'b0;
    defparam \c0.i4201_3_lut_LC_3_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4201_3_lut_LC_3_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4201_3_lut_LC_3_25_6  (
            .in0(N__15521),
            .in1(N__13448),
            .in2(_gnd_net_),
            .in3(N__9743),
            .lcout(\c0.n4556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_320_LC_3_26_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_320_LC_3_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_320_LC_3_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_320_LC_3_26_0  (
            .in0(N__10131),
            .in1(N__9895),
            .in2(N__13722),
            .in3(N__13598),
            .lcout(),
            .ltout(\c0.n10_adj_874_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_322_LC_3_26_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_322_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_322_LC_3_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_322_LC_3_26_1  (
            .in0(N__13645),
            .in1(N__10341),
            .in2(N__9716),
            .in3(N__9851),
            .lcout(\c0.n4469 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4212_3_lut_LC_3_26_2 .C_ON=1'b0;
    defparam \c0.i4212_3_lut_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4212_3_lut_LC_3_26_2 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \c0.i4212_3_lut_LC_3_26_2  (
            .in0(N__15513),
            .in1(N__10454),
            .in2(N__11663),
            .in3(_gnd_net_),
            .lcout(\c0.n4567 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i7_LC_3_26_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i7_LC_3_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i7_LC_3_26_3 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i7_LC_3_26_3  (
            .in0(N__9704),
            .in1(N__11661),
            .in2(N__14501),
            .in3(N__15027),
            .lcout(\c0.data_in_field_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22884),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_338_LC_3_26_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_338_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_338_LC_3_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_338_LC_3_26_4  (
            .in0(N__11474),
            .in1(N__10173),
            .in2(N__13265),
            .in3(N__10309),
            .lcout(\c0.n15_adj_885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4186_3_lut_LC_3_26_5 .C_ON=1'b0;
    defparam \c0.i4186_3_lut_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4186_3_lut_LC_3_26_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i4186_3_lut_LC_3_26_5  (
            .in0(N__10478),
            .in1(N__13297),
            .in2(_gnd_net_),
            .in3(N__15515),
            .lcout(\c0.n4541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4189_3_lut_LC_3_26_6 .C_ON=1'b0;
    defparam \c0.i4189_3_lut_LC_3_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4189_3_lut_LC_3_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4189_3_lut_LC_3_26_6  (
            .in0(N__15514),
            .in1(N__13530),
            .in2(_gnd_net_),
            .in3(N__10061),
            .lcout(\c0.n4544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_303_LC_3_27_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_303_LC_3_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_303_LC_3_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_303_LC_3_27_0  (
            .in0(N__11654),
            .in1(N__9887),
            .in2(_gnd_net_),
            .in3(N__9865),
            .lcout(\c0.n4408 ),
            .ltout(\c0.n4408_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_3_27_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_3_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_3_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_3_27_1  (
            .in0(N__11592),
            .in1(N__10018),
            .in2(N__9854),
            .in3(N__9850),
            .lcout(\c0.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_337_LC_3_27_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_337_LC_3_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_337_LC_3_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_337_LC_3_27_2  (
            .in0(N__11636),
            .in1(N__13151),
            .in2(N__16133),
            .in3(N__11771),
            .lcout(\c0.n16_adj_884 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_302_LC_3_27_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_302_LC_3_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_302_LC_3_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_302_LC_3_27_3  (
            .in0(N__9977),
            .in1(N__10266),
            .in2(N__12878),
            .in3(N__11684),
            .lcout(\c0.n4468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i19_LC_3_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i19_LC_3_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i19_LC_3_27_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i19_LC_3_27_5  (
            .in0(N__9839),
            .in1(N__15042),
            .in2(N__10277),
            .in3(N__14653),
            .lcout(\c0.data_in_field_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22890),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i26_LC_3_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i26_LC_3_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i26_LC_3_27_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i26_LC_3_27_6  (
            .in0(N__14652),
            .in1(N__15038),
            .in2(N__9809),
            .in3(N__13531),
            .lcout(\c0.data_in_field_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22890),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i21_LC_3_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i21_LC_3_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i21_LC_3_27_7 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i21_LC_3_27_7  (
            .in0(N__9776),
            .in1(N__11685),
            .in2(N__15047),
            .in3(N__14654),
            .lcout(\c0.data_in_field_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22890),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_308_LC_3_28_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_308_LC_3_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_308_LC_3_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_308_LC_3_28_0  (
            .in0(N__13636),
            .in1(N__10330),
            .in2(_gnd_net_),
            .in3(N__11172),
            .lcout(\c0.n1271 ),
            .ltout(\c0.n1271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_357_LC_3_28_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_357_LC_3_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_357_LC_3_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_357_LC_3_28_1  (
            .in0(N__11756),
            .in1(N__10120),
            .in2(N__9746),
            .in3(N__10060),
            .lcout(\c0.n4429 ),
            .ltout(\c0.n4429_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_341_LC_3_28_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_341_LC_3_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_341_LC_3_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_341_LC_3_28_2  (
            .in0(N__13022),
            .in1(N__10211),
            .in2(N__10034),
            .in3(N__12895),
            .lcout(\c0.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_339_LC_3_28_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_339_LC_3_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_339_LC_3_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_339_LC_3_28_3  (
            .in0(N__10031),
            .in1(N__10020),
            .in2(N__9992),
            .in3(N__9978),
            .lcout(\c0.n4430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i25_LC_3_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i25_LC_3_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i25_LC_3_28_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i25_LC_3_28_4  (
            .in0(N__10552),
            .in1(N__14997),
            .in2(N__14713),
            .in3(N__13284),
            .lcout(\c0.data_in_field_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22895),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_297_LC_3_28_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_297_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_297_LC_3_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_297_LC_3_28_6  (
            .in0(N__14005),
            .in1(N__13283),
            .in2(N__10422),
            .in3(N__9956),
            .lcout(\c0.n1296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i34_LC_3_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i34_LC_3_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i34_LC_3_28_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i34_LC_3_28_7  (
            .in0(N__10331),
            .in1(N__11383),
            .in2(N__15043),
            .in3(N__14665),
            .lcout(\c0.data_in_field_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22895),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i4_LC_3_29_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i4_LC_3_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i4_LC_3_29_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i4_LC_3_29_0  (
            .in0(N__9950),
            .in1(N__14935),
            .in2(N__14712),
            .in3(N__11761),
            .lcout(\c0.data_in_field_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22901),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_310_LC_3_29_1 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_310_LC_3_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_310_LC_3_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_310_LC_3_29_1  (
            .in0(N__10987),
            .in1(N__9919),
            .in2(_gnd_net_),
            .in3(N__10470),
            .lcout(\c0.n1261 ),
            .ltout(\c0.n1261_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_312_LC_3_29_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_312_LC_3_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_312_LC_3_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_312_LC_3_29_2  (
            .in0(N__13553),
            .in1(N__10445),
            .in2(N__9899),
            .in3(N__11892),
            .lcout(\c0.n4390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i53_LC_3_29_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i53_LC_3_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i53_LC_3_29_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i53_LC_3_29_3  (
            .in0(N__14934),
            .in1(N__14655),
            .in2(N__10202),
            .in3(N__12284),
            .lcout(\c0.data_in_frame_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22901),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i43_LC_3_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i43_LC_3_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i43_LC_3_29_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i43_LC_3_29_4  (
            .in0(N__13554),
            .in1(N__16562),
            .in2(N__14711),
            .in3(N__14936),
            .lcout(\c0.data_in_field_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22901),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_294_LC_3_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_294_LC_3_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_294_LC_3_29_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_294_LC_3_29_5  (
            .in0(N__12817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13432),
            .lcout(\c0.n4411 ),
            .ltout(\c0.n4411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_354_LC_3_29_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_354_LC_3_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_354_LC_3_29_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_354_LC_3_29_6  (
            .in0(N__11624),
            .in1(N__10233),
            .in2(N__10205),
            .in3(N__12779),
            .lcout(\c0.n4399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4240_3_lut_LC_3_29_7 .C_ON=1'b0;
    defparam \c0.i4240_3_lut_LC_3_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4240_3_lut_LC_3_29_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.i4240_3_lut_LC_3_29_7  (
            .in0(N__10198),
            .in1(N__15528),
            .in2(_gnd_net_),
            .in3(N__10357),
            .lcout(\c0.n4595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_298_LC_3_30_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_298_LC_3_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_298_LC_3_30_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_298_LC_3_30_0  (
            .in0(N__10119),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11757),
            .lcout(),
            .ltout(\c0.n1340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_324_LC_3_30_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_324_LC_3_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_324_LC_3_30_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_324_LC_3_30_1  (
            .in0(N__13045),
            .in1(N__10250),
            .in2(N__10178),
            .in3(N__13068),
            .lcout(\c0.n4445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_306_LC_3_30_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_306_LC_3_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_306_LC_3_30_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_306_LC_3_30_2  (
            .in0(N__10154),
            .in1(N__10295),
            .in2(N__10130),
            .in3(N__10052),
            .lcout(\c0.n8_adj_872 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i1_LC_3_30_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i1_LC_3_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i1_LC_3_30_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i1_LC_3_30_3  (
            .in0(N__15009),
            .in1(N__14694),
            .in2(N__12834),
            .in3(N__10685),
            .lcout(\c0.data_in_field_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22909),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i18_LC_3_30_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i18_LC_3_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i18_LC_3_30_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i18_LC_3_30_4  (
            .in0(N__10091),
            .in1(N__15012),
            .in2(N__14724),
            .in3(N__10053),
            .lcout(\c0.data_in_field_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22909),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i32_LC_3_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i32_LC_3_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i32_LC_3_30_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i32_LC_3_30_5  (
            .in0(N__15010),
            .in1(N__14255),
            .in2(N__10999),
            .in3(N__14695),
            .lcout(\c0.data_in_field_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22909),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i17_LC_3_30_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i17_LC_3_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i17_LC_3_30_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i17_LC_3_30_6  (
            .in0(N__10505),
            .in1(N__15011),
            .in2(N__14723),
            .in3(N__10474),
            .lcout(\c0.data_in_field_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22909),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_317_LC_3_30_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_317_LC_3_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_317_LC_3_30_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_317_LC_3_30_7  (
            .in0(N__11339),
            .in1(N__10446),
            .in2(N__14014),
            .in3(N__11272),
            .lcout(\c0.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4192_3_lut_LC_3_31_0 .C_ON=1'b0;
    defparam \c0.i4192_3_lut_LC_3_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4192_3_lut_LC_3_31_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4192_3_lut_LC_3_31_0  (
            .in0(N__15545),
            .in1(N__10423),
            .in2(_gnd_net_),
            .in3(N__10276),
            .lcout(\c0.n4547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i3_LC_3_31_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i3_LC_3_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i3_LC_3_31_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i3_LC_3_31_1  (
            .in0(N__10302),
            .in1(N__10382),
            .in2(N__14669),
            .in3(N__14978),
            .lcout(\c0.data_in_field_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22916),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i61_LC_3_31_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i61_LC_3_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i61_LC_3_31_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i61_LC_3_31_2  (
            .in0(N__14977),
            .in1(N__14570),
            .in2(N__12311),
            .in3(N__10358),
            .lcout(\c0.data_in_frame_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22916),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_314_LC_3_31_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_314_LC_3_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_314_LC_3_31_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_314_LC_3_31_4  (
            .in0(N__10342),
            .in1(N__10301),
            .in2(N__12310),
            .in3(N__10275),
            .lcout(\c0.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i45_LC_3_31_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i45_LC_3_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i45_LC_3_31_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i45_LC_3_31_5  (
            .in0(N__11983),
            .in1(N__17024),
            .in2(_gnd_net_),
            .in3(N__12180),
            .lcout(data_in_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22916),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_349_LC_3_31_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_349_LC_3_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_349_LC_3_31_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_349_LC_3_31_6  (
            .in0(N__13433),
            .in1(N__10232),
            .in2(_gnd_net_),
            .in3(N__12818),
            .lcout(\c0.n1280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_3_31_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_3_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_3_31_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_3_31_7  (
            .in0(N__15142),
            .in1(N__15110),
            .in2(N__10700),
            .in3(N__17711),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22916),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i46_LC_3_32_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i46_LC_3_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i46_LC_3_32_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i46_LC_3_32_1  (
            .in0(N__17058),
            .in1(N__10653),
            .in2(_gnd_net_),
            .in3(N__12273),
            .lcout(data_in_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22923),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i2_LC_3_32_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i2_LC_3_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i2_LC_3_32_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i2_LC_3_32_2  (
            .in0(N__11805),
            .in1(N__17059),
            .in2(_gnd_net_),
            .in3(N__10684),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22923),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i38_LC_3_32_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i38_LC_3_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i38_LC_3_32_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i38_LC_3_32_3  (
            .in0(N__17057),
            .in1(N__10654),
            .in2(_gnd_net_),
            .in3(N__10621),
            .lcout(data_in_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22923),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_3_32_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_3_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_3_32_4 .LUT_INIT=16'b0111101001110000;
    LogicCell40 \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_3_32_4  (
            .in0(N__17555),
            .in1(N__17378),
            .in2(N__17778),
            .in3(N__16046),
            .lcout(),
            .ltout(\c0.rx.n4873_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.n4873_bdd_4_lut_4_lut_LC_3_32_5 .C_ON=1'b0;
    defparam \c0.rx.n4873_bdd_4_lut_4_lut_LC_3_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.n4873_bdd_4_lut_4_lut_LC_3_32_5 .LUT_INIT=16'b1111000111000001;
    LogicCell40 \c0.rx.n4873_bdd_4_lut_4_lut_LC_3_32_5  (
            .in0(N__17686),
            .in1(N__17556),
            .in2(N__10610),
            .in3(N__17816),
            .lcout(\c0.rx.n4876 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i32_LC_3_32_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i32_LC_3_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i32_LC_3_32_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i32_LC_3_32_6  (
            .in0(N__10603),
            .in1(N__11531),
            .in2(_gnd_net_),
            .in3(N__17060),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22923),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i26_LC_3_32_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i26_LC_3_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i26_LC_3_32_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i26_LC_3_32_7  (
            .in0(N__17056),
            .in1(N__10573),
            .in2(_gnd_net_),
            .in3(N__10545),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22923),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_2_lut_LC_4_21_0 .C_ON=1'b1;
    defparam \c0.tx2.add_59_2_lut_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_2_lut_LC_4_21_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_2_lut_LC_4_21_0  (
            .in0(N__10946),
            .in1(N__10945),
            .in2(N__12455),
            .in3(N__10517),
            .lcout(n1768),
            .ltout(),
            .carryin(bfn_4_21_0_),
            .carryout(\c0.tx2.n3891 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_3_lut_LC_4_21_1 .C_ON=1'b1;
    defparam \c0.tx2.add_59_3_lut_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_3_lut_LC_4_21_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_3_lut_LC_4_21_1  (
            .in0(N__10897),
            .in1(N__10896),
            .in2(N__12459),
            .in3(N__10508),
            .lcout(n1710),
            .ltout(),
            .carryin(\c0.tx2.n3891 ),
            .carryout(\c0.tx2.n3892 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_4_lut_LC_4_21_2 .C_ON=1'b1;
    defparam \c0.tx2.add_59_4_lut_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_4_lut_LC_4_21_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_4_lut_LC_4_21_2  (
            .in0(N__10934),
            .in1(N__10933),
            .in2(N__12456),
            .in3(N__10742),
            .lcout(n1707),
            .ltout(),
            .carryin(\c0.tx2.n3892 ),
            .carryout(\c0.tx2.n3893 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_5_lut_LC_4_21_3 .C_ON=1'b1;
    defparam \c0.tx2.add_59_5_lut_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_5_lut_LC_4_21_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_5_lut_LC_4_21_3  (
            .in0(N__10877),
            .in1(N__10876),
            .in2(N__12460),
            .in3(N__10739),
            .lcout(n1704),
            .ltout(),
            .carryin(\c0.tx2.n3893 ),
            .carryout(\c0.tx2.n3894 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_6_lut_LC_4_21_4 .C_ON=1'b1;
    defparam \c0.tx2.add_59_6_lut_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_6_lut_LC_4_21_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_6_lut_LC_4_21_4  (
            .in0(N__10850),
            .in1(N__10849),
            .in2(N__12457),
            .in3(N__10736),
            .lcout(n1701),
            .ltout(),
            .carryin(\c0.tx2.n3894 ),
            .carryout(\c0.tx2.n3895 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_7_lut_LC_4_21_5 .C_ON=1'b1;
    defparam \c0.tx2.add_59_7_lut_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_7_lut_LC_4_21_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_7_lut_LC_4_21_5  (
            .in0(N__10916),
            .in1(N__10915),
            .in2(N__12461),
            .in3(N__10727),
            .lcout(n1698),
            .ltout(),
            .carryin(\c0.tx2.n3895 ),
            .carryout(\c0.tx2.n3896 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_8_lut_LC_4_21_6 .C_ON=1'b1;
    defparam \c0.tx2.add_59_8_lut_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_8_lut_LC_4_21_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_8_lut_LC_4_21_6  (
            .in0(N__15194),
            .in1(N__15193),
            .in2(N__12458),
            .in3(N__10724),
            .lcout(n1695),
            .ltout(),
            .carryin(\c0.tx2.n3896 ),
            .carryout(\c0.tx2.n3897 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_9_lut_LC_4_21_7 .C_ON=1'b1;
    defparam \c0.tx2.add_59_9_lut_LC_4_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_9_lut_LC_4_21_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_9_lut_LC_4_21_7  (
            .in0(N__10823),
            .in1(N__10822),
            .in2(N__12462),
            .in3(N__10721),
            .lcout(n1692),
            .ltout(),
            .carryin(\c0.tx2.n3897 ),
            .carryout(\c0.tx2.n3898 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_10_lut_LC_4_22_0 .C_ON=1'b0;
    defparam \c0.tx2.add_59_10_lut_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_10_lut_LC_4_22_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_10_lut_LC_4_22_0  (
            .in0(N__10800),
            .in1(N__10801),
            .in2(N__12448),
            .in3(N__10718),
            .lcout(n1689),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i3_LC_4_22_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i3_LC_4_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i3_LC_4_22_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i3_LC_4_22_1  (
            .in0(N__15227),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10709),
            .lcout(\c0.tx2.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22874),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i2_LC_4_22_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i2_LC_4_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i2_LC_4_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i2_LC_4_22_2  (
            .in0(_gnd_net_),
            .in1(N__10958),
            .in2(_gnd_net_),
            .in3(N__15226),
            .lcout(\c0.tx2.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22874),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i0_LC_4_22_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i0_LC_4_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i0_LC_4_22_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i0_LC_4_22_3  (
            .in0(N__15225),
            .in1(N__10952),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.tx2.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22874),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_LC_4_22_4 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_LC_4_22_4 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \c0.tx2.i1_4_lut_LC_4_22_4  (
            .in0(N__10932),
            .in1(N__10914),
            .in2(N__10898),
            .in3(N__10875),
            .lcout(),
            .ltout(\c0.tx2.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2675_4_lut_LC_4_22_5 .C_ON=1'b0;
    defparam \c0.tx2.i2675_4_lut_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2675_4_lut_LC_4_22_5 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.tx2.i2675_4_lut_LC_4_22_5  (
            .in0(N__15192),
            .in1(N__10848),
            .in2(N__10859),
            .in3(N__10821),
            .lcout(\c0.tx2.n2902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i4_LC_4_22_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i4_LC_4_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i4_LC_4_22_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i4_LC_4_22_6  (
            .in0(_gnd_net_),
            .in1(N__10856),
            .in2(_gnd_net_),
            .in3(N__15228),
            .lcout(\c0.tx2.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22874),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i7_LC_4_22_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i7_LC_4_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i7_LC_4_22_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.tx2.r_Clock_Count__i7_LC_4_22_7  (
            .in0(N__15229),
            .in1(_gnd_net_),
            .in2(N__10832),
            .in3(_gnd_net_),
            .lcout(\c0.tx2.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22874),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2677_2_lut_LC_4_23_0 .C_ON=1'b0;
    defparam \c0.tx2.i2677_2_lut_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2677_2_lut_LC_4_23_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx2.i2677_2_lut_LC_4_23_0  (
            .in0(_gnd_net_),
            .in1(N__10797),
            .in2(_gnd_net_),
            .in3(N__10766),
            .lcout(r_SM_Main_2_N_759_1),
            .ltout(r_SM_Main_2_N_759_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i2_LC_4_23_1 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i2_LC_4_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i2_LC_4_23_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.tx2.r_SM_Main_i2_LC_4_23_1  (
            .in0(N__12623),
            .in1(N__12524),
            .in2(N__10805),
            .in3(N__12409),
            .lcout(r_SM_Main_2_adj_952),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22878),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_3_lut_4_lut_LC_4_23_2 .C_ON=1'b0;
    defparam \c0.tx2.i1_3_lut_4_lut_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_3_lut_4_lut_LC_4_23_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx2.i1_3_lut_4_lut_LC_4_23_2  (
            .in0(N__12407),
            .in1(N__10798),
            .in2(N__12553),
            .in3(N__10767),
            .lcout(n4_adj_965),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4188_3_lut_LC_4_23_3 .C_ON=1'b0;
    defparam \c0.i4188_3_lut_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4188_3_lut_LC_4_23_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4188_3_lut_LC_4_23_3  (
            .in0(N__15430),
            .in1(N__14315),
            .in2(_gnd_net_),
            .in3(N__11897),
            .lcout(\c0.n4543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i1_LC_4_23_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i1_LC_4_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i1_LC_4_23_4 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \c0.tx2.r_SM_Main_i1_LC_4_23_4  (
            .in0(N__12408),
            .in1(N__12624),
            .in2(N__12554),
            .in3(N__11411),
            .lcout(r_SM_Main_1_adj_953),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22878),
            .ce(),
            .sr(_gnd_net_));
    defparam i4164_4_lut_LC_4_23_6.C_ON=1'b0;
    defparam i4164_4_lut_LC_4_23_6.SEQ_MODE=4'b0000;
    defparam i4164_4_lut_LC_4_23_6.LUT_INIT=16'b1101110101000000;
    LogicCell40 i4164_4_lut_LC_4_23_6 (
            .in0(N__11113),
            .in1(N__11134),
            .in2(N__11069),
            .in3(N__11089),
            .lcout(n4519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4165_4_lut_LC_4_23_7.C_ON=1'b0;
    defparam i4165_4_lut_LC_4_23_7.SEQ_MODE=4'b0000;
    defparam i4165_4_lut_LC_4_23_7.LUT_INIT=16'b1111110111100000;
    LogicCell40 i4165_4_lut_LC_4_23_7 (
            .in0(N__11135),
            .in1(N__11114),
            .in2(N__11093),
            .in3(N__11068),
            .lcout(n4520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_4_24_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_4_24_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_LC_4_24_0  (
            .in0(N__15604),
            .in1(N__11045),
            .in2(N__15777),
            .in3(N__10964),
            .lcout(),
            .ltout(\c0.n4855_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4855_bdd_4_lut_LC_4_24_1 .C_ON=1'b0;
    defparam \c0.n4855_bdd_4_lut_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.n4855_bdd_4_lut_LC_4_24_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n4855_bdd_4_lut_LC_4_24_1  (
            .in0(N__11030),
            .in1(N__15747),
            .in2(N__11018),
            .in3(N__11576),
            .lcout(),
            .ltout(tx2_data_0_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i0_LC_4_24_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i0_LC_4_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i0_LC_4_24_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx2.r_Tx_Data_i0_LC_4_24_2  (
            .in0(_gnd_net_),
            .in1(N__11229),
            .in2(N__11015),
            .in3(N__11012),
            .lcout(r_Tx_Data_0_adj_964),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22881),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4224_3_lut_LC_4_24_3 .C_ON=1'b0;
    defparam \c0.i4224_3_lut_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4224_3_lut_LC_4_24_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4224_3_lut_LC_4_24_3  (
            .in0(N__15469),
            .in1(N__13976),
            .in2(_gnd_net_),
            .in3(N__11000),
            .lcout(\c0.n4579 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4194_3_lut_LC_4_24_4 .C_ON=1'b0;
    defparam \c0.i4194_3_lut_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4194_3_lut_LC_4_24_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4194_3_lut_LC_4_24_4  (
            .in0(N__15432),
            .in1(N__14018),
            .in2(_gnd_net_),
            .in3(N__11765),
            .lcout(),
            .ltout(\c0.n4549_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4819_bdd_4_lut_LC_4_24_5 .C_ON=1'b0;
    defparam \c0.n4819_bdd_4_lut_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n4819_bdd_4_lut_LC_4_24_5 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \c0.n4819_bdd_4_lut_LC_4_24_5  (
            .in0(N__11261),
            .in1(N__15746),
            .in2(N__11255),
            .in3(N__11156),
            .lcout(),
            .ltout(tx2_data_4_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i4_LC_4_24_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i4_LC_4_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i4_LC_4_24_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx2.r_Tx_Data_i4_LC_4_24_6  (
            .in0(_gnd_net_),
            .in1(N__11230),
            .in2(N__11204),
            .in3(N__11201),
            .lcout(r_Tx_Data_4_adj_960),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22881),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4242_3_lut_LC_4_24_7 .C_ON=1'b0;
    defparam \c0.i4242_3_lut_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4242_3_lut_LC_4_24_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4242_3_lut_LC_4_24_7  (
            .in0(N__15468),
            .in1(N__12164),
            .in2(_gnd_net_),
            .in3(N__13613),
            .lcout(\c0.n4597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4397_2_lut_LC_4_25_0 .C_ON=1'b0;
    defparam \c0.i4397_2_lut_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4397_2_lut_LC_4_25_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \c0.i4397_2_lut_LC_4_25_0  (
            .in0(_gnd_net_),
            .in1(N__14405),
            .in2(_gnd_net_),
            .in3(N__13091),
            .lcout(\c0.n1675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i48_LC_4_25_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i48_LC_4_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i48_LC_4_25_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i48_LC_4_25_1  (
            .in0(N__17087),
            .in1(N__11487),
            .in2(_gnd_net_),
            .in3(N__13681),
            .lcout(data_in_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22885),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4195_3_lut_LC_4_25_2 .C_ON=1'b0;
    defparam \c0.i4195_3_lut_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4195_3_lut_LC_4_25_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4195_3_lut_LC_4_25_2  (
            .in0(N__15431),
            .in1(N__13223),
            .in2(_gnd_net_),
            .in3(N__11183),
            .lcout(\c0.n4550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_wait_for_transmission_621_LC_4_25_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_wait_for_transmission_621_LC_4_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_wait_for_transmission_621_LC_4_25_3 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \c0.FRAME_MATCHER_wait_for_transmission_621_LC_4_25_3  (
            .in0(N__14406),
            .in1(N__12710),
            .in2(N__13099),
            .in3(N__15332),
            .lcout(\c0.FRAME_MATCHER_wait_for_transmission ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22885),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i639_4_lut_LC_4_25_4 .C_ON=1'b0;
    defparam \c0.tx2.i639_4_lut_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i639_4_lut_LC_4_25_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.tx2.i639_4_lut_LC_4_25_4  (
            .in0(N__11150),
            .in1(N__12559),
            .in2(N__12694),
            .in3(N__11412),
            .lcout(),
            .ltout(n865_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i0_LC_4_25_5 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i0_LC_4_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i0_LC_4_25_5 .LUT_INIT=16'b0000000001110100;
    LogicCell40 \c0.tx2.r_SM_Main_i0_LC_4_25_5  (
            .in0(N__11414),
            .in1(N__12619),
            .in2(N__11144),
            .in3(N__12463),
            .lcout(r_SM_Main_0_adj_954),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22885),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4383_3_lut_4_lut_4_lut_LC_4_25_6 .C_ON=1'b0;
    defparam \c0.tx2.i4383_3_lut_4_lut_4_lut_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4383_3_lut_4_lut_4_lut_LC_4_25_6 .LUT_INIT=16'b1100001000000010;
    LogicCell40 \c0.tx2.i4383_3_lut_4_lut_4_lut_LC_4_25_6  (
            .in0(N__12688),
            .in1(N__12560),
            .in2(N__12638),
            .in3(N__11413),
            .lcout(),
            .ltout(n4366_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_47_LC_4_25_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_47_LC_4_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_47_LC_4_25_7 .LUT_INIT=16'b1100110001011100;
    LogicCell40 \c0.tx2.r_Tx_Active_47_LC_4_25_7  (
            .in0(N__12561),
            .in1(N__12725),
            .in2(N__11387),
            .in3(N__12464),
            .lcout(tx2_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22885),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i64_LC_4_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i64_LC_4_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i64_LC_4_26_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i64_LC_4_26_0  (
            .in0(N__13712),
            .in1(N__12065),
            .in2(_gnd_net_),
            .in3(N__17089),
            .lcout(data_in_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22891),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i35_LC_4_26_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i35_LC_4_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i35_LC_4_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i35_LC_4_26_1  (
            .in0(N__17088),
            .in1(N__14173),
            .in2(_gnd_net_),
            .in3(N__11373),
            .lcout(data_in_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22891),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_329_LC_4_26_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_329_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_329_LC_4_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_329_LC_4_26_2  (
            .in0(N__13752),
            .in1(N__11356),
            .in2(N__13907),
            .in3(N__13526),
            .lcout(),
            .ltout(\c0.n8_adj_879_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_adj_331_LC_4_26_3 .C_ON=1'b0;
    defparam \c0.i4_3_lut_adj_331_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_adj_331_LC_4_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i4_3_lut_adj_331_LC_4_26_3  (
            .in0(_gnd_net_),
            .in1(N__11979),
            .in2(N__11312),
            .in3(N__13263),
            .lcout(),
            .ltout(\c0.n4451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_336_LC_4_26_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_336_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_336_LC_4_26_4 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i5_4_lut_adj_336_LC_4_26_4  (
            .in0(N__15853),
            .in1(N__11702),
            .in2(N__11309),
            .in3(N__11306),
            .lcout(\c0.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_295_LC_4_26_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_295_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_295_LC_4_26_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_295_LC_4_26_5  (
            .in0(N__13184),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13222),
            .lcout(),
            .ltout(\c0.n1357_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_333_LC_4_26_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_333_LC_4_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_333_LC_4_26_6 .LUT_INIT=16'b1011011101111011;
    LogicCell40 \c0.i6_4_lut_adj_333_LC_4_26_6  (
            .in0(N__11297),
            .in1(N__11288),
            .in2(N__11282),
            .in3(N__11279),
            .lcout(\c0.n22_adj_881 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_346_LC_4_27_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_346_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_346_LC_4_27_0 .LUT_INIT=16'b1011011101111011;
    LogicCell40 \c0.i1_4_lut_adj_346_LC_4_27_0  (
            .in0(N__11564),
            .in1(N__11558),
            .in2(N__11552),
            .in3(N__11543),
            .lcout(),
            .ltout(\c0.n17_adj_889_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_352_LC_4_27_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_352_LC_4_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_352_LC_4_27_1 .LUT_INIT=16'b1111011111111101;
    LogicCell40 \c0.i9_4_lut_adj_352_LC_4_27_1  (
            .in0(N__13382),
            .in1(N__11453),
            .in2(N__11537),
            .in3(N__12752),
            .lcout(\c0.n25_adj_893 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_300_LC_4_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_300_LC_4_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_300_LC_4_27_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_300_LC_4_27_2  (
            .in0(N__13972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12037),
            .lcout(),
            .ltout(\c0.n4387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_325_LC_4_27_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_325_LC_4_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_325_LC_4_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_325_LC_4_27_3  (
            .in0(N__13185),
            .in1(N__12283),
            .in2(N__11534),
            .in3(N__11470),
            .lcout(\c0.n4388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i39_LC_4_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i39_LC_4_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i39_LC_4_27_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i39_LC_4_27_4  (
            .in0(N__14464),
            .in1(N__15035),
            .in2(N__11530),
            .in3(N__12038),
            .lcout(\c0.data_in_field_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22896),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i47_LC_4_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i47_LC_4_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i47_LC_4_27_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i47_LC_4_27_5  (
            .in0(N__15034),
            .in1(N__14465),
            .in2(N__12877),
            .in3(N__11497),
            .lcout(\c0.data_in_field_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22896),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_345_LC_4_27_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_345_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_345_LC_4_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_345_LC_4_27_7  (
            .in0(N__13076),
            .in1(N__13264),
            .in2(N__17276),
            .in3(N__11469),
            .lcout(\c0.n11_adj_888 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i23_LC_4_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i23_LC_4_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i23_LC_4_28_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i23_LC_4_28_0  (
            .in0(N__13367),
            .in1(N__15031),
            .in2(N__11447),
            .in3(N__14472),
            .lcout(\c0.data_in_field_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22902),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i28_LC_4_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i28_LC_4_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i28_LC_4_28_1 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i28_LC_4_28_1  (
            .in0(N__15029),
            .in1(N__12139),
            .in2(N__14578),
            .in3(N__13221),
            .lcout(\c0.data_in_field_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22902),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i9_LC_4_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i9_LC_4_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i9_LC_4_28_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i9_LC_4_28_2  (
            .in0(N__13481),
            .in1(N__15032),
            .in2(N__11813),
            .in3(N__14473),
            .lcout(\c0.data_in_field_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22902),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_304_LC_4_28_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_304_LC_4_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_304_LC_4_28_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_304_LC_4_28_3  (
            .in0(_gnd_net_),
            .in1(N__13525),
            .in2(_gnd_net_),
            .in3(N__13366),
            .lcout(),
            .ltout(\c0.n8_adj_871_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_4_28_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_4_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_4_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_LC_4_28_4  (
            .in0(N__13480),
            .in1(N__13742),
            .in2(N__11780),
            .in3(N__11777),
            .lcout(\c0.n1418 ),
            .ltout(\c0.n1418_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_309_LC_4_28_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_309_LC_4_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_309_LC_4_28_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_309_LC_4_28_5  (
            .in0(N__11755),
            .in1(N__15943),
            .in2(N__11729),
            .in3(N__13393),
            .lcout(\c0.n4474 ),
            .ltout(\c0.n4474_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_4_28_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_4_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_4_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_LC_4_28_6  (
            .in0(_gnd_net_),
            .in1(N__13673),
            .in2(N__11726),
            .in3(N__13183),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i38_LC_4_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i38_LC_4_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i38_LC_4_28_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i38_LC_4_28_7  (
            .in0(N__15030),
            .in1(N__11723),
            .in2(N__14579),
            .in3(N__12007),
            .lcout(\c0.data_in_field_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22902),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_299_LC_4_29_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_299_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_299_LC_4_29_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_299_LC_4_29_0  (
            .in0(_gnd_net_),
            .in1(N__12003),
            .in2(_gnd_net_),
            .in3(N__11602),
            .lcout(\c0.n4396 ),
            .ltout(\c0.n4396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_316_LC_4_29_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_316_LC_4_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_316_LC_4_29_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_316_LC_4_29_1  (
            .in0(N__16751),
            .in1(N__11692),
            .in2(N__11666),
            .in3(N__11662),
            .lcout(\c0.n12_adj_873 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4215_3_lut_LC_4_29_2 .C_ON=1'b0;
    defparam \c0.i4215_3_lut_LC_4_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4215_3_lut_LC_4_29_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4215_3_lut_LC_4_29_2  (
            .in0(N__15510),
            .in1(N__11635),
            .in2(_gnd_net_),
            .in3(N__11603),
            .lcout(\c0.n4570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i29_LC_4_29_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i29_LC_4_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i29_LC_4_29_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i29_LC_4_29_3  (
            .in0(N__11943),
            .in1(N__17062),
            .in2(_gnd_net_),
            .in3(N__12137),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22910),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_353_LC_4_29_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_353_LC_4_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_353_LC_4_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_353_LC_4_29_4  (
            .in0(N__12042),
            .in1(N__12002),
            .in2(N__14311),
            .in3(N__13963),
            .lcout(\c0.n1290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i53_LC_4_29_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i53_LC_4_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i53_LC_4_29_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i53_LC_4_29_5  (
            .in0(N__11978),
            .in1(N__13821),
            .in2(_gnd_net_),
            .in3(N__17063),
            .lcout(data_in_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22910),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i37_LC_4_29_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i37_LC_4_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i37_LC_4_29_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i37_LC_4_29_6  (
            .in0(N__17061),
            .in1(N__12191),
            .in2(_gnd_net_),
            .in3(N__11944),
            .lcout(data_in_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22910),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_LC_4_29_7 .C_ON=1'b0;
    defparam \c0.i4_3_lut_LC_4_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_LC_4_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_3_lut_LC_4_29_7  (
            .in0(N__11891),
            .in1(N__12159),
            .in2(_gnd_net_),
            .in3(N__11927),
            .lcout(\c0.n1267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i2_LC_4_30_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i2_LC_4_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i2_LC_4_30_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i2_LC_4_30_0  (
            .in0(N__11921),
            .in1(N__15016),
            .in2(N__14590),
            .in3(N__11896),
            .lcout(\c0.data_in_field_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22917),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i57_LC_4_30_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i57_LC_4_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i57_LC_4_30_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i57_LC_4_30_1  (
            .in0(N__15015),
            .in1(N__14486),
            .in2(N__11870),
            .in3(N__17272),
            .lcout(\c0.data_in_frame_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22917),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4252_3_lut_LC_4_30_2 .C_ON=1'b0;
    defparam \c0.i4252_3_lut_LC_4_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4252_3_lut_LC_4_30_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4252_3_lut_LC_4_30_2  (
            .in0(N__15544),
            .in1(N__11866),
            .in2(_gnd_net_),
            .in3(N__12202),
            .lcout(\c0.n4607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i30_LC_4_30_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i30_LC_4_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i30_LC_4_30_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i30_LC_4_30_3  (
            .in0(N__15013),
            .in1(N__11843),
            .in2(N__13447),
            .in3(N__14493),
            .lcout(\c0.data_in_field_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22917),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i49_LC_4_30_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i49_LC_4_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i49_LC_4_30_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i49_LC_4_30_4  (
            .in0(N__12203),
            .in1(N__16762),
            .in2(N__14591),
            .in3(N__15018),
            .lcout(\c0.data_in_frame_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22917),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i44_LC_4_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i44_LC_4_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i44_LC_4_30_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i44_LC_4_30_5  (
            .in0(N__15014),
            .in1(N__14485),
            .in2(N__12190),
            .in3(N__12163),
            .lcout(\c0.data_in_field_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22917),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i40_LC_4_30_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i40_LC_4_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i40_LC_4_30_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i40_LC_4_30_6  (
            .in0(N__14484),
            .in1(N__15017),
            .in2(N__14276),
            .in3(N__13971),
            .lcout(\c0.data_in_field_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22917),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i21_LC_4_30_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i21_LC_4_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i21_LC_4_30_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i21_LC_4_30_7  (
            .in0(N__12138),
            .in1(N__16996),
            .in2(_gnd_net_),
            .in3(N__12104),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22917),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_4_31_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_4_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_4_31_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_4_31_0  (
            .in0(N__15127),
            .in1(N__14142),
            .in2(N__13852),
            .in3(N__17707),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22924),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_4_31_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_4_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_4_31_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_4_31_1  (
            .in0(N__17705),
            .in1(N__15128),
            .in2(N__12077),
            .in3(N__15105),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22924),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i62_LC_4_31_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i62_LC_4_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i62_LC_4_31_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i62_LC_4_31_2  (
            .in0(N__17023),
            .in1(N__12073),
            .in2(_gnd_net_),
            .in3(N__12308),
            .lcout(data_in_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22924),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i57_LC_4_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i57_LC_4_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i57_LC_4_31_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i57_LC_4_31_3  (
            .in0(N__17022),
            .in1(N__15155),
            .in2(_gnd_net_),
            .in3(N__16118),
            .lcout(data_in_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22924),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_4_31_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_4_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_4_31_4 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_4_31_4  (
            .in0(N__15106),
            .in1(N__14288),
            .in2(N__12064),
            .in3(N__17708),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22924),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_4_31_5 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_4_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_4_31_5 .LUT_INIT=16'b1101110110011001;
    LogicCell40 \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_4_31_5  (
            .in0(N__12639),
            .in1(N__12571),
            .in2(_gnd_net_),
            .in3(N__12476),
            .lcout(),
            .ltout(n3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_31_6 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_31_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.tx2.o_Tx_Serial_45_LC_4_31_6  (
            .in0(N__12449),
            .in1(_gnd_net_),
            .in2(N__12341),
            .in3(N__14049),
            .lcout(tx2_o_adj_949),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22924),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_4_31_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_4_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_4_31_7 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_4_31_7  (
            .in0(N__17706),
            .in1(N__12334),
            .in2(N__14149),
            .in3(N__14287),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22924),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_4_32_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_4_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_4_32_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_4_32_1  (
            .in0(_gnd_net_),
            .in1(N__17639),
            .in2(_gnd_net_),
            .in3(N__12323),
            .lcout(\c0.rx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22931),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_5 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_5  (
            .in0(N__17158),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i54_LC_4_32_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i54_LC_4_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i54_LC_4_32_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i54_LC_4_32_7  (
            .in0(N__17049),
            .in1(N__12272),
            .in2(_gnd_net_),
            .in3(N__12309),
            .lcout(data_in_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22931),
            .ce(),
            .sr(_gnd_net_));
    defparam i4166_3_lut_LC_5_23_4.C_ON=1'b0;
    defparam i4166_3_lut_LC_5_23_4.SEQ_MODE=4'b0000;
    defparam i4166_3_lut_LC_5_23_4.LUT_INIT=16'b0011001101010101;
    LogicCell40 i4166_3_lut_LC_5_23_4 (
            .in0(N__12248),
            .in1(N__12242),
            .in2(_gnd_net_),
            .in3(N__12236),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_325_326__i1_LC_5_24_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_325_326__i1_LC_5_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_325_326__i1_LC_5_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_325_326__i1_LC_5_24_0  (
            .in0(_gnd_net_),
            .in1(N__15327),
            .in2(N__15495),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter2_0 ),
            .ltout(),
            .carryin(bfn_5_24_0_),
            .carryout(\c0.n3921 ),
            .clk(N__22886),
            .ce(N__12734),
            .sr(N__12743));
    defparam \c0.byte_transmit_counter2_325_326__i2_LC_5_24_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_325_326__i2_LC_5_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_325_326__i2_LC_5_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_325_326__i2_LC_5_24_1  (
            .in0(_gnd_net_),
            .in1(N__15608),
            .in2(_gnd_net_),
            .in3(N__12206),
            .lcout(\c0.byte_transmit_counter2_1 ),
            .ltout(),
            .carryin(\c0.n3921 ),
            .carryout(\c0.n3922 ),
            .clk(N__22886),
            .ce(N__12734),
            .sr(N__12743));
    defparam \c0.byte_transmit_counter2_325_326__i3_LC_5_24_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_325_326__i3_LC_5_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_325_326__i3_LC_5_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_325_326__i3_LC_5_24_2  (
            .in0(_gnd_net_),
            .in1(N__15705),
            .in2(_gnd_net_),
            .in3(N__12746),
            .lcout(\c0.byte_transmit_counter2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22886),
            .ce(N__12734),
            .sr(N__12743));
    defparam \c0.i288_3_lut_4_lut_LC_5_25_0 .C_ON=1'b0;
    defparam \c0.i288_3_lut_4_lut_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i288_3_lut_4_lut_LC_5_25_0 .LUT_INIT=16'b0000010100100111;
    LogicCell40 \c0.i288_3_lut_4_lut_LC_5_25_0  (
            .in0(N__14404),
            .in1(N__12724),
            .in2(N__13100),
            .in3(N__12693),
            .lcout(\c0.n688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i4_LC_5_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i4_LC_5_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i4_LC_5_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i4_LC_5_25_2  (
            .in0(_gnd_net_),
            .in1(N__21520),
            .in2(_gnd_net_),
            .in3(N__19457),
            .lcout(\c0.byte_transmit_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22892),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i7_LC_5_25_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i7_LC_5_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i7_LC_5_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.byte_transmit_counter__i7_LC_5_25_3  (
            .in0(N__21519),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19847),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22892),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i6_LC_5_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i6_LC_5_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i6_LC_5_25_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i6_LC_5_25_4  (
            .in0(_gnd_net_),
            .in1(N__21521),
            .in2(_gnd_net_),
            .in3(N__19379),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22892),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i5_LC_5_25_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i5_LC_5_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i5_LC_5_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.byte_transmit_counter__i5_LC_5_25_5  (
            .in0(N__21518),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19418),
            .lcout(\c0.byte_transmit_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22892),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2421_2_lut_LC_5_25_6 .C_ON=1'b0;
    defparam \c0.i2421_2_lut_LC_5_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2421_2_lut_LC_5_25_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i2421_2_lut_LC_5_25_6  (
            .in0(_gnd_net_),
            .in1(N__12723),
            .in2(_gnd_net_),
            .in3(N__12692),
            .lcout(\c0.n2643 ),
            .ltout(\c0.n2643_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_619_LC_5_25_7 .C_ON=1'b0;
    defparam \c0.tx2_transmit_619_LC_5_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_619_LC_5_25_7 .LUT_INIT=16'b0000100001011101;
    LogicCell40 \c0.tx2_transmit_619_LC_5_25_7  (
            .in0(N__14428),
            .in1(N__15328),
            .in2(N__12704),
            .in3(N__13098),
            .lcout(\c0.tx2_transmit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22892),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_351_LC_5_26_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_351_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_351_LC_5_26_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_351_LC_5_26_0  (
            .in0(N__12665),
            .in1(N__13457),
            .in2(N__12659),
            .in3(N__12965),
            .lcout(),
            .ltout(\c0.n30_adj_892_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2415_4_lut_LC_5_26_1 .C_ON=1'b0;
    defparam \c0.i2415_4_lut_LC_5_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2415_4_lut_LC_5_26_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2415_4_lut_LC_5_26_1  (
            .in0(N__15026),
            .in1(N__12938),
            .in2(N__13109),
            .in3(N__13106),
            .lcout(\c0.n2637 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_5_26_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_5_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_5_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_5_26_2  (
            .in0(N__13075),
            .in1(N__13232),
            .in2(N__13046),
            .in3(N__13004),
            .lcout(),
            .ltout(\c0.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_5_26_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_5_26_3 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i8_4_lut_LC_5_26_3  (
            .in0(N__13571),
            .in1(N__12995),
            .in2(N__12983),
            .in3(N__12980),
            .lcout(\c0.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_348_LC_5_26_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_348_LC_5_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_348_LC_5_26_6 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i10_4_lut_adj_348_LC_5_26_6  (
            .in0(N__12842),
            .in1(N__12959),
            .in2(N__12953),
            .in3(N__15932),
            .lcout(\c0.n26_adj_890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i50_LC_5_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i50_LC_5_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i50_LC_5_27_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i50_LC_5_27_0  (
            .in0(N__15037),
            .in1(N__12928),
            .in2(N__15852),
            .in3(N__14495),
            .lcout(\c0.data_in_frame_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22903),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_326_LC_5_27_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_326_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_326_LC_5_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_326_LC_5_27_1  (
            .in0(N__12914),
            .in1(N__12899),
            .in2(N__14129),
            .in3(N__12866),
            .lcout(\c0.n4391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i42_LC_5_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i42_LC_5_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i42_LC_5_27_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i42_LC_5_27_4  (
            .in0(N__15036),
            .in1(N__14494),
            .in2(N__14177),
            .in3(N__13189),
            .lcout(\c0.data_in_field_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22903),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_342_LC_5_27_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_342_LC_5_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_342_LC_5_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_342_LC_5_27_5  (
            .in0(N__13121),
            .in1(N__12835),
            .in2(N__12794),
            .in3(N__12758),
            .lcout(\c0.n12_adj_887 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i56_LC_5_27_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i56_LC_5_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i56_LC_5_27_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i56_LC_5_27_6  (
            .in0(N__13724),
            .in1(N__16998),
            .in2(_gnd_net_),
            .in3(N__13674),
            .lcout(data_in_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22903),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_319_LC_5_27_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_319_LC_5_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_319_LC_5_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_319_LC_5_27_7  (
            .in0(N__13369),
            .in1(N__13341),
            .in2(N__13652),
            .in3(N__13608),
            .lcout(\c0.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_332_LC_5_28_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_332_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_332_LC_5_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_332_LC_5_28_0  (
            .in0(N__13865),
            .in1(N__13120),
            .in2(N__13565),
            .in3(N__13535),
            .lcout(),
            .ltout(\c0.n4415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_335_LC_5_28_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_335_LC_5_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_335_LC_5_28_1 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i7_4_lut_adj_335_LC_5_28_1  (
            .in0(N__16577),
            .in1(N__13304),
            .in2(N__13499),
            .in3(N__13485),
            .lcout(\c0.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_344_LC_5_28_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_344_LC_5_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_344_LC_5_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_344_LC_5_28_2  (
            .in0(N__13443),
            .in1(N__13406),
            .in2(N__13831),
            .in3(N__13394),
            .lcout(\c0.n4421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_334_LC_5_28_3 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_334_LC_5_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_334_LC_5_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_334_LC_5_28_3  (
            .in0(N__13250),
            .in1(N__13368),
            .in2(N__13298),
            .in3(N__13343),
            .lcout(\c0.n8_adj_883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_301_LC_5_28_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_301_LC_5_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_301_LC_5_28_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_301_LC_5_28_4  (
            .in0(_gnd_net_),
            .in1(N__13293),
            .in2(_gnd_net_),
            .in3(N__13249),
            .lcout(\c0.n4441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_355_LC_5_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_355_LC_5_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_355_LC_5_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_355_LC_5_28_5  (
            .in0(N__13214),
            .in1(N__13182),
            .in2(_gnd_net_),
            .in3(N__13147),
            .lcout(\c0.n4414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i52_LC_5_28_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i52_LC_5_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i52_LC_5_28_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i52_LC_5_28_7  (
            .in0(N__16578),
            .in1(N__17096),
            .in2(_gnd_net_),
            .in3(N__14128),
            .lcout(data_in_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22911),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i55_LC_5_29_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i55_LC_5_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i55_LC_5_29_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i55_LC_5_29_0  (
            .in0(N__16986),
            .in1(N__13928),
            .in2(_gnd_net_),
            .in3(N__14090),
            .lcout(data_in_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22918),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i41_LC_5_29_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i41_LC_5_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i41_LC_5_29_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i41_LC_5_29_1  (
            .in0(N__16086),
            .in1(N__14271),
            .in2(_gnd_net_),
            .in3(N__16988),
            .lcout(data_in_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22918),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_5_29_2 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_5_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_5_29_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_5_29_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14056),
            .lcout(tx2_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_328_LC_5_29_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_328_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_328_LC_5_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_328_LC_5_29_3  (
            .in0(N__14013),
            .in1(N__13964),
            .in2(N__13935),
            .in3(N__13896),
            .lcout(\c0.n12_adj_878 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i61_LC_5_29_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i61_LC_5_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i61_LC_5_29_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i61_LC_5_29_4  (
            .in0(N__16987),
            .in1(N__13856),
            .in2(_gnd_net_),
            .in3(N__13820),
            .lcout(data_in_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22918),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i24_LC_5_29_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i24_LC_5_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i24_LC_5_29_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i24_LC_5_29_5  (
            .in0(N__13796),
            .in1(N__15045),
            .in2(N__14685),
            .in3(N__13751),
            .lcout(\c0.data_in_field_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22918),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i36_LC_5_29_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i36_LC_5_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i36_LC_5_29_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i36_LC_5_29_6  (
            .in0(N__16985),
            .in1(N__16561),
            .in2(_gnd_net_),
            .in3(N__14226),
            .lcout(data_in_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22918),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i10_LC_5_29_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i10_LC_5_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i10_LC_5_29_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i10_LC_5_29_7  (
            .in0(N__15080),
            .in1(N__15044),
            .in2(N__14684),
            .in3(N__14310),
            .lcout(\c0.data_in_field_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22918),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i50_LC_5_30_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i50_LC_5_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i50_LC_5_30_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i50_LC_5_30_0  (
            .in0(N__17265),
            .in1(N__16973),
            .in2(_gnd_net_),
            .in3(N__16752),
            .lcout(data_in_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22925),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2429_2_lut_LC_5_30_1 .C_ON=1'b0;
    defparam \c0.rx.i2429_2_lut_LC_5_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2429_2_lut_LC_5_30_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i2429_2_lut_LC_5_30_1  (
            .in0(_gnd_net_),
            .in1(N__16360),
            .in2(_gnd_net_),
            .in3(N__16393),
            .lcout(n2651),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_5_30_2 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_5_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_5_30_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_5_30_2  (
            .in0(N__16032),
            .in1(N__16158),
            .in2(_gnd_net_),
            .in3(N__16143),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22925),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_5_30_3 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_5_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_5_30_3 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_5_30_3  (
            .in0(N__16144),
            .in1(N__16361),
            .in2(N__16163),
            .in3(N__16033),
            .lcout(\c0.rx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22925),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i33_LC_5_30_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i33_LC_5_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i33_LC_5_30_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i33_LC_5_30_4  (
            .in0(N__17097),
            .in1(N__14272),
            .in2(_gnd_net_),
            .in3(N__14247),
            .lcout(data_in_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22925),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i28_LC_5_30_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i28_LC_5_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i28_LC_5_30_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i28_LC_5_30_5  (
            .in0(N__16971),
            .in1(N__14227),
            .in2(_gnd_net_),
            .in3(N__14201),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22925),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_5_30_6 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_5_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_5_30_6 .LUT_INIT=16'b0110101000000000;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_5_30_6  (
            .in0(N__16394),
            .in1(N__16162),
            .in2(N__16004),
            .in3(N__16145),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22925),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i43_LC_5_30_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i43_LC_5_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i43_LC_5_30_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i43_LC_5_30_7  (
            .in0(N__16972),
            .in1(N__14161),
            .in2(_gnd_net_),
            .in3(N__15854),
            .lcout(data_in_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22925),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_LC_5_31_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_LC_5_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_LC_5_31_0 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_LC_5_31_0  (
            .in0(N__15119),
            .in1(N__17557),
            .in2(N__16034),
            .in3(N__17637),
            .lcout(n1222),
            .ltout(n1222_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_5_31_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_5_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_5_31_1 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_5_31_1  (
            .in0(N__15154),
            .in1(N__16327),
            .in2(N__15158),
            .in3(N__17709),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22932),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_27_i4_2_lut_LC_5_31_2 .C_ON=1'b0;
    defparam \c0.rx.equal_27_i4_2_lut_LC_5_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_27_i4_2_lut_LC_5_31_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.rx.equal_27_i4_2_lut_LC_5_31_2  (
            .in0(N__16396),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16363),
            .lcout(n4_adj_950),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_25_i4_2_lut_LC_5_31_3 .C_ON=1'b0;
    defparam \c0.rx.equal_25_i4_2_lut_LC_5_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_25_i4_2_lut_LC_5_31_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.equal_25_i4_2_lut_LC_5_31_3  (
            .in0(_gnd_net_),
            .in1(N__16362),
            .in2(_gnd_net_),
            .in3(N__16395),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_5_31_5 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_5_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_5_31_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.i1_2_lut_LC_5_31_5  (
            .in0(_gnd_net_),
            .in1(N__17756),
            .in2(_gnd_net_),
            .in3(N__17372),
            .lcout(\c0.rx.n2269 ),
            .ltout(\c0.rx.n2269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_adj_279_LC_5_31_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_adj_279_LC_5_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_adj_279_LC_5_31_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_adj_279_LC_5_31_6  (
            .in0(N__16031),
            .in1(N__17558),
            .in2(N__15113),
            .in3(N__17638),
            .lcout(n1227),
            .ltout(n1227_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_31_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_31_7 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_5_31_7  (
            .in0(N__17287),
            .in1(N__16328),
            .in2(N__15092),
            .in3(N__17710),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22932),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_5_32_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_5_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_5_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_2_lut_LC_5_32_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16226),
            .in3(N__15089),
            .lcout(n226),
            .ltout(),
            .carryin(bfn_5_32_0_),
            .carryout(\c0.rx.n3884 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_3_lut_LC_5_32_1 .C_ON=1'b1;
    defparam \c0.rx.add_62_3_lut_LC_5_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_3_lut_LC_5_32_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_3_lut_LC_5_32_1  (
            .in0(N__16517),
            .in1(N__16306),
            .in2(_gnd_net_),
            .in3(N__15086),
            .lcout(\c0.rx.n4679 ),
            .ltout(),
            .carryin(\c0.rx.n3884 ),
            .carryout(\c0.rx.n3885 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_4_lut_LC_5_32_2 .C_ON=1'b1;
    defparam \c0.rx.add_62_4_lut_LC_5_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_4_lut_LC_5_32_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_4_lut_LC_5_32_2  (
            .in0(_gnd_net_),
            .in1(N__17423),
            .in2(_gnd_net_),
            .in3(N__15083),
            .lcout(n224),
            .ltout(),
            .carryin(\c0.rx.n3885 ),
            .carryout(\c0.rx.n3886 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_5_lut_LC_5_32_3 .C_ON=1'b1;
    defparam \c0.rx.add_62_5_lut_LC_5_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_5_lut_LC_5_32_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_5_lut_LC_5_32_3  (
            .in0(_gnd_net_),
            .in1(N__16428),
            .in2(_gnd_net_),
            .in3(N__15260),
            .lcout(n223),
            .ltout(),
            .carryin(\c0.rx.n3886 ),
            .carryout(\c0.rx.n3887 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_6_lut_LC_5_32_4 .C_ON=1'b1;
    defparam \c0.rx.add_62_6_lut_LC_5_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_6_lut_LC_5_32_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_6_lut_LC_5_32_4  (
            .in0(_gnd_net_),
            .in1(N__16180),
            .in2(_gnd_net_),
            .in3(N__15257),
            .lcout(n222),
            .ltout(),
            .carryin(\c0.rx.n3887 ),
            .carryout(\c0.rx.n3888 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_7_lut_LC_5_32_5 .C_ON=1'b1;
    defparam \c0.rx.add_62_7_lut_LC_5_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_7_lut_LC_5_32_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_7_lut_LC_5_32_5  (
            .in0(_gnd_net_),
            .in1(N__16474),
            .in2(_gnd_net_),
            .in3(N__15254),
            .lcout(n221),
            .ltout(),
            .carryin(\c0.rx.n3888 ),
            .carryout(\c0.rx.n3889 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_8_lut_LC_5_32_6 .C_ON=1'b1;
    defparam \c0.rx.add_62_8_lut_LC_5_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_8_lut_LC_5_32_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_8_lut_LC_5_32_6  (
            .in0(_gnd_net_),
            .in1(N__17855),
            .in2(_gnd_net_),
            .in3(N__15251),
            .lcout(n220),
            .ltout(),
            .carryin(\c0.rx.n3889 ),
            .carryout(\c0.rx.n3890 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_9_lut_LC_5_32_7 .C_ON=1'b0;
    defparam \c0.rx.add_62_9_lut_LC_5_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_9_lut_LC_5_32_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_9_lut_LC_5_32_7  (
            .in0(_gnd_net_),
            .in1(N__16273),
            .in2(_gnd_net_),
            .in3(N__15248),
            .lcout(n219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i1_LC_6_23_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i1_LC_6_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i1_LC_6_23_0 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.data_out_0__i1_LC_6_23_0  (
            .in0(N__22427),
            .in1(N__21540),
            .in2(_gnd_net_),
            .in3(N__21257),
            .lcout(data_out_field_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22887),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i6_LC_6_23_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i6_LC_6_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i6_LC_6_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i6_LC_6_23_4  (
            .in0(_gnd_net_),
            .in1(N__15245),
            .in2(_gnd_net_),
            .in3(N__15233),
            .lcout(\c0.tx2.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22887),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i0_LC_6_25_0 .C_ON=1'b1;
    defparam \c0.data_327__i0_LC_6_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i0_LC_6_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i0_LC_6_25_0  (
            .in0(_gnd_net_),
            .in1(N__18277),
            .in2(_gnd_net_),
            .in3(N__15164),
            .lcout(\c0.data_0 ),
            .ltout(),
            .carryin(bfn_6_25_0_),
            .carryout(\c0.n3906 ),
            .clk(N__22897),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i1_LC_6_25_1 .C_ON=1'b1;
    defparam \c0.data_327__i1_LC_6_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i1_LC_6_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i1_LC_6_25_1  (
            .in0(_gnd_net_),
            .in1(N__15898),
            .in2(_gnd_net_),
            .in3(N__15161),
            .lcout(\c0.data_1 ),
            .ltout(),
            .carryin(\c0.n3906 ),
            .carryout(\c0.n3907 ),
            .clk(N__22897),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i2_LC_6_25_2 .C_ON=1'b1;
    defparam \c0.data_327__i2_LC_6_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i2_LC_6_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i2_LC_6_25_2  (
            .in0(_gnd_net_),
            .in1(N__19060),
            .in2(_gnd_net_),
            .in3(N__15287),
            .lcout(\c0.data_2 ),
            .ltout(),
            .carryin(\c0.n3907 ),
            .carryout(\c0.n3908 ),
            .clk(N__22897),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i3_LC_6_25_3 .C_ON=1'b1;
    defparam \c0.data_327__i3_LC_6_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i3_LC_6_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i3_LC_6_25_3  (
            .in0(_gnd_net_),
            .in1(N__18613),
            .in2(_gnd_net_),
            .in3(N__15284),
            .lcout(\c0.data_3 ),
            .ltout(),
            .carryin(\c0.n3908 ),
            .carryout(\c0.n3909 ),
            .clk(N__22897),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i4_LC_6_25_4 .C_ON=1'b1;
    defparam \c0.data_327__i4_LC_6_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i4_LC_6_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i4_LC_6_25_4  (
            .in0(_gnd_net_),
            .in1(N__18658),
            .in2(_gnd_net_),
            .in3(N__15281),
            .lcout(\c0.data_4 ),
            .ltout(),
            .carryin(\c0.n3909 ),
            .carryout(\c0.n3910 ),
            .clk(N__22897),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i5_LC_6_25_5 .C_ON=1'b1;
    defparam \c0.data_327__i5_LC_6_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i5_LC_6_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i5_LC_6_25_5  (
            .in0(_gnd_net_),
            .in1(N__18814),
            .in2(_gnd_net_),
            .in3(N__15278),
            .lcout(\c0.data_5 ),
            .ltout(),
            .carryin(\c0.n3910 ),
            .carryout(\c0.n3911 ),
            .clk(N__22897),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i6_LC_6_25_6 .C_ON=1'b1;
    defparam \c0.data_327__i6_LC_6_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i6_LC_6_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i6_LC_6_25_6  (
            .in0(_gnd_net_),
            .in1(N__18106),
            .in2(_gnd_net_),
            .in3(N__15275),
            .lcout(\c0.data_6 ),
            .ltout(),
            .carryin(\c0.n3911 ),
            .carryout(\c0.n3912 ),
            .clk(N__22897),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i7_LC_6_25_7 .C_ON=1'b1;
    defparam \c0.data_327__i7_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i7_LC_6_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i7_LC_6_25_7  (
            .in0(_gnd_net_),
            .in1(N__18088),
            .in2(_gnd_net_),
            .in3(N__15272),
            .lcout(\c0.data_7 ),
            .ltout(),
            .carryin(\c0.n3912 ),
            .carryout(\c0.n3913 ),
            .clk(N__22897),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i8_LC_6_26_0 .C_ON=1'b1;
    defparam \c0.data_327__i8_LC_6_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i8_LC_6_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i8_LC_6_26_0  (
            .in0(_gnd_net_),
            .in1(N__18028),
            .in2(_gnd_net_),
            .in3(N__15269),
            .lcout(\c0.data_8 ),
            .ltout(),
            .carryin(bfn_6_26_0_),
            .carryout(\c0.n3914 ),
            .clk(N__22904),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i9_LC_6_26_1 .C_ON=1'b1;
    defparam \c0.data_327__i9_LC_6_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i9_LC_6_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i9_LC_6_26_1  (
            .in0(_gnd_net_),
            .in1(N__15301),
            .in2(_gnd_net_),
            .in3(N__15266),
            .lcout(\c0.data_9 ),
            .ltout(),
            .carryin(\c0.n3914 ),
            .carryout(\c0.n3915 ),
            .clk(N__22904),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i10_LC_6_26_2 .C_ON=1'b1;
    defparam \c0.data_327__i10_LC_6_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i10_LC_6_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i10_LC_6_26_2  (
            .in0(_gnd_net_),
            .in1(N__18184),
            .in2(_gnd_net_),
            .in3(N__15263),
            .lcout(\c0.data_10 ),
            .ltout(),
            .carryin(\c0.n3915 ),
            .carryout(\c0.n3916 ),
            .clk(N__22904),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i11_LC_6_26_3 .C_ON=1'b1;
    defparam \c0.data_327__i11_LC_6_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i11_LC_6_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i11_LC_6_26_3  (
            .in0(_gnd_net_),
            .in1(N__18634),
            .in2(_gnd_net_),
            .in3(N__15803),
            .lcout(\c0.data_11 ),
            .ltout(),
            .carryin(\c0.n3916 ),
            .carryout(\c0.n3917 ),
            .clk(N__22904),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i12_LC_6_26_4 .C_ON=1'b1;
    defparam \c0.data_327__i12_LC_6_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i12_LC_6_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i12_LC_6_26_4  (
            .in0(_gnd_net_),
            .in1(N__19297),
            .in2(_gnd_net_),
            .in3(N__15800),
            .lcout(\c0.data_12 ),
            .ltout(),
            .carryin(\c0.n3917 ),
            .carryout(\c0.n3918 ),
            .clk(N__22904),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i13_LC_6_26_5 .C_ON=1'b1;
    defparam \c0.data_327__i13_LC_6_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i13_LC_6_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i13_LC_6_26_5  (
            .in0(_gnd_net_),
            .in1(N__21619),
            .in2(_gnd_net_),
            .in3(N__15797),
            .lcout(\c0.data_13 ),
            .ltout(),
            .carryin(\c0.n3918 ),
            .carryout(\c0.n3919 ),
            .clk(N__22904),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i14_LC_6_26_6 .C_ON=1'b1;
    defparam \c0.data_327__i14_LC_6_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i14_LC_6_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i14_LC_6_26_6  (
            .in0(_gnd_net_),
            .in1(N__18067),
            .in2(_gnd_net_),
            .in3(N__15794),
            .lcout(\c0.data_14 ),
            .ltout(),
            .carryin(\c0.n3919 ),
            .carryout(\c0.n3920 ),
            .clk(N__22904),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_327__i15_LC_6_26_7 .C_ON=1'b0;
    defparam \c0.data_327__i15_LC_6_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_327__i15_LC_6_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_327__i15_LC_6_26_7  (
            .in0(_gnd_net_),
            .in1(N__17977),
            .in2(_gnd_net_),
            .in3(N__15791),
            .lcout(\c0.data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22904),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4401_3_lut_LC_6_27_1 .C_ON=1'b0;
    defparam \c0.i4401_3_lut_LC_6_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4401_3_lut_LC_6_27_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \c0.i4401_3_lut_LC_6_27_1  (
            .in0(N__15767),
            .in1(N__15637),
            .in2(_gnd_net_),
            .in3(N__15527),
            .lcout(\c0.FRAME_MATCHER_wait_for_transmission_N_423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i34_LC_6_27_2 .C_ON=1'b0;
    defparam \c0.data_out_0__i34_LC_6_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i34_LC_6_27_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0__i34_LC_6_27_2  (
            .in0(N__18894),
            .in1(N__21562),
            .in2(N__15305),
            .in3(N__21255),
            .lcout(\c0.data_out_field_47_N_682_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22912),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4264_3_lut_LC_6_27_3 .C_ON=1'b0;
    defparam \c0.i4264_3_lut_LC_6_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4264_3_lut_LC_6_27_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4264_3_lut_LC_6_27_3  (
            .in0(N__18383),
            .in1(N__20288),
            .in2(_gnd_net_),
            .in3(N__20551),
            .lcout(),
            .ltout(\c0.n4619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4435_LC_6_27_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4435_LC_6_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4435_LC_6_27_4 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_4435_LC_6_27_4  (
            .in0(N__20783),
            .in1(N__20693),
            .in2(N__15290),
            .in3(N__19565),
            .lcout(\c0.n4789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_6_27_5 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_6_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_6_27_5 .LUT_INIT=16'b0011010000110000;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_6_27_5  (
            .in0(N__23249),
            .in1(N__21852),
            .in2(N__19210),
            .in3(N__23207),
            .lcout(\c0.tx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22912),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_318_LC_6_27_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_318_LC_6_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_318_LC_6_27_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_318_LC_6_27_6  (
            .in0(N__18558),
            .in1(N__18172),
            .in2(_gnd_net_),
            .in3(N__18888),
            .lcout(\c0.n4380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i42_LC_6_27_7 .C_ON=1'b0;
    defparam \c0.data_out_0__i42_LC_6_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i42_LC_6_27_7 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0__i42_LC_6_27_7  (
            .in0(N__21256),
            .in1(N__18585),
            .in2(N__15905),
            .in3(N__21554),
            .lcout(\c0.data_out_field_47_N_682_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22912),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i51_LC_6_28_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i51_LC_6_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i51_LC_6_28_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i51_LC_6_28_0  (
            .in0(N__16997),
            .in1(N__15845),
            .in2(_gnd_net_),
            .in3(N__15887),
            .lcout(data_in_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22919),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4162_3_lut_LC_6_28_2 .C_ON=1'b0;
    defparam \c0.i4162_3_lut_LC_6_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4162_3_lut_LC_6_28_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4162_3_lut_LC_6_28_2  (
            .in0(N__20550),
            .in1(N__18137),
            .in2(_gnd_net_),
            .in3(N__18233),
            .lcout(),
            .ltout(\c0.n4517_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_6_28_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_6_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_6_28_3 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_6_28_3  (
            .in0(N__19589),
            .in1(N__15917),
            .in2(N__15818),
            .in3(N__20706),
            .lcout(),
            .ltout(\c0.n4867_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4867_bdd_4_lut_LC_6_28_4 .C_ON=1'b0;
    defparam \c0.n4867_bdd_4_lut_LC_6_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.n4867_bdd_4_lut_LC_6_28_4 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n4867_bdd_4_lut_LC_6_28_4  (
            .in0(N__15809),
            .in1(N__18395),
            .in2(N__15815),
            .in3(N__19590),
            .lcout(),
            .ltout(tx_data_2_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_6_28_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_6_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_6_28_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_6_28_5  (
            .in0(_gnd_net_),
            .in1(N__22116),
            .in2(N__15812),
            .in3(N__17191),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22919),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4209_3_lut_LC_6_28_6 .C_ON=1'b0;
    defparam \c0.i4209_3_lut_LC_6_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4209_3_lut_LC_6_28_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4209_3_lut_LC_6_28_6  (
            .in0(N__20549),
            .in1(N__22001),
            .in2(_gnd_net_),
            .in3(N__21680),
            .lcout(\c0.n4564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_327_LC_6_29_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_327_LC_6_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_327_LC_6_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_327_LC_6_29_0  (
            .in0(N__16087),
            .in1(N__15962),
            .in2(_gnd_net_),
            .in3(N__15950),
            .lcout(\c0.n4409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4354_2_lut_LC_6_29_1 .C_ON=1'b0;
    defparam \c0.rx.i4354_2_lut_LC_6_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4354_2_lut_LC_6_29_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.i4354_2_lut_LC_6_29_1  (
            .in0(N__17363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17618),
            .lcout(\c0.rx.n4677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_LC_6_29_2 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_LC_6_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_LC_6_29_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i2_2_lut_LC_6_29_2  (
            .in0(N__16225),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17856),
            .lcout(\c0.rx.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i223_3_lut_LC_6_29_3 .C_ON=1'b0;
    defparam \c0.rx.i223_3_lut_LC_6_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i223_3_lut_LC_6_29_3 .LUT_INIT=16'b1100100011001000;
    LogicCell40 \c0.rx.i223_3_lut_LC_6_29_3  (
            .in0(N__17419),
            .in1(N__16430),
            .in2(N__16310),
            .in3(_gnd_net_),
            .lcout(\c0.rx.n232 ),
            .ltout(\c0.rx.n232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_6_29_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_6_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_6_29_4 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_6_29_4  (
            .in0(N__15977),
            .in1(N__17857),
            .in2(N__15920),
            .in3(N__16277),
            .lcout(\c0.rx.r_SM_Main_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22926),
            .ce(),
            .sr(N__17330));
    defparam \c0.i4161_3_lut_LC_6_29_5 .C_ON=1'b0;
    defparam \c0.i4161_3_lut_LC_6_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4161_3_lut_LC_6_29_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4161_3_lut_LC_6_29_5  (
            .in0(N__20341),
            .in1(N__18563),
            .in2(_gnd_net_),
            .in3(N__20519),
            .lcout(\c0.n4516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4171_3_lut_LC_6_29_7 .C_ON=1'b0;
    defparam \c0.i4171_3_lut_LC_6_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4171_3_lut_LC_6_29_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i4171_3_lut_LC_6_29_7  (
            .in0(N__18173),
            .in1(N__19772),
            .in2(_gnd_net_),
            .in3(N__20518),
            .lcout(\c0.n4526 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13_4_lut_4_lut_LC_6_30_0 .C_ON=1'b0;
    defparam \c0.rx.i13_4_lut_4_lut_LC_6_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13_4_lut_4_lut_LC_6_30_0 .LUT_INIT=16'b0010010100000101;
    LogicCell40 \c0.rx.i13_4_lut_4_lut_LC_6_30_0  (
            .in0(N__17553),
            .in1(N__17620),
            .in2(N__17789),
            .in3(N__17368),
            .lcout(),
            .ltout(\c0.rx.n1464_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_6_30_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_6_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_6_30_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_6_30_1  (
            .in0(N__17621),
            .in1(N__16906),
            .in2(N__15908),
            .in3(N__17554),
            .lcout(rx_data_ready_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22933),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_4_lut_LC_6_30_2 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_4_lut_LC_6_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_4_lut_LC_6_30_2 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \c0.rx.i2_4_lut_4_lut_LC_6_30_2  (
            .in0(N__17551),
            .in1(N__17619),
            .in2(N__17788),
            .in3(N__17367),
            .lcout(n1527),
            .ltout(n1527_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_3_lut_4_lut_LC_6_30_3 .C_ON=1'b0;
    defparam \c0.rx.i1_3_lut_4_lut_LC_6_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_3_lut_4_lut_LC_6_30_3 .LUT_INIT=16'b0111111100001111;
    LogicCell40 \c0.rx.i1_3_lut_4_lut_LC_6_30_3  (
            .in0(N__16392),
            .in1(N__16000),
            .in2(N__16148),
            .in3(N__17552),
            .lcout(n2142),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i49_LC_6_30_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i49_LC_6_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i49_LC_6_30_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i49_LC_6_30_4  (
            .in0(N__16905),
            .in1(N__16085),
            .in2(_gnd_net_),
            .in3(N__16131),
            .lcout(data_in_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22933),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_276_LC_6_30_5 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_276_LC_6_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_276_LC_6_30_5 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.rx.i1_4_lut_adj_276_LC_6_30_5  (
            .in0(N__17858),
            .in1(N__15973),
            .in2(N__16058),
            .in3(N__16272),
            .lcout(\c0.rx.r_SM_Main_2_N_816_2 ),
            .ltout(\c0.rx.r_SM_Main_2_N_816_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4336_2_lut_3_lut_4_lut_LC_6_30_6 .C_ON=1'b0;
    defparam \c0.rx.i4336_2_lut_3_lut_4_lut_LC_6_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4336_2_lut_3_lut_4_lut_LC_6_30_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i4336_2_lut_3_lut_4_lut_LC_6_30_6  (
            .in0(N__16358),
            .in1(N__16026),
            .in2(N__16049),
            .in3(N__16391),
            .lcout(\c0.rx.n4678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_274_LC_6_30_7 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_274_LC_6_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_274_LC_6_30_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_274_LC_6_30_7  (
            .in0(N__16027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16359),
            .lcout(n4_adj_943),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i3_LC_6_31_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i3_LC_6_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_6_31_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_6_31_0  (
            .in0(N__16429),
            .in1(N__17925),
            .in2(N__15989),
            .in3(N__17888),
            .lcout(r_Clock_Count_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_289_LC_6_31_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_289_LC_6_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_289_LC_6_31_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_289_LC_6_31_1  (
            .in0(_gnd_net_),
            .in1(N__18562),
            .in2(_gnd_net_),
            .in3(N__20198),
            .lcout(n4_adj_942),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_275_LC_6_31_2 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_275_LC_6_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_275_LC_6_31_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_adj_275_LC_6_31_2  (
            .in0(_gnd_net_),
            .in1(N__16473),
            .in2(_gnd_net_),
            .in3(N__16179),
            .lcout(\c0.rx.n214 ),
            .ltout(\c0.rx.n214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_268_LC_6_31_3 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_268_LC_6_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_268_LC_6_31_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.i1_4_lut_adj_268_LC_6_31_3  (
            .in0(N__16424),
            .in1(N__16270),
            .in2(N__16403),
            .in3(N__16304),
            .lcout(\c0.rx.n4 ),
            .ltout(\c0.rx.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_LC_6_31_4 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_LC_6_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_LC_6_31_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_LC_6_31_4  (
            .in0(N__17837),
            .in1(N__16217),
            .in2(N__16400),
            .in3(N__17416),
            .lcout(\c0.rx.n2179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_28_i4_2_lut_LC_6_31_5 .C_ON=1'b0;
    defparam \c0.rx.equal_28_i4_2_lut_LC_6_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_28_i4_2_lut_LC_6_31_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.equal_28_i4_2_lut_LC_6_31_5  (
            .in0(N__16397),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16364),
            .lcout(n4_adj_951),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_6_31_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i1_LC_6_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_6_31_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_6_31_6  (
            .in0(N__16305),
            .in1(N__16316),
            .in2(_gnd_net_),
            .in3(N__17924),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i7_LC_6_31_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_6_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_6_31_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_6_31_7  (
            .in0(N__17889),
            .in1(N__16283),
            .in2(N__17933),
            .in3(N__16271),
            .lcout(r_Clock_Count_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2038_4_lut_LC_6_32_0 .C_ON=1'b0;
    defparam \c0.rx.i2038_4_lut_LC_6_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2038_4_lut_LC_6_32_0 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \c0.rx.i2038_4_lut_LC_6_32_0  (
            .in0(N__17306),
            .in1(N__16247),
            .in2(N__17550),
            .in3(N__16490),
            .lcout(n573),
            .ltout(n573_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_6_32_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_6_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_6_32_1 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_6_32_1  (
            .in0(N__16238),
            .in1(N__16224),
            .in2(N__16229),
            .in3(N__17929),
            .lcout(r_Clock_Count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22944),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i4_LC_6_32_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i4_LC_6_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_6_32_2 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_6_32_2  (
            .in0(N__17930),
            .in1(N__16184),
            .in2(N__16196),
            .in3(N__17886),
            .lcout(r_Clock_Count_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22944),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4353_3_lut_LC_6_32_3 .C_ON=1'b0;
    defparam \c0.rx.i4353_3_lut_LC_6_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4353_3_lut_LC_6_32_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.rx.i4353_3_lut_LC_6_32_3  (
            .in0(N__17766),
            .in1(N__17685),
            .in2(_gnd_net_),
            .in3(N__17809),
            .lcout(),
            .ltout(\c0.rx.n4641_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_269_LC_6_32_4 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_269_LC_6_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_269_LC_6_32_4 .LUT_INIT=16'b1101110011111110;
    LogicCell40 \c0.rx.i1_4_lut_adj_269_LC_6_32_4  (
            .in0(N__17524),
            .in1(N__17632),
            .in2(N__16520),
            .in3(N__17374),
            .lcout(\c0.rx.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4_4_lut_LC_6_32_5 .C_ON=1'b0;
    defparam \c0.rx.i4_4_lut_LC_6_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4_4_lut_LC_6_32_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \c0.rx.i4_4_lut_LC_6_32_5  (
            .in0(N__16511),
            .in1(N__17417),
            .in2(N__16505),
            .in3(N__17304),
            .lcout(\c0.rx.n4093 ),
            .ltout(\c0.rx.n4093_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i82_3_lut_4_lut_LC_6_32_6 .C_ON=1'b0;
    defparam \c0.rx.i82_3_lut_4_lut_LC_6_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i82_3_lut_4_lut_LC_6_32_6 .LUT_INIT=16'b0101010111010001;
    LogicCell40 \c0.rx.i82_3_lut_4_lut_LC_6_32_6  (
            .in0(N__17305),
            .in1(N__17767),
            .in2(N__16493),
            .in3(N__17631),
            .lcout(\c0.rx.n2246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i5_LC_6_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i5_LC_6_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_6_32_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_6_32_7  (
            .in0(N__17887),
            .in1(N__17931),
            .in2(N__16484),
            .in3(N__16475),
            .lcout(r_Clock_Count_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22944),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i25_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i25_LC_7_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i25_LC_7_24_0 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.data_out_0__i25_LC_7_24_0  (
            .in0(N__21525),
            .in1(N__18314),
            .in2(_gnd_net_),
            .in3(N__21249),
            .lcout(data_out_field_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22898),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4430_LC_7_25_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4430_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4430_LC_7_25_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_4430_LC_7_25_1  (
            .in0(N__16607),
            .in1(N__19602),
            .in2(N__16439),
            .in3(N__20705),
            .lcout(),
            .ltout(\c0.n4783_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4783_bdd_4_lut_LC_7_25_2 .C_ON=1'b0;
    defparam \c0.n4783_bdd_4_lut_LC_7_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.n4783_bdd_4_lut_LC_7_25_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n4783_bdd_4_lut_LC_7_25_2  (
            .in0(N__19603),
            .in1(N__16601),
            .in2(N__16457),
            .in3(N__16454),
            .lcout(),
            .ltout(tx_data_3_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_7_25_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_7_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_7_25_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_7_25_3  (
            .in0(_gnd_net_),
            .in1(N__22151),
            .in2(N__16442),
            .in3(N__17206),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22905),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4267_3_lut_LC_7_26_0 .C_ON=1'b0;
    defparam \c0.i4267_3_lut_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4267_3_lut_LC_7_26_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4267_3_lut_LC_7_26_0  (
            .in0(N__20546),
            .in1(N__18056),
            .in2(_gnd_net_),
            .in3(N__18793),
            .lcout(\c0.n4622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4266_3_lut_LC_7_26_1 .C_ON=1'b0;
    defparam \c0.i4266_3_lut_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4266_3_lut_LC_7_26_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4266_3_lut_LC_7_26_1  (
            .in0(N__21957),
            .in1(N__19822),
            .in2(_gnd_net_),
            .in3(N__20547),
            .lcout(\c0.n4621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4170_3_lut_LC_7_26_2 .C_ON=1'b0;
    defparam \c0.i4170_3_lut_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4170_3_lut_LC_7_26_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4170_3_lut_LC_7_26_2  (
            .in0(N__20548),
            .in1(N__18479),
            .in2(_gnd_net_),
            .in3(N__18364),
            .lcout(\c0.n4525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i44_LC_7_26_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i44_LC_7_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i44_LC_7_26_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i44_LC_7_26_3  (
            .in0(N__16548),
            .in1(N__17092),
            .in2(_gnd_net_),
            .in3(N__16591),
            .lcout(data_in_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22913),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4765_bdd_4_lut_LC_7_26_4 .C_ON=1'b0;
    defparam \c0.n4765_bdd_4_lut_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.n4765_bdd_4_lut_LC_7_26_4 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \c0.n4765_bdd_4_lut_LC_7_26_4  (
            .in0(N__20369),
            .in1(N__19286),
            .in2(N__21931),
            .in3(N__20708),
            .lcout(),
            .ltout(\c0.n4768_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i277446_i1_3_lut_LC_7_26_5 .C_ON=1'b0;
    defparam \c0.i277446_i1_3_lut_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i277446_i1_3_lut_LC_7_26_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.i277446_i1_3_lut_LC_7_26_5  (
            .in0(_gnd_net_),
            .in1(N__17963),
            .in2(N__16532),
            .in3(N__19585),
            .lcout(),
            .ltout(tx_data_7_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_7_26_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_7_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_7_26_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_7_26_6  (
            .in0(_gnd_net_),
            .in1(N__22150),
            .in2(N__16529),
            .in3(N__16658),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22913),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4488_LC_7_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4488_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4488_LC_7_27_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_4488_LC_7_27_0  (
            .in0(N__16646),
            .in1(N__19566),
            .in2(N__16625),
            .in3(N__20694),
            .lcout(),
            .ltout(\c0.n4843_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4843_bdd_4_lut_LC_7_27_1 .C_ON=1'b0;
    defparam \c0.n4843_bdd_4_lut_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n4843_bdd_4_lut_LC_7_27_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n4843_bdd_4_lut_LC_7_27_1  (
            .in0(N__19567),
            .in1(N__19082),
            .in2(N__16526),
            .in3(N__18245),
            .lcout(),
            .ltout(tx_data_1_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_7_27_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_7_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_7_27_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_7_27_2  (
            .in0(_gnd_net_),
            .in1(N__22141),
            .in2(N__16523),
            .in3(N__17236),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22920),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4234_3_lut_LC_7_27_3 .C_ON=1'b0;
    defparam \c0.tx.i4234_3_lut_LC_7_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4234_3_lut_LC_7_27_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.i4234_3_lut_LC_7_27_3  (
            .in0(N__19185),
            .in1(N__16657),
            .in2(_gnd_net_),
            .in3(N__16639),
            .lcout(\c0.tx.n4589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4230_3_lut_LC_7_27_4 .C_ON=1'b0;
    defparam \c0.i4230_3_lut_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4230_3_lut_LC_7_27_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i4230_3_lut_LC_7_27_4  (
            .in0(N__18887),
            .in1(N__18584),
            .in2(_gnd_net_),
            .in3(N__20554),
            .lcout(\c0.n4585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1361_2_lut_LC_7_27_5 .C_ON=1'b0;
    defparam \c0.tx.i1361_2_lut_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1361_2_lut_LC_7_27_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.tx.i1361_2_lut_LC_7_27_5  (
            .in0(N__23244),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23205),
            .lcout(\c0.tx.n1588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_7_27_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_7_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_7_27_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_7_27_6  (
            .in0(N__16640),
            .in1(N__22142),
            .in2(_gnd_net_),
            .in3(N__19334),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22920),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4493_LC_7_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4493_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4493_LC_7_28_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_4493_LC_7_28_0  (
            .in0(N__16712),
            .in1(N__19596),
            .in2(N__19676),
            .in3(N__20701),
            .lcout(),
            .ltout(\c0.n4861_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4861_bdd_4_lut_LC_7_28_1 .C_ON=1'b0;
    defparam \c0.n4861_bdd_4_lut_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.n4861_bdd_4_lut_LC_7_28_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n4861_bdd_4_lut_LC_7_28_1  (
            .in0(N__19597),
            .in1(N__16616),
            .in2(N__16631),
            .in3(N__18200),
            .lcout(),
            .ltout(tx_data_0_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_7_28_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_7_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_7_28_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_7_28_2  (
            .in0(_gnd_net_),
            .in1(N__22114),
            .in2(N__16628),
            .in3(N__17221),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22927),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4231_3_lut_LC_7_28_3 .C_ON=1'b0;
    defparam \c0.i4231_3_lut_LC_7_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4231_3_lut_LC_7_28_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4231_3_lut_LC_7_28_3  (
            .in0(N__18214),
            .in1(N__17999),
            .in2(_gnd_net_),
            .in3(N__20553),
            .lcout(\c0.n4586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4233_3_lut_LC_7_28_4 .C_ON=1'b0;
    defparam \c0.tx.i4233_3_lut_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4233_3_lut_LC_7_28_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.i4233_3_lut_LC_7_28_4  (
            .in0(N__19199),
            .in1(N__16687),
            .in2(_gnd_net_),
            .in3(N__16723),
            .lcout(\c0.tx.n4588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4218_3_lut_LC_7_28_5 .C_ON=1'b0;
    defparam \c0.i4218_3_lut_LC_7_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4218_3_lut_LC_7_28_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i4218_3_lut_LC_7_28_5  (
            .in0(N__22431),
            .in1(N__22232),
            .in2(_gnd_net_),
            .in3(N__20552),
            .lcout(\c0.n4573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4789_bdd_4_lut_LC_7_28_6 .C_ON=1'b0;
    defparam \c0.n4789_bdd_4_lut_LC_7_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.n4789_bdd_4_lut_LC_7_28_6 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n4789_bdd_4_lut_LC_7_28_6  (
            .in0(N__18419),
            .in1(N__16733),
            .in2(N__19604),
            .in3(N__17387),
            .lcout(),
            .ltout(tx_data_4_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_7_28_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_7_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_7_28_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_7_28_7  (
            .in0(N__22115),
            .in1(_gnd_net_),
            .in2(N__16727),
            .in3(N__16724),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22927),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4221_3_lut_LC_7_29_0 .C_ON=1'b0;
    defparam \c0.i4221_3_lut_LC_7_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4221_3_lut_LC_7_29_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4221_3_lut_LC_7_29_0  (
            .in0(N__19112),
            .in1(N__18515),
            .in2(_gnd_net_),
            .in3(N__20516),
            .lcout(\c0.n4576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_7_29_2 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_7_29_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_7_29_2  (
            .in0(N__19226),
            .in1(N__16706),
            .in2(N__19261),
            .in3(N__16697),
            .lcout(\c0.tx.n4837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4795_bdd_4_lut_LC_7_29_3 .C_ON=1'b0;
    defparam \c0.n4795_bdd_4_lut_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.n4795_bdd_4_lut_LC_7_29_3 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n4795_bdd_4_lut_LC_7_29_3  (
            .in0(N__20084),
            .in1(N__18998),
            .in2(N__19721),
            .in3(N__19601),
            .lcout(),
            .ltout(tx_data_5_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_7_29_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_7_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_7_29_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_7_29_4  (
            .in0(N__22143),
            .in1(_gnd_net_),
            .in2(N__16691),
            .in3(N__16688),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22934),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_7_29_5 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_7_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_7_29_5 .LUT_INIT=16'b0111001110000000;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_7_29_5  (
            .in0(N__19209),
            .in1(N__21853),
            .in2(N__16676),
            .in3(N__19228),
            .lcout(\c0.tx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22934),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4360_2_lut_LC_7_29_6 .C_ON=1'b0;
    defparam \c0.tx.i4360_2_lut_LC_7_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4360_2_lut_LC_7_29_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx.i4360_2_lut_LC_7_29_6  (
            .in0(N__19227),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19208),
            .lcout(),
            .ltout(\c0.tx.n4715_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_7_29_7 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_7_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_7_29_7 .LUT_INIT=16'b0011101110000000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_7_29_7  (
            .in0(N__16675),
            .in1(N__21854),
            .in2(N__16661),
            .in3(N__19256),
            .lcout(\c0.tx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22934),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i58_LC_7_30_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i58_LC_7_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i58_LC_7_30_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i58_LC_7_30_0  (
            .in0(N__16970),
            .in1(N__17294),
            .in2(_gnd_net_),
            .in3(N__17261),
            .lcout(data_in_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22939),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_375_LC_7_30_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_375_LC_7_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_375_LC_7_30_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_375_LC_7_30_1  (
            .in0(N__19139),
            .in1(N__18365),
            .in2(N__21740),
            .in3(N__19768),
            .lcout(n4_adj_970),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4203_3_lut_LC_7_30_2 .C_ON=1'b0;
    defparam \c0.tx.i4203_3_lut_LC_7_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4203_3_lut_LC_7_30_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx.i4203_3_lut_LC_7_30_2  (
            .in0(N__17237),
            .in1(N__17222),
            .in2(_gnd_net_),
            .in3(N__19206),
            .lcout(\c0.tx.n4558 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_7_30_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_7_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_7_30_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_LC_7_30_3  (
            .in0(_gnd_net_),
            .in1(N__19767),
            .in2(_gnd_net_),
            .in3(N__19132),
            .lcout(\c0.n1333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4204_3_lut_LC_7_30_4 .C_ON=1'b0;
    defparam \c0.tx.i4204_3_lut_LC_7_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4204_3_lut_LC_7_30_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx.i4204_3_lut_LC_7_30_4  (
            .in0(N__17207),
            .in1(N__17192),
            .in2(_gnd_net_),
            .in3(N__19207),
            .lcout(),
            .ltout(\c0.tx.n4559_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n4837_bdd_4_lut_LC_7_30_5 .C_ON=1'b0;
    defparam \c0.tx.n4837_bdd_4_lut_LC_7_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n4837_bdd_4_lut_LC_7_30_5 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.tx.n4837_bdd_4_lut_LC_7_30_5  (
            .in0(N__19257),
            .in1(N__17177),
            .in2(N__17171),
            .in3(N__17168),
            .lcout(\c0.tx.o_Tx_Serial_N_790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i26_LC_7_30_6 .C_ON=1'b0;
    defparam \c0.data_out_0__i26_LC_7_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i26_LC_7_30_6 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.data_out_0__i26_LC_7_30_6  (
            .in0(N__21560),
            .in1(N__19140),
            .in2(_gnd_net_),
            .in3(N__21259),
            .lcout(data_out_field_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22939),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_7_31_0 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_7_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_7_31_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_7_31_0  (
            .in0(N__17145),
            .in1(N__23501),
            .in2(_gnd_net_),
            .in3(N__17315),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22945),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i42_LC_7_31_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i42_LC_7_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i42_LC_7_31_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i42_LC_7_31_1  (
            .in0(N__16907),
            .in1(N__17451),
            .in2(_gnd_net_),
            .in3(N__16763),
            .lcout(data_in_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22945),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i2_LC_7_31_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i2_LC_7_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_7_31_2 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_7_31_2  (
            .in0(N__17418),
            .in1(N__17932),
            .in2(N__17438),
            .in3(N__17891),
            .lcout(r_Clock_Count_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22945),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4173_3_lut_LC_7_31_3 .C_ON=1'b0;
    defparam \c0.i4173_3_lut_LC_7_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4173_3_lut_LC_7_31_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4173_3_lut_LC_7_31_3  (
            .in0(N__20150),
            .in1(N__18452),
            .in2(_gnd_net_),
            .in3(N__20555),
            .lcout(\c0.n4528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4346_2_lut_LC_7_31_4 .C_ON=1'b0;
    defparam \c0.rx.i4346_2_lut_LC_7_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4346_2_lut_LC_7_31_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i4346_2_lut_LC_7_31_4  (
            .in0(N__17780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17373),
            .lcout(\c0.rx.n4667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i13_LC_7_31_5 .C_ON=1'b0;
    defparam \c0.data_out_0__i13_LC_7_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i13_LC_7_31_5 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \c0.data_out_0__i13_LC_7_31_5  (
            .in0(N__20151),
            .in1(N__21561),
            .in2(_gnd_net_),
            .in3(N__21260),
            .lcout(data_out_field_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22945),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4404_2_lut_3_lut_LC_7_31_6 .C_ON=1'b0;
    defparam \c0.rx.i4404_2_lut_3_lut_LC_7_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4404_2_lut_3_lut_LC_7_31_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.rx.i4404_2_lut_3_lut_LC_7_31_6  (
            .in0(N__17781),
            .in1(N__17633),
            .in2(_gnd_net_),
            .in3(N__17542),
            .lcout(\c0.rx.n1024 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i26_3_lut_LC_7_31_7 .C_ON=1'b0;
    defparam \c0.tx.i26_3_lut_LC_7_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i26_3_lut_LC_7_31_7 .LUT_INIT=16'b0100010001100110;
    LogicCell40 \c0.tx.i26_3_lut_LC_7_31_7  (
            .in0(N__23206),
            .in1(N__23018),
            .in2(_gnd_net_),
            .in3(N__17321),
            .lcout(\c0.tx.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_277_LC_7_32_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_277_LC_7_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_277_LC_7_32_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.i1_2_lut_adj_277_LC_7_32_0  (
            .in0(N__17762),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17517),
            .lcout(\c0.rx.n4378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_adj_271_LC_7_32_1 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_adj_271_LC_7_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_adj_271_LC_7_32_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.rx.i2_2_lut_adj_271_LC_7_32_1  (
            .in0(_gnd_net_),
            .in1(N__17684),
            .in2(_gnd_net_),
            .in3(N__17807),
            .lcout(\c0.rx.n6 ),
            .ltout(\c0.rx.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_272_LC_7_32_2 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_272_LC_7_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_272_LC_7_32_2 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \c0.rx.i1_4_lut_adj_272_LC_7_32_2  (
            .in0(N__17760),
            .in1(N__17516),
            .in2(N__17309),
            .in3(N__17627),
            .lcout(\c0.rx.n357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_adj_278_LC_7_32_3 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_adj_278_LC_7_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_adj_278_LC_7_32_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_adj_278_LC_7_32_3  (
            .in0(N__17628),
            .in1(N__17761),
            .in2(N__17544),
            .in3(N__17954),
            .lcout(),
            .ltout(\c0.rx.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_273_LC_7_32_4 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_273_LC_7_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_273_LC_7_32_4 .LUT_INIT=16'b1111001011110011;
    LogicCell40 \c0.rx.i1_4_lut_adj_273_LC_7_32_4  (
            .in0(N__17948),
            .in1(N__17629),
            .in2(N__17942),
            .in3(N__17939),
            .lcout(n1554),
            .ltout(n1554_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i6_LC_7_32_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i6_LC_7_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_7_32_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_7_32_5  (
            .in0(N__17900),
            .in1(N__17890),
            .in2(N__17861),
            .in3(N__17846),
            .lcout(r_Clock_Count_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22951),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4356_3_lut_LC_7_32_6 .C_ON=1'b0;
    defparam \c0.rx.i4356_3_lut_LC_7_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4356_3_lut_LC_7_32_6 .LUT_INIT=16'b1111111110101111;
    LogicCell40 \c0.rx.i4356_3_lut_LC_7_32_6  (
            .in0(N__17808),
            .in1(_gnd_net_),
            .in2(N__17779),
            .in3(N__17687),
            .lcout(),
            .ltout(\c0.rx.n4666_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_7_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_7_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_7_32_7 .LUT_INIT=16'b0000000101000101;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_7_32_7  (
            .in0(N__17630),
            .in1(N__17543),
            .in2(N__17567),
            .in3(N__17564),
            .lcout(\c0.rx.r_SM_Main_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22951),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_328__i0_LC_9_25_0 .C_ON=1'b1;
    defparam \c0.delay_counter_328__i0_LC_9_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_328__i0_LC_9_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_328__i0_LC_9_25_0  (
            .in0(_gnd_net_),
            .in1(N__18122),
            .in2(N__18764),
            .in3(_gnd_net_),
            .lcout(\c0.delay_counter_0 ),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(\c0.n3899 ),
            .clk(N__22921),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_328__i1_LC_9_25_1 .C_ON=1'b1;
    defparam \c0.delay_counter_328__i1_LC_9_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_328__i1_LC_9_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_328__i1_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__18710),
            .in2(_gnd_net_),
            .in3(N__17474),
            .lcout(\c0.delay_counter_1 ),
            .ltout(),
            .carryin(\c0.n3899 ),
            .carryout(\c0.n3900 ),
            .clk(N__22921),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_328__i2_LC_9_25_2 .C_ON=1'b1;
    defparam \c0.delay_counter_328__i2_LC_9_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_328__i2_LC_9_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_328__i2_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__18748),
            .in2(_gnd_net_),
            .in3(N__17471),
            .lcout(\c0.delay_counter_2 ),
            .ltout(),
            .carryin(\c0.n3900 ),
            .carryout(\c0.n3901 ),
            .clk(N__22921),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_328__i3_LC_9_25_3 .C_ON=1'b1;
    defparam \c0.delay_counter_328__i3_LC_9_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_328__i3_LC_9_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_328__i3_LC_9_25_3  (
            .in0(_gnd_net_),
            .in1(N__18683),
            .in2(_gnd_net_),
            .in3(N__18014),
            .lcout(\c0.delay_counter_3 ),
            .ltout(),
            .carryin(\c0.n3901 ),
            .carryout(\c0.n3902 ),
            .clk(N__22921),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_328__i4_LC_9_25_4 .C_ON=1'b1;
    defparam \c0.delay_counter_328__i4_LC_9_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_328__i4_LC_9_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_328__i4_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(N__18734),
            .in2(_gnd_net_),
            .in3(N__18011),
            .lcout(\c0.delay_counter_4 ),
            .ltout(),
            .carryin(\c0.n3902 ),
            .carryout(\c0.n3903 ),
            .clk(N__22921),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_328__i5_LC_9_25_5 .C_ON=1'b1;
    defparam \c0.delay_counter_328__i5_LC_9_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_328__i5_LC_9_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_328__i5_LC_9_25_5  (
            .in0(_gnd_net_),
            .in1(N__18722),
            .in2(_gnd_net_),
            .in3(N__18008),
            .lcout(\c0.delay_counter_5 ),
            .ltout(),
            .carryin(\c0.n3903 ),
            .carryout(\c0.n3904 ),
            .clk(N__22921),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_328__i6_LC_9_25_6 .C_ON=1'b1;
    defparam \c0.delay_counter_328__i6_LC_9_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_328__i6_LC_9_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_328__i6_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__18776),
            .in2(_gnd_net_),
            .in3(N__18005),
            .lcout(\c0.delay_counter_6 ),
            .ltout(),
            .carryin(\c0.n3904 ),
            .carryout(\c0.n3905 ),
            .clk(N__22921),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_328__i7_LC_9_25_7 .C_ON=1'b0;
    defparam \c0.delay_counter_328__i7_LC_9_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_328__i7_LC_9_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_328__i7_LC_9_25_7  (
            .in0(_gnd_net_),
            .in1(N__18697),
            .in2(_gnd_net_),
            .in3(N__18002),
            .lcout(\c0.delay_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22921),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i50_LC_9_26_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i50_LC_9_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i50_LC_9_26_0 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_out_0__i50_LC_9_26_0  (
            .in0(N__21577),
            .in1(N__17995),
            .in2(N__20723),
            .in3(N__21136),
            .lcout(data_out_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22928),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i40_LC_9_26_1 .C_ON=1'b0;
    defparam \c0.data_out_0__i40_LC_9_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i40_LC_9_26_1 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_out_0__i40_LC_9_26_1  (
            .in0(N__21133),
            .in1(N__17981),
            .in2(N__21735),
            .in3(N__21583),
            .lcout(\c0.data_out_field_47_N_682_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22928),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4885_bdd_4_lut_LC_9_26_2 .C_ON=1'b0;
    defparam \c0.n4885_bdd_4_lut_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.n4885_bdd_4_lut_LC_9_26_2 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n4885_bdd_4_lut_LC_9_26_2  (
            .in0(N__22324),
            .in1(N__21724),
            .in2(N__18830),
            .in3(N__20707),
            .lcout(\c0.n4888 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_612_LC_9_26_3 .C_ON=1'b0;
    defparam \c0.tx_transmit_612_LC_9_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_612_LC_9_26_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.tx_transmit_612_LC_9_26_3  (
            .in0(N__22270),
            .in1(N__22458),
            .in2(_gnd_net_),
            .in3(N__21213),
            .lcout(\c0.tx_transmit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22928),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_340_LC_9_26_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_340_LC_9_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_340_LC_9_26_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.i2_3_lut_adj_340_LC_9_26_4  (
            .in0(N__22457),
            .in1(N__21131),
            .in2(_gnd_net_),
            .in3(N__22269),
            .lcout(\c0.n2429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i47_LC_9_26_5 .C_ON=1'b0;
    defparam \c0.data_out_0__i47_LC_9_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i47_LC_9_26_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_0__i47_LC_9_26_5  (
            .in0(N__21134),
            .in1(N__21579),
            .in2(N__18116),
            .in3(N__19877),
            .lcout(\c0.data_out_field_47_N_682_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22928),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i48_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.data_out_0__i48_LC_9_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i48_LC_9_26_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.data_out_0__i48_LC_9_26_6  (
            .in0(N__22325),
            .in1(N__18095),
            .in2(N__21584),
            .in3(N__21135),
            .lcout(\c0.data_out_field_47_N_682_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22928),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i39_LC_9_26_7 .C_ON=1'b0;
    defparam \c0.data_out_0__i39_LC_9_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i39_LC_9_26_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_0__i39_LC_9_26_7  (
            .in0(N__21132),
            .in1(N__21578),
            .in2(N__18077),
            .in3(N__21814),
            .lcout(data_out_field_38),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22928),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i27_LC_9_27_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i27_LC_9_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i27_LC_9_27_0 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.data_out_0__i27_LC_9_27_0  (
            .in0(N__21542),
            .in1(N__22042),
            .in2(_gnd_net_),
            .in3(N__21145),
            .lcout(data_out_field_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22935),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i60_LC_9_27_1 .C_ON=1'b0;
    defparam \c0.data_out_0__i60_LC_9_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i60_LC_9_27_1 .LUT_INIT=16'b1100110001001110;
    LogicCell40 \c0.data_out_0__i60_LC_9_27_1  (
            .in0(N__21148),
            .in1(N__18055),
            .in2(N__22301),
            .in3(N__21545),
            .lcout(data_out_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22935),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i12_LC_9_27_2 .C_ON=1'b0;
    defparam \c0.data_out_0__i12_LC_9_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i12_LC_9_27_2 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.data_out_0__i12_LC_9_27_2  (
            .in0(N__21541),
            .in1(N__18356),
            .in2(_gnd_net_),
            .in3(N__21144),
            .lcout(data_out_field_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22935),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i33_LC_9_27_3 .C_ON=1'b0;
    defparam \c0.data_out_0__i33_LC_9_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i33_LC_9_27_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0__i33_LC_9_27_3  (
            .in0(N__21147),
            .in1(N__18508),
            .in2(N__18038),
            .in3(N__21544),
            .lcout(\c0.data_out_field_47_N_682_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22935),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_adj_359_LC_9_27_4 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_359_LC_9_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_359_LC_9_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_adj_359_LC_9_27_4  (
            .in0(N__20583),
            .in1(N__20882),
            .in2(_gnd_net_),
            .in3(N__22547),
            .lcout(),
            .ltout(n8_adj_932_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i59_LC_9_27_5 .C_ON=1'b0;
    defparam \c0.data_out_0__i59_LC_9_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i59_LC_9_27_5 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \c0.data_out_0__i59_LC_9_27_5  (
            .in0(N__18602),
            .in1(N__18229),
            .in2(N__18017),
            .in3(N__20070),
            .lcout(data_out_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22935),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i5_LC_9_27_6 .C_ON=1'b0;
    defparam \c0.data_out_0__i5_LC_9_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i5_LC_9_27_6 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.data_out_0__i5_LC_9_27_6  (
            .in0(N__21543),
            .in1(N__18450),
            .in2(_gnd_net_),
            .in3(N__21146),
            .lcout(data_out_field_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22935),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_9_27_7 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_9_27_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_LC_9_27_7  (
            .in0(N__21692),
            .in1(N__18328),
            .in2(_gnd_net_),
            .in3(N__20816),
            .lcout(n8_adj_936),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i32_LC_9_28_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i32_LC_9_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i32_LC_9_28_0 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \c0.data_out_0__i32_LC_9_28_0  (
            .in0(N__21537),
            .in1(_gnd_net_),
            .in2(N__20590),
            .in3(N__21178),
            .lcout(data_out_field_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22940),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i58_LC_9_28_1 .C_ON=1'b0;
    defparam \c0.data_out_0__i58_LC_9_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i58_LC_9_28_1 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \c0.data_out_0__i58_LC_9_28_1  (
            .in0(N__20056),
            .in1(N__18215),
            .in2(N__19322),
            .in3(N__19004),
            .lcout(data_out_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22940),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i18_LC_9_28_2 .C_ON=1'b0;
    defparam \c0.data_out_0__i18_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i18_LC_9_28_2 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.data_out_0__i18_LC_9_28_2  (
            .in0(N__21536),
            .in1(N__18265),
            .in2(_gnd_net_),
            .in3(N__21176),
            .lcout(data_out_field_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22940),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4219_3_lut_LC_9_28_3 .C_ON=1'b0;
    defparam \c0.i4219_3_lut_LC_9_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4219_3_lut_LC_9_28_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4219_3_lut_LC_9_28_3  (
            .in0(N__18327),
            .in1(N__18964),
            .in2(_gnd_net_),
            .in3(N__20495),
            .lcout(\c0.n4574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i35_LC_9_28_4 .C_ON=1'b0;
    defparam \c0.data_out_0__i35_LC_9_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i35_LC_9_28_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \c0.data_out_0__i35_LC_9_28_4  (
            .in0(N__21538),
            .in1(N__18191),
            .in2(N__18557),
            .in3(N__21179),
            .lcout(\c0.data_out_field_47_N_682_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22940),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i20_LC_9_28_5 .C_ON=1'b0;
    defparam \c0.data_out_0__i20_LC_9_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i20_LC_9_28_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \c0.data_out_0__i20_LC_9_28_5  (
            .in0(N__21177),
            .in1(N__18165),
            .in2(_gnd_net_),
            .in3(N__21539),
            .lcout(data_out_field_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22940),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i51_LC_9_28_6 .C_ON=1'b0;
    defparam \c0.data_out_0__i51_LC_9_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i51_LC_9_28_6 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \c0.data_out_0__i51_LC_9_28_6  (
            .in0(N__18143),
            .in1(N__18136),
            .in2(N__20075),
            .in3(N__18407),
            .lcout(data_out_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22940),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4210_3_lut_LC_9_28_7 .C_ON=1'b0;
    defparam \c0.i4210_3_lut_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4210_3_lut_LC_9_28_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4210_3_lut_LC_9_28_7  (
            .in0(N__22031),
            .in1(N__20235),
            .in2(_gnd_net_),
            .in3(N__20496),
            .lcout(\c0.n4565 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_385_LC_9_29_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_385_LC_9_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_385_LC_9_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_385_LC_9_29_1  (
            .in0(N__20578),
            .in1(N__18261),
            .in2(_gnd_net_),
            .in3(N__18509),
            .lcout(\c0.n1312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_4_lut_adj_384_LC_9_29_2 .C_ON=1'b0;
    defparam \c0.i4_3_lut_4_lut_adj_384_LC_9_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_4_lut_adj_384_LC_9_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_3_lut_4_lut_adj_384_LC_9_29_2  (
            .in0(N__18510),
            .in1(N__20579),
            .in2(N__20237),
            .in3(N__18475),
            .lcout(),
            .ltout(n11_adj_967_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i61_LC_9_29_3 .C_ON=1'b0;
    defparam \c0.data_out_0__i61_LC_9_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i61_LC_9_29_3 .LUT_INIT=16'b1110110100100001;
    LogicCell40 \c0.data_out_0__i61_LC_9_29_3  (
            .in0(N__18857),
            .in1(N__20062),
            .in2(N__18386),
            .in3(N__18379),
            .lcout(data_out_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22946),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_9_29_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_9_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_9_29_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_9_29_4  (
            .in0(N__21815),
            .in1(N__18357),
            .in2(_gnd_net_),
            .in3(N__21728),
            .lcout(),
            .ltout(\c0.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_9_29_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_9_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_9_29_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_LC_9_29_5  (
            .in0(N__21672),
            .in1(N__22038),
            .in2(N__18332),
            .in3(N__18329),
            .lcout(\c0.n4456 ),
            .ltout(\c0.n4456_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_386_LC_9_29_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_386_LC_9_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_386_LC_9_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_386_LC_9_29_6  (
            .in0(_gnd_net_),
            .in1(N__18592),
            .in2(N__18290),
            .in3(N__19105),
            .lcout(n1255),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i41_LC_9_29_7 .C_ON=1'b0;
    defparam \c0.data_out_0__i41_LC_9_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i41_LC_9_29_7 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0__i41_LC_9_29_7  (
            .in0(N__19106),
            .in1(N__21576),
            .in2(N__18287),
            .in3(N__21246),
            .lcout(\c0.data_out_field_47_N_682_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22946),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4207_3_lut_LC_9_30_0 .C_ON=1'b0;
    defparam \c0.i4207_3_lut_LC_9_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4207_3_lut_LC_9_30_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.i4207_3_lut_LC_9_30_0  (
            .in0(N__20494),
            .in1(N__18266),
            .in2(_gnd_net_),
            .in3(N__19142),
            .lcout(\c0.n4562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_9_30_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_9_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_9_30_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_9_30_1  (
            .in0(N__18596),
            .in1(N__19110),
            .in2(N__20345),
            .in3(N__20162),
            .lcout(n4462),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i4_LC_9_30_2 .C_ON=1'b0;
    defparam \c0.data_out_0__i4_LC_9_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i4_LC_9_30_2 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \c0.data_out_0__i4_LC_9_30_2  (
            .in0(N__21242),
            .in1(N__18471),
            .in2(_gnd_net_),
            .in3(N__21524),
            .lcout(data_out_field_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22952),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_364_LC_9_30_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_364_LC_9_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_364_LC_9_30_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_364_LC_9_30_3  (
            .in0(_gnd_net_),
            .in1(N__18556),
            .in2(_gnd_net_),
            .in3(N__18901),
            .lcout(),
            .ltout(\c0.n1384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_350_LC_9_30_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_350_LC_9_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_350_LC_9_30_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_350_LC_9_30_4  (
            .in0(N__19886),
            .in1(N__18446),
            .in2(N__18518),
            .in3(N__18511),
            .lcout(n10_adj_947),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_365_LC_9_30_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_365_LC_9_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_365_LC_9_30_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_365_LC_9_30_5  (
            .in0(N__18470),
            .in1(N__18926),
            .in2(N__18451),
            .in3(N__22348),
            .lcout(\c0.n4465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4174_3_lut_LC_9_30_7 .C_ON=1'b0;
    defparam \c0.i4174_3_lut_LC_9_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4174_3_lut_LC_9_30_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4174_3_lut_LC_9_30_7  (
            .in0(N__20891),
            .in1(N__20194),
            .in2(_gnd_net_),
            .in3(N__20493),
            .lcout(\c0.n4529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i14_LC_10_23_7 .C_ON=1'b0;
    defparam \c0.data_out_0__i14_LC_10_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i14_LC_10_23_7 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \c0.data_out_0__i14_LC_10_23_7  (
            .in0(N__20913),
            .in1(N__21522),
            .in2(_gnd_net_),
            .in3(N__21258),
            .lcout(data_out_field_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i10_LC_10_24_6 .C_ON=1'b0;
    defparam \c0.data_out_0__i10_LC_10_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i10_LC_10_24_6 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.data_out_0__i10_LC_10_24_6  (
            .in0(N__21433),
            .in1(N__21768),
            .in2(_gnd_net_),
            .in3(N__21234),
            .lcout(data_out_field_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_10_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__19632),
            .in2(_gnd_net_),
            .in3(N__22231),
            .lcout(n7_adj_937),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i16_LC_10_25_2 .C_ON=1'b0;
    defparam \c0.data_out_0__i16_LC_10_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i16_LC_10_25_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \c0.data_out_0__i16_LC_10_25_2  (
            .in0(N__21917),
            .in1(N__21444),
            .in2(_gnd_net_),
            .in3(N__21214),
            .lcout(data_out_field_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22922),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_374_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_374_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_374_LC_10_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_374_LC_10_25_3  (
            .in0(N__18775),
            .in1(N__18760),
            .in2(N__18749),
            .in3(N__18733),
            .lcout(\c0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_373_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_373_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_373_LC_10_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_373_LC_10_25_4  (
            .in0(N__18721),
            .in1(N__18709),
            .in2(N__18698),
            .in3(N__18682),
            .lcout(),
            .ltout(\c0.n14_adj_902_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_10_25_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_10_25_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_10_25_5  (
            .in0(N__22459),
            .in1(N__18671),
            .in2(N__18665),
            .in3(N__22271),
            .lcout(n3580),
            .ltout(n3580_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i45_LC_10_25_6 .C_ON=1'b0;
    defparam \c0.data_out_0__i45_LC_10_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i45_LC_10_25_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.data_out_0__i45_LC_10_25_6  (
            .in0(N__20849),
            .in1(N__18662),
            .in2(N__18647),
            .in3(N__21215),
            .lcout(\c0.data_out_field_47_N_682_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22922),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i36_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i36_LC_10_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i36_LC_10_26_0 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_out_0__i36_LC_10_26_0  (
            .in0(N__21436),
            .in1(N__19821),
            .in2(N__18644),
            .in3(N__21152),
            .lcout(\c0.data_out_field_47_N_682_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22929),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i44_LC_10_26_1 .C_ON=1'b0;
    defparam \c0.data_out_0__i44_LC_10_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i44_LC_10_26_1 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0__i44_LC_10_26_1  (
            .in0(N__21153),
            .in1(N__21956),
            .in2(N__18623),
            .in3(N__21438),
            .lcout(data_out_field_43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22929),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_10_26_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_10_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_10_26_2  (
            .in0(N__21891),
            .in1(N__18966),
            .in2(_gnd_net_),
            .in3(N__19876),
            .lcout(n7_adj_933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_363_LC_10_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_363_LC_10_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_363_LC_10_26_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_363_LC_10_26_3  (
            .in0(_gnd_net_),
            .in1(N__21992),
            .in2(_gnd_net_),
            .in3(N__21890),
            .lcout(\c0.n4393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i23_LC_10_26_4 .C_ON=1'b0;
    defparam \c0.data_out_0__i23_LC_10_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i23_LC_10_26_4 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.data_out_0__i23_LC_10_26_4  (
            .in0(N__21434),
            .in1(N__19633),
            .in2(_gnd_net_),
            .in3(N__21149),
            .lcout(data_out_field_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22929),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_10_26_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_10_26_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_LC_10_26_5  (
            .in0(N__18845),
            .in1(N__20644),
            .in2(N__19037),
            .in3(N__20438),
            .lcout(\c0.n4885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i29_LC_10_26_6 .C_ON=1'b0;
    defparam \c0.data_out_0__i29_LC_10_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i29_LC_10_26_6 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.data_out_0__i29_LC_10_26_6  (
            .in0(N__21435),
            .in1(N__20883),
            .in2(_gnd_net_),
            .in3(N__21150),
            .lcout(data_out_field_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22929),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i31_LC_10_26_7 .C_ON=1'b0;
    defparam \c0.data_out_0__i31_LC_10_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i31_LC_10_26_7 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \c0.data_out_0__i31_LC_10_26_7  (
            .in0(N__21151),
            .in1(N__21892),
            .in2(_gnd_net_),
            .in3(N__21437),
            .lcout(data_out_field_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22929),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i46_LC_10_27_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i46_LC_10_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i46_LC_10_27_0 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \c0.data_out_0__i46_LC_10_27_0  (
            .in0(N__21143),
            .in1(N__18821),
            .in2(N__21526),
            .in3(N__19945),
            .lcout(\c0.data_out_field_47_N_682_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i17_LC_10_27_1 .C_ON=1'b0;
    defparam \c0.data_out_0__i17_LC_10_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i17_LC_10_27_1 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \c0.data_out_0__i17_LC_10_27_1  (
            .in0(N__18967),
            .in1(N__21464),
            .in2(_gnd_net_),
            .in3(N__21142),
            .lcout(data_out_field_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_376_LC_10_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_376_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_376_LC_10_27_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_376_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(N__19483),
            .in2(_gnd_net_),
            .in3(N__19837),
            .lcout(),
            .ltout(\c0.n6_adj_904_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_377_LC_10_27_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_377_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_377_LC_10_27_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_377_LC_10_27_3  (
            .in0(N__19447),
            .in1(N__19408),
            .in2(N__18803),
            .in3(N__19369),
            .lcout(n7_adj_938),
            .ltout(n7_adj_938_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i52_LC_10_27_4 .C_ON=1'b0;
    defparam \c0.data_out_0__i52_LC_10_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i52_LC_10_27_4 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_0__i52_LC_10_27_4  (
            .in0(N__21462),
            .in1(N__21644),
            .in2(N__18800),
            .in3(N__18797),
            .lcout(data_out_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i11_LC_10_27_5 .C_ON=1'b0;
    defparam \c0.data_out_0__i11_LC_10_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i11_LC_10_27_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.data_out_0__i11_LC_10_27_5  (
            .in0(N__21671),
            .in1(N__21463),
            .in2(_gnd_net_),
            .in3(N__21141),
            .lcout(data_out_field_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_370_LC_10_27_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_370_LC_10_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_370_LC_10_27_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_370_LC_10_27_6  (
            .in0(N__18925),
            .in1(N__19817),
            .in2(_gnd_net_),
            .in3(N__20809),
            .lcout(n7_adj_935),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_356_LC_10_27_7 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_356_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_356_LC_10_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_356_LC_10_27_7  (
            .in0(N__20856),
            .in1(N__18905),
            .in2(N__18866),
            .in3(N__18965),
            .lcout(n12_adj_966),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_379_LC_10_28_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_379_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_379_LC_10_28_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_379_LC_10_28_0  (
            .in0(_gnd_net_),
            .in1(N__21448),
            .in2(_gnd_net_),
            .in3(N__21137),
            .lcout(n1677),
            .ltout(n1677_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i56_LC_10_28_1 .C_ON=1'b0;
    defparam \c0.data_out_0__i56_LC_10_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i56_LC_10_28_1 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \c0.data_out_0__i56_LC_10_28_1  (
            .in0(N__22490),
            .in1(N__18844),
            .in2(N__18848),
            .in3(N__18989),
            .lcout(data_out_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22941),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i22_LC_10_28_2 .C_ON=1'b0;
    defparam \c0.data_out_0__i22_LC_10_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i22_LC_10_28_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \c0.data_out_0__i22_LC_10_28_2  (
            .in0(N__20759),
            .in1(N__21449),
            .in2(_gnd_net_),
            .in3(N__21139),
            .lcout(data_out_field_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22941),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i21_LC_10_28_3 .C_ON=1'b0;
    defparam \c0.data_out_0__i21_LC_10_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i21_LC_10_28_3 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \c0.data_out_0__i21_LC_10_28_3  (
            .in0(N__21138),
            .in1(N__21466),
            .in2(_gnd_net_),
            .in3(N__20193),
            .lcout(data_out_field_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22941),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i6_LC_10_28_4 .C_ON=1'b0;
    defparam \c0.data_out_0__i6_LC_10_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i6_LC_10_28_4 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.data_out_0__i6_LC_10_28_4  (
            .in0(N__21465),
            .in1(N__20263),
            .in2(_gnd_net_),
            .in3(N__21140),
            .lcout(data_out_field_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22941),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_366_LC_10_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_366_LC_10_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_366_LC_10_28_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_366_LC_10_28_5  (
            .in0(_gnd_net_),
            .in1(N__20755),
            .in2(_gnd_net_),
            .in3(N__22329),
            .lcout(\c0.n4483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_LC_10_28_6 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_LC_10_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_LC_10_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_LC_10_28_6  (
            .in0(N__22330),
            .in1(N__19664),
            .in2(N__20764),
            .in3(N__20262),
            .lcout(),
            .ltout(n8_adj_934_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i64_LC_10_28_7 .C_ON=1'b0;
    defparam \c0.data_out_0__i64_LC_10_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i64_LC_10_28_7 .LUT_INIT=16'b1100110010100101;
    LogicCell40 \c0.data_out_0__i64_LC_10_28_7  (
            .in0(N__19046),
            .in1(N__19033),
            .in2(N__19040),
            .in3(N__20063),
            .lcout(data_out_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22941),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_361_LC_10_29_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_361_LC_10_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_361_LC_10_29_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_361_LC_10_29_0  (
            .in0(N__19019),
            .in1(N__20299),
            .in2(N__20990),
            .in3(N__20092),
            .lcout(\c0.n4447 ),
            .ltout(\c0.n4447_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_10_29_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_10_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_10_29_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i3_2_lut_LC_10_29_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19007),
            .in3(N__19982),
            .lcout(n9_adj_972),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4473_LC_10_29_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4473_LC_10_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_4473_LC_10_29_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_4473_LC_10_29_2  (
            .in0(N__20689),
            .in1(N__19148),
            .in2(N__19568),
            .in3(N__19922),
            .lcout(\c0.n4795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_4_lut_LC_10_29_3 .C_ON=1'b0;
    defparam \c0.i4_3_lut_4_lut_LC_10_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_4_lut_LC_10_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_3_lut_4_lut_LC_10_29_3  (
            .in0(N__20093),
            .in1(N__20858),
            .in2(N__19955),
            .in3(N__19983),
            .lcout(n11_adj_945),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i54_LC_10_29_4 .C_ON=1'b0;
    defparam \c0.data_out_0__i54_LC_10_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i54_LC_10_29_4 .LUT_INIT=16'b1111011000000110;
    LogicCell40 \c0.data_out_0__i54_LC_10_29_4  (
            .in0(N__22063),
            .in1(N__18980),
            .in2(N__20074),
            .in3(N__19160),
            .lcout(data_out_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22947),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_368_LC_10_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_368_LC_10_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_368_LC_10_29_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_368_LC_10_29_5  (
            .in0(_gnd_net_),
            .in1(N__19878),
            .in2(_gnd_net_),
            .in3(N__18968),
            .lcout(\c0.n4417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_383_LC_10_29_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_383_LC_10_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_383_LC_10_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_383_LC_10_29_6  (
            .in0(N__19984),
            .in1(N__19953),
            .in2(_gnd_net_),
            .in3(N__18935),
            .lcout(),
            .ltout(n7_adj_969_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i57_LC_10_29_7 .C_ON=1'b0;
    defparam \c0.data_out_0__i57_LC_10_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i57_LC_10_29_7 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \c0.data_out_0__i57_LC_10_29_7  (
            .in0(N__20055),
            .in1(N__19706),
            .in2(N__18929),
            .in3(N__19697),
            .lcout(data_out_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22947),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i19_LC_10_30_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i19_LC_10_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i19_LC_10_30_0 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.data_out_0__i19_LC_10_30_0  (
            .in0(N__21523),
            .in1(N__20234),
            .in2(_gnd_net_),
            .in3(N__21238),
            .lcout(data_out_field_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22953),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_LC_10_30_2 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_LC_10_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_LC_10_30_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i2_3_lut_LC_10_30_2  (
            .in0(N__19265),
            .in1(N__19235),
            .in2(_gnd_net_),
            .in3(N__19211),
            .lcout(\c0.tx.n84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4261_3_lut_LC_10_30_3 .C_ON=1'b0;
    defparam \c0.i4261_3_lut_LC_10_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4261_3_lut_LC_10_30_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4261_3_lut_LC_10_30_3  (
            .in0(N__19966),
            .in1(N__19159),
            .in2(_gnd_net_),
            .in3(N__20479),
            .lcout(\c0.n4616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_287_LC_10_30_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_287_LC_10_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_287_LC_10_30_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_287_LC_10_30_6  (
            .in0(N__19141),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19111),
            .lcout(n4480),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4206_3_lut_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.i4206_3_lut_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4206_3_lut_LC_11_24_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i4206_3_lut_LC_11_24_1  (
            .in0(N__20989),
            .in1(N__21767),
            .in2(_gnd_net_),
            .in3(N__20478),
            .lcout(\c0.n4561 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i43_LC_11_25_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i43_LC_11_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i43_LC_11_25_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0__i43_LC_11_25_0  (
            .in0(N__21248),
            .in1(N__20328),
            .in2(N__19067),
            .in3(N__21447),
            .lcout(\c0.data_out_field_47_N_682_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22930),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i3_LC_11_25_3 .C_ON=1'b0;
    defparam \c0.data_out_0__i3_LC_11_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i3_LC_11_25_3 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.data_out_0__i3_LC_11_25_3  (
            .in0(N__21996),
            .in1(N__21445),
            .in2(_gnd_net_),
            .in3(N__21247),
            .lcout(data_out_field_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22930),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4502_LC_11_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4502_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4502_LC_11_25_4 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_4502_LC_11_25_4  (
            .in0(N__20477),
            .in1(N__21872),
            .in2(N__19634),
            .in3(N__20681),
            .lcout(),
            .ltout(\c0.n4771_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4771_bdd_4_lut_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.n4771_bdd_4_lut_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.n4771_bdd_4_lut_LC_11_25_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n4771_bdd_4_lut_LC_11_25_5  (
            .in0(N__20682),
            .in1(N__20360),
            .in2(N__19049),
            .in3(N__19657),
            .lcout(),
            .ltout(\c0.n4774_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i276843_i1_3_lut_LC_11_25_6 .C_ON=1'b0;
    defparam \c0.i276843_i1_3_lut_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i276843_i1_3_lut_LC_11_25_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.i276843_i1_3_lut_LC_11_25_6  (
            .in0(_gnd_net_),
            .in1(N__20930),
            .in2(N__19337),
            .in3(N__19561),
            .lcout(tx_data_6_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_360_LC_11_25_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_360_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_360_LC_11_25_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_360_LC_11_25_7  (
            .in0(N__22081),
            .in1(N__22391),
            .in2(N__22000),
            .in3(N__20845),
            .lcout(n10_adj_971),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i8_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i8_LC_11_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i8_LC_11_26_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \c0.data_out_0__i8_LC_11_26_0  (
            .in0(N__19281),
            .in1(N__21446),
            .in2(_gnd_net_),
            .in3(N__21184),
            .lcout(data_out_field_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i7_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.data_out_0__i7_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i7_LC_11_26_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.data_out_0__i7_LC_11_26_1  (
            .in0(N__21183),
            .in1(N__21442),
            .in2(_gnd_net_),
            .in3(N__19656),
            .lcout(data_out_field_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i37_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.data_out_0__i37_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i37_LC_11_26_2 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_out_0__i37_LC_11_26_2  (
            .in0(N__21440),
            .in1(N__20807),
            .in2(N__19307),
            .in3(N__21185),
            .lcout(\c0.data_out_field_47_N_682_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i3_LC_11_26_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i3_LC_11_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i3_LC_11_26_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i3_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(N__21441),
            .in2(_gnd_net_),
            .in3(N__19484),
            .lcout(\c0.byte_transmit_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i2_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.data_out_0__i2_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i2_LC_11_26_4 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.data_out_0__i2_LC_11_26_4  (
            .in0(N__21439),
            .in1(N__20984),
            .in2(_gnd_net_),
            .in3(N__21182),
            .lcout(data_out_field_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i55_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.data_out_0__i55_LC_11_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i55_LC_11_26_5 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0__i55_LC_11_26_5  (
            .in0(N__21186),
            .in1(N__19916),
            .in2(N__22010),
            .in3(N__21443),
            .lcout(data_out_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_380_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_380_LC_11_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_380_LC_11_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_380_LC_11_26_6  (
            .in0(N__21602),
            .in1(N__19813),
            .in2(N__19285),
            .in3(N__20806),
            .lcout(n1246),
            .ltout(n1246_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_11_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_11_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_LC_11_26_7  (
            .in0(_gnd_net_),
            .in1(N__19655),
            .in2(N__19637),
            .in3(N__19628),
            .lcout(n4438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i0_LC_11_27_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter__i0_LC_11_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i0_LC_11_27_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \c0.byte_transmit_counter__i0_LC_11_27_0  (
            .in0(_gnd_net_),
            .in1(N__22283),
            .in2(N__20453),
            .in3(N__20054),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(bfn_11_27_0_),
            .carryout(\c0.n3844 ),
            .clk(N__22942),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i1_LC_11_27_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter__i1_LC_11_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i1_LC_11_27_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.byte_transmit_counter__i1_LC_11_27_1  (
            .in0(N__20053),
            .in1(N__20643),
            .in2(_gnd_net_),
            .in3(N__19607),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(\c0.n3844 ),
            .carryout(\c0.n3845 ),
            .clk(N__22942),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i2_LC_11_27_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter__i2_LC_11_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i2_LC_11_27_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.byte_transmit_counter__i2_LC_11_27_2  (
            .in0(N__20061),
            .in1(N__19522),
            .in2(_gnd_net_),
            .in3(N__19493),
            .lcout(\c0.byte_transmit_counter_2 ),
            .ltout(),
            .carryin(\c0.n3845 ),
            .carryout(\c0.n3846 ),
            .clk(N__22942),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_637_5_lut_LC_11_27_3 .C_ON=1'b1;
    defparam \c0.add_637_5_lut_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_637_5_lut_LC_11_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_637_5_lut_LC_11_27_3  (
            .in0(_gnd_net_),
            .in1(N__19490),
            .in2(_gnd_net_),
            .in3(N__19472),
            .lcout(\c0.tx_transmit_N_274_3 ),
            .ltout(),
            .carryin(\c0.n3846 ),
            .carryout(\c0.n3847 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_637_6_lut_LC_11_27_4 .C_ON=1'b1;
    defparam \c0.add_637_6_lut_LC_11_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_637_6_lut_LC_11_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_637_6_lut_LC_11_27_4  (
            .in0(_gnd_net_),
            .in1(N__19469),
            .in2(_gnd_net_),
            .in3(N__19436),
            .lcout(\c0.tx_transmit_N_274_4 ),
            .ltout(),
            .carryin(\c0.n3847 ),
            .carryout(\c0.n3848 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_637_7_lut_LC_11_27_5 .C_ON=1'b1;
    defparam \c0.add_637_7_lut_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_637_7_lut_LC_11_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_637_7_lut_LC_11_27_5  (
            .in0(_gnd_net_),
            .in1(N__19433),
            .in2(_gnd_net_),
            .in3(N__19397),
            .lcout(\c0.tx_transmit_N_274_5 ),
            .ltout(),
            .carryin(\c0.n3848 ),
            .carryout(\c0.n3849 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_637_8_lut_LC_11_27_6 .C_ON=1'b1;
    defparam \c0.add_637_8_lut_LC_11_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_637_8_lut_LC_11_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_637_8_lut_LC_11_27_6  (
            .in0(_gnd_net_),
            .in1(N__19394),
            .in2(_gnd_net_),
            .in3(N__19358),
            .lcout(\c0.tx_transmit_N_274_6 ),
            .ltout(),
            .carryin(\c0.n3849 ),
            .carryout(\c0.n3850 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_637_9_lut_LC_11_27_7 .C_ON=1'b0;
    defparam \c0.add_637_9_lut_LC_11_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_637_9_lut_LC_11_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_637_9_lut_LC_11_27_7  (
            .in0(_gnd_net_),
            .in1(N__19355),
            .in2(_gnd_net_),
            .in3(N__19340),
            .lcout(\c0.tx_transmit_N_274_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_4_lut_LC_11_28_0 .C_ON=1'b0;
    defparam \c0.i3_2_lut_4_lut_LC_11_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_4_lut_LC_11_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_2_lut_4_lut_LC_11_28_0  (
            .in0(N__20236),
            .in1(N__20192),
            .in2(N__20264),
            .in3(N__19826),
            .lcout(),
            .ltout(n9_adj_948_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i63_LC_11_28_1 .C_ON=1'b0;
    defparam \c0.data_out_0__i63_LC_11_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i63_LC_11_28_1 .LUT_INIT=16'b1110101101000001;
    LogicCell40 \c0.data_out_0__i63_LC_11_28_1  (
            .in0(N__20057),
            .in1(N__19787),
            .in2(N__19775),
            .in3(N__19903),
            .lcout(data_out_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22948),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i24_LC_11_28_2 .C_ON=1'b0;
    defparam \c0.data_out_0__i24_LC_11_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i24_LC_11_28_2 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.data_out_0__i24_LC_11_28_2  (
            .in0(N__21485),
            .in1(N__22192),
            .in2(_gnd_net_),
            .in3(N__21180),
            .lcout(data_out_field_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22948),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i28_LC_11_28_3 .C_ON=1'b0;
    defparam \c0.data_out_0__i28_LC_11_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i28_LC_11_28_3 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \c0.data_out_0__i28_LC_11_28_3  (
            .in0(N__21181),
            .in1(N__19758),
            .in2(_gnd_net_),
            .in3(N__21486),
            .lcout(data_out_field_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22948),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i49_LC_11_28_4 .C_ON=1'b0;
    defparam \c0.data_out_0__i49_LC_11_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i49_LC_11_28_4 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \c0.data_out_0__i49_LC_11_28_4  (
            .in0(N__19685),
            .in1(N__20108),
            .in2(N__19736),
            .in3(N__20058),
            .lcout(data_out_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22948),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4176_3_lut_LC_11_28_5 .C_ON=1'b0;
    defparam \c0.i4176_3_lut_LC_11_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4176_3_lut_LC_11_28_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.i4176_3_lut_LC_11_28_5  (
            .in0(N__20923),
            .in1(N__20452),
            .in2(_gnd_net_),
            .in3(N__20258),
            .lcout(\c0.n4531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_adj_362_LC_11_28_6 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_362_LC_11_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_362_LC_11_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_adj_362_LC_11_28_6  (
            .in0(N__22373),
            .in1(N__22439),
            .in2(_gnd_net_),
            .in3(N__20924),
            .lcout(n8_adj_968),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4222_3_lut_LC_11_28_7 .C_ON=1'b0;
    defparam \c0.i4222_3_lut_LC_11_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4222_3_lut_LC_11_28_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.i4222_3_lut_LC_11_28_7  (
            .in0(N__19696),
            .in1(N__20451),
            .in2(_gnd_net_),
            .in3(N__19684),
            .lcout(\c0.n4577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i53_LC_11_29_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i53_LC_11_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i53_LC_11_29_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_out_0__i53_LC_11_29_0  (
            .in0(N__20284),
            .in1(_gnd_net_),
            .in2(N__20306),
            .in3(N__20060),
            .lcout(data_out_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22954),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_367_LC_11_29_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_367_LC_11_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_367_LC_11_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_367_LC_11_29_1  (
            .in0(N__20257),
            .in1(N__20224),
            .in2(_gnd_net_),
            .in3(N__20185),
            .lcout(),
            .ltout(\c0.n4432_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_369_LC_11_29_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_369_LC_11_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_369_LC_11_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_369_LC_11_29_2  (
            .in0(N__21775),
            .in1(N__20161),
            .in2(N__20129),
            .in3(N__20126),
            .lcout(),
            .ltout(\c0.n10_adj_900_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_371_LC_11_29_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_371_LC_11_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_371_LC_11_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_371_LC_11_29_3  (
            .in0(N__20120),
            .in1(N__22162),
            .in2(N__20111),
            .in3(N__20107),
            .lcout(\c0.n4489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4177_3_lut_LC_11_29_4 .C_ON=1'b0;
    defparam \c0.i4177_3_lut_LC_11_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4177_3_lut_LC_11_29_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i4177_3_lut_LC_11_29_4  (
            .in0(N__20954),
            .in1(N__20760),
            .in2(_gnd_net_),
            .in3(N__20466),
            .lcout(\c0.n4532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i62_LC_11_29_5 .C_ON=1'b0;
    defparam \c0.data_out_0__i62_LC_11_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i62_LC_11_29_5 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \c0.data_out_0__i62_LC_11_29_5  (
            .in0(N__20059),
            .in1(N__19967),
            .in2(N__19954),
            .in3(N__19991),
            .lcout(\c0.data_out_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22954),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4260_3_lut_LC_11_29_6 .C_ON=1'b0;
    defparam \c0.i4260_3_lut_LC_11_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4260_3_lut_LC_11_29_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i4260_3_lut_LC_11_29_6  (
            .in0(N__21608),
            .in1(N__19946),
            .in2(_gnd_net_),
            .in3(N__20465),
            .lcout(\c0.n4615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4507_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4507_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4507_LC_12_25_2 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_4507_LC_12_25_2  (
            .in0(N__19915),
            .in1(N__20679),
            .in2(N__20517),
            .in3(N__19904),
            .lcout(),
            .ltout(\c0.n4879_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n4879_bdd_4_lut_LC_12_25_3 .C_ON=1'b0;
    defparam \c0.n4879_bdd_4_lut_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.n4879_bdd_4_lut_LC_12_25_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n4879_bdd_4_lut_LC_12_25_3  (
            .in0(N__20680),
            .in1(N__21823),
            .in2(N__19889),
            .in3(N__19885),
            .lcout(\c0.n4882 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_290_LC_12_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_290_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_290_LC_12_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_290_LC_12_25_5  (
            .in0(N__21918),
            .in1(N__21990),
            .in2(_gnd_net_),
            .in3(N__21893),
            .lcout(\c0.n1378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_387_LC_12_25_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_387_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_387_LC_12_25_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_387_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(N__20922),
            .in2(_gnd_net_),
            .in3(N__20890),
            .lcout(n4423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i15_LC_12_26_0 .C_ON=1'b0;
    defparam \c0.data_out_0__i15_LC_12_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i15_LC_12_26_0 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.data_out_0__i15_LC_12_26_0  (
            .in0(N__20359),
            .in1(N__21555),
            .in2(_gnd_net_),
            .in3(N__21250),
            .lcout(data_out_field_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22943),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4263_3_lut_LC_12_26_1 .C_ON=1'b0;
    defparam \c0.i4263_3_lut_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4263_3_lut_LC_12_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i4263_3_lut_LC_12_26_1  (
            .in0(N__20423),
            .in1(N__20857),
            .in2(_gnd_net_),
            .in3(N__20808),
            .lcout(\c0.n4618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4368_4_lut_LC_12_26_2.C_ON=1'b0;
    defparam i4368_4_lut_LC_12_26_2.SEQ_MODE=4'b0000;
    defparam i4368_4_lut_LC_12_26_2.LUT_INIT=16'b0110100110010110;
    LogicCell40 i4368_4_lut_LC_12_26_2 (
            .in0(N__20768),
            .in1(N__22166),
            .in2(N__20735),
            .in3(N__21822),
            .lcout(n4663),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i30_LC_12_26_3 .C_ON=1'b0;
    defparam \c0.data_out_0__i30_LC_12_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i30_LC_12_26_3 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \c0.data_out_0__i30_LC_12_26_3  (
            .in0(N__21251),
            .in1(N__20950),
            .in2(_gnd_net_),
            .in3(N__21559),
            .lcout(data_out_field_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22943),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4417_LC_12_26_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4417_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_4417_LC_12_26_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_4417_LC_12_26_4  (
            .in0(N__22193),
            .in1(N__20660),
            .in2(N__20594),
            .in3(N__20424),
            .lcout(\c0.n4765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_372_LC_12_26_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_372_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_372_LC_12_26_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_372_LC_12_26_5  (
            .in0(_gnd_net_),
            .in1(N__20358),
            .in2(_gnd_net_),
            .in3(N__20327),
            .lcout(\c0.n1421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4372_4_lut_LC_12_26_6.C_ON=1'b0;
    defparam i4372_4_lut_LC_12_26_6.SEQ_MODE=4'b0000;
    defparam i4372_4_lut_LC_12_26_6.LUT_INIT=16'b0110100110010110;
    LogicCell40 i4372_4_lut_LC_12_26_6 (
            .in0(N__21959),
            .in1(N__22082),
            .in2(N__22067),
            .in3(N__22043),
            .lcout(n4655),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_12_26_7  (
            .in0(N__21991),
            .in1(N__21958),
            .in2(N__21935),
            .in3(N__21889),
            .lcout(\c0.n4453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_LC_12_27_0 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.tx.i1_4_lut_LC_12_27_0  (
            .in0(N__23014),
            .in1(N__23453),
            .in2(N__23201),
            .in3(N__23069),
            .lcout(\c0.tx.n1514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_12_27_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_12_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_LC_12_27_1  (
            .in0(N__21824),
            .in1(N__21606),
            .in2(N__21779),
            .in3(N__21736),
            .lcout(n4426),
            .ltout(n4426_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4370_4_lut_LC_12_27_2.C_ON=1'b0;
    defparam i4370_4_lut_LC_12_27_2.SEQ_MODE=4'b0000;
    defparam i4370_4_lut_LC_12_27_2.LUT_INIT=16'b0110100110010110;
    LogicCell40 i4370_4_lut_LC_12_27_2 (
            .in0(N__22191),
            .in1(N__22525),
            .in2(N__21683),
            .in3(N__21676),
            .lcout(n4659),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i38_LC_12_27_3 .C_ON=1'b0;
    defparam \c0.data_out_0__i38_LC_12_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i38_LC_12_27_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_0__i38_LC_12_27_3  (
            .in0(N__21220),
            .in1(N__21564),
            .in2(N__21632),
            .in3(N__21607),
            .lcout(\c0.data_out_field_47_N_682_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22949),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__i9_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.data_out_0__i9_LC_12_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__i9_LC_12_27_4 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.data_out_0__i9_LC_12_27_4  (
            .in0(N__21563),
            .in1(N__22221),
            .in2(_gnd_net_),
            .in3(N__21219),
            .lcout(data_out_field_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22949),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_378_LC_12_27_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_378_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_378_LC_12_27_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_378_LC_12_27_6  (
            .in0(N__20985),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20946),
            .lcout(\c0.n1306 ),
            .ltout(\c0.n1306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_358_LC_12_27_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_358_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_358_LC_12_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_358_LC_12_27_7  (
            .in0(N__22369),
            .in1(N__22355),
            .in2(N__22337),
            .in3(N__22334),
            .lcout(n4454),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_prev_611_LC_12_28_0 .C_ON=1'b0;
    defparam \c0.tx_active_prev_611_LC_12_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx_active_prev_611_LC_12_28_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.tx_active_prev_611_LC_12_28_0  (
            .in0(N__22254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.tx_active_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22955),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_343_LC_12_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_343_LC_12_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_343_LC_12_28_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i1_2_lut_adj_343_LC_12_28_1  (
            .in0(_gnd_net_),
            .in1(N__22289),
            .in2(_gnd_net_),
            .in3(N__22252),
            .lcout(\c0.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_12_28_2 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_12_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_12_28_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx.i1_2_lut_LC_12_28_2  (
            .in0(_gnd_net_),
            .in1(N__22992),
            .in2(_gnd_net_),
            .in3(N__23072),
            .lcout(),
            .ltout(\c0.tx.n2908_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_LC_12_28_3 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_LC_12_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_LC_12_28_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.tx.i2_4_lut_LC_12_28_3  (
            .in0(N__23161),
            .in1(N__22088),
            .in2(N__22277),
            .in3(N__23472),
            .lcout(),
            .ltout(\c0.tx.n1457_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_12_28_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_12_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_12_28_4 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_12_28_4  (
            .in0(N__22253),
            .in1(_gnd_net_),
            .in2(N__22274),
            .in3(N__23162),
            .lcout(\c0.tx_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22955),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_288_LC_12_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_288_LC_12_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_288_LC_12_28_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_288_LC_12_28_5  (
            .in0(N__22214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22187),
            .lcout(n1325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_4_lut_LC_12_28_6 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_4_lut_LC_12_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_4_lut_LC_12_28_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx.i2_3_lut_4_lut_LC_12_28_6  (
            .in0(N__23471),
            .in1(N__23160),
            .in2(N__22481),
            .in3(N__22993),
            .lcout(n1025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_280_LC_12_28_7 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_280_LC_12_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_280_LC_12_28_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_280_LC_12_28_7  (
            .in0(N__22991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22477),
            .lcout(\c0.tx.n752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_284_LC_12_29_5 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_284_LC_12_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_284_LC_12_29_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.i1_2_lut_adj_284_LC_12_29_5  (
            .in0(_gnd_net_),
            .in1(N__22471),
            .in2(_gnd_net_),
            .in3(N__23473),
            .lcout(\c0.tx.n3643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_LC_13_26_0 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_LC_13_26_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i2_2_lut_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__23574),
            .in2(_gnd_net_),
            .in3(N__23631),
            .lcout(\c0.tx.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i2_LC_13_26_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i2_LC_13_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_13_26_1 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_13_26_1  (
            .in0(N__22604),
            .in1(N__23315),
            .in2(N__23100),
            .in3(N__23463),
            .lcout(\c0.tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22950),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_13_26_2 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_13_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_13_26_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_13_26_2  (
            .in0(N__23080),
            .in1(N__23189),
            .in2(N__23493),
            .in3(N__23013),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22950),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i6_LC_13_26_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i6_LC_13_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_13_26_5 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_13_26_5  (
            .in0(N__23558),
            .in1(N__23317),
            .in2(N__23102),
            .in3(N__23465),
            .lcout(\c0.tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22950),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i4_LC_13_26_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i4_LC_13_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_13_26_7 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_13_26_7  (
            .in0(N__23615),
            .in1(N__23316),
            .in2(N__23101),
            .in3(N__23464),
            .lcout(\c0.tx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22950),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_381_LC_13_27_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_381_LC_13_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_381_LC_13_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_381_LC_13_27_0  (
            .in0(N__22438),
            .in1(N__22390),
            .in2(_gnd_net_),
            .in3(N__22379),
            .lcout(\c0.n4477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_13_27_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i1_LC_13_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_13_27_1 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_13_27_1  (
            .in0(N__23309),
            .in1(N__22634),
            .in2(N__23099),
            .in3(N__23469),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22956),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_adj_283_LC_13_27_2 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_adj_283_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_adj_283_LC_13_27_2 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \c0.tx.i1_4_lut_adj_283_LC_13_27_2  (
            .in0(N__22593),
            .in1(N__23604),
            .in2(N__22625),
            .in3(N__22650),
            .lcout(),
            .ltout(\c0.tx.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_adj_285_LC_13_27_3 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_adj_285_LC_13_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_adj_285_LC_13_27_3 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \c0.tx.i1_4_lut_adj_285_LC_13_27_3  (
            .in0(N__23522),
            .in1(N__22568),
            .in2(N__22562),
            .in3(N__23547),
            .lcout(\c0.tx.n17 ),
            .ltout(\c0.tx.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i7_LC_13_27_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i7_LC_13_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_13_27_4 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_13_27_4  (
            .in0(N__23466),
            .in1(N__23531),
            .in2(N__22559),
            .in3(N__23314),
            .lcout(\c0.tx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22956),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_13_27_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_13_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_13_27_5 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_13_27_5  (
            .in0(N__23308),
            .in1(N__22661),
            .in2(N__23098),
            .in3(N__23468),
            .lcout(\c0.tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22956),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i5_LC_13_27_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i5_LC_13_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_13_27_6 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_13_27_6  (
            .in0(N__23078),
            .in1(N__23313),
            .in2(N__23588),
            .in3(N__23470),
            .lcout(\c0.tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22956),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i3_LC_13_27_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i3_LC_13_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_13_27_7 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_13_27_7  (
            .in0(N__22577),
            .in1(N__23467),
            .in2(N__23318),
            .in3(N__23079),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22956),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_281_LC_13_28_2 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_281_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_281_LC_13_28_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_281_LC_13_28_2  (
            .in0(_gnd_net_),
            .in1(N__23474),
            .in2(_gnd_net_),
            .in3(N__23070),
            .lcout(n4375),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i8_LC_13_28_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_13_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_13_28_6 .LUT_INIT=16'b1000100011001000;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_13_28_6  (
            .in0(N__23475),
            .in1(N__23327),
            .in2(N__23307),
            .in3(N__23071),
            .lcout(\c0.tx.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22957),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_382_LC_13_28_7 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_382_LC_13_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_382_LC_13_28_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_382_LC_13_28_7  (
            .in0(N__22556),
            .in1(N__22540),
            .in2(N__22529),
            .in3(N__22502),
            .lcout(n12_adj_944),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_13_29_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_13_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_13_29_0 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_13_29_0  (
            .in0(N__23002),
            .in1(N__23478),
            .in2(N__23200),
            .in3(N__23096),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22958),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i605_2_lut_LC_13_29_1 .C_ON=1'b0;
    defparam \c0.tx.i605_2_lut_LC_13_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i605_2_lut_LC_13_29_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i605_2_lut_LC_13_29_1  (
            .in0(_gnd_net_),
            .in1(N__23182),
            .in2(_gnd_net_),
            .in3(N__23000),
            .lcout(n88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_LC_13_29_3.C_ON=1'b0;
    defparam i1_4_lut_4_lut_LC_13_29_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_LC_13_29_3.LUT_INIT=16'b1110100011100000;
    LogicCell40 i1_4_lut_4_lut_LC_13_29_3 (
            .in0(N__23172),
            .in1(N__23001),
            .in2(N__23264),
            .in3(N__23114),
            .lcout(),
            .ltout(n4_adj_946_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Done_44_LC_13_29_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Done_44_LC_13_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Done_44_LC_13_29_4 .LUT_INIT=16'b1111100011111100;
    LogicCell40 \c0.tx.r_Tx_Done_44_LC_13_29_4  (
            .in0(N__23263),
            .in1(N__23476),
            .in2(N__23321),
            .in3(N__23306),
            .lcout(tx_done),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22958),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i25_4_lut_LC_13_29_5 .C_ON=1'b0;
    defparam \c0.tx.i25_4_lut_LC_13_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i25_4_lut_LC_13_29_5 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.tx.i25_4_lut_LC_13_29_5  (
            .in0(N__23245),
            .in1(N__23213),
            .in2(N__23193),
            .in3(N__23113),
            .lcout(),
            .ltout(\c0.tx.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_13_29_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_13_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_13_29_6 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_13_29_6  (
            .in0(N__23003),
            .in1(N__23477),
            .in2(N__23105),
            .in3(N__23097),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22958),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_14_27_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_14_27_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_2_lut_LC_14_27_0  (
            .in0(N__22673),
            .in1(N__22672),
            .in2(N__23479),
            .in3(N__22655),
            .lcout(\c0.tx.n1979 ),
            .ltout(),
            .carryin(bfn_14_27_0_),
            .carryout(\c0.tx.n3876 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_3_lut_LC_14_27_1 .C_ON=1'b1;
    defparam \c0.tx.add_59_3_lut_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_3_lut_LC_14_27_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_3_lut_LC_14_27_1  (
            .in0(N__22652),
            .in1(N__22651),
            .in2(N__23483),
            .in3(N__22628),
            .lcout(\c0.tx.n1754 ),
            .ltout(),
            .carryin(\c0.tx.n3876 ),
            .carryout(\c0.tx.n3877 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_4_lut_LC_14_27_2 .C_ON=1'b1;
    defparam \c0.tx.add_59_4_lut_LC_14_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_4_lut_LC_14_27_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_4_lut_LC_14_27_2  (
            .in0(N__22624),
            .in1(N__22623),
            .in2(N__23480),
            .in3(N__22598),
            .lcout(\c0.tx.n1751 ),
            .ltout(),
            .carryin(\c0.tx.n3877 ),
            .carryout(\c0.tx.n3878 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_5_lut_LC_14_27_3 .C_ON=1'b1;
    defparam \c0.tx.add_59_5_lut_LC_14_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_5_lut_LC_14_27_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_5_lut_LC_14_27_3  (
            .in0(N__22595),
            .in1(N__22594),
            .in2(N__23484),
            .in3(N__22571),
            .lcout(\c0.tx.n1748 ),
            .ltout(),
            .carryin(\c0.tx.n3878 ),
            .carryout(\c0.tx.n3879 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_6_lut_LC_14_27_4 .C_ON=1'b1;
    defparam \c0.tx.add_59_6_lut_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_6_lut_LC_14_27_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_6_lut_LC_14_27_4  (
            .in0(N__23633),
            .in1(N__23632),
            .in2(N__23481),
            .in3(N__23609),
            .lcout(\c0.tx.n1745 ),
            .ltout(),
            .carryin(\c0.tx.n3879 ),
            .carryout(\c0.tx.n3880 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_7_lut_LC_14_27_5 .C_ON=1'b1;
    defparam \c0.tx.add_59_7_lut_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_7_lut_LC_14_27_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_7_lut_LC_14_27_5  (
            .in0(N__23606),
            .in1(N__23605),
            .in2(N__23485),
            .in3(N__23579),
            .lcout(\c0.tx.n1742 ),
            .ltout(),
            .carryin(\c0.tx.n3880 ),
            .carryout(\c0.tx.n3881 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_8_lut_LC_14_27_6 .C_ON=1'b1;
    defparam \c0.tx.add_59_8_lut_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_8_lut_LC_14_27_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_8_lut_LC_14_27_6  (
            .in0(N__23576),
            .in1(N__23575),
            .in2(N__23482),
            .in3(N__23552),
            .lcout(\c0.tx.n1739 ),
            .ltout(),
            .carryin(\c0.tx.n3881 ),
            .carryout(\c0.tx.n3882 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_9_lut_LC_14_27_7 .C_ON=1'b1;
    defparam \c0.tx.add_59_9_lut_LC_14_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_9_lut_LC_14_27_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_9_lut_LC_14_27_7  (
            .in0(N__23549),
            .in1(N__23548),
            .in2(N__23486),
            .in3(N__23525),
            .lcout(\c0.tx.n1736 ),
            .ltout(),
            .carryin(\c0.tx.n3882 ),
            .carryout(\c0.tx.n3883 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_10_lut_LC_14_28_0 .C_ON=1'b0;
    defparam \c0.tx.add_59_10_lut_LC_14_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_10_lut_LC_14_28_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_10_lut_LC_14_28_0  (
            .in0(N__23520),
            .in1(N__23521),
            .in2(N__23494),
            .in3(N__23330),
            .lcout(\c0.tx.n1733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
