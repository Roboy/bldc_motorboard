-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 16 2019 20:28:05

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : inout std_logic;
    PIN_5 : inout std_logic;
    PIN_4 : inout std_logic;
    PIN_3 : out std_logic;
    PIN_24 : out std_logic;
    PIN_23 : out std_logic;
    PIN_22 : out std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : out std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : inout std_logic;
    PIN_10 : inout std_logic;
    PIN_1 : out std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__81286\ : std_logic;
signal \N__81285\ : std_logic;
signal \N__81284\ : std_logic;
signal \N__81277\ : std_logic;
signal \N__81276\ : std_logic;
signal \N__81275\ : std_logic;
signal \N__81268\ : std_logic;
signal \N__81267\ : std_logic;
signal \N__81266\ : std_logic;
signal \N__81259\ : std_logic;
signal \N__81258\ : std_logic;
signal \N__81257\ : std_logic;
signal \N__81250\ : std_logic;
signal \N__81249\ : std_logic;
signal \N__81248\ : std_logic;
signal \N__81241\ : std_logic;
signal \N__81240\ : std_logic;
signal \N__81239\ : std_logic;
signal \N__81232\ : std_logic;
signal \N__81231\ : std_logic;
signal \N__81230\ : std_logic;
signal \N__81223\ : std_logic;
signal \N__81222\ : std_logic;
signal \N__81221\ : std_logic;
signal \N__81214\ : std_logic;
signal \N__81213\ : std_logic;
signal \N__81212\ : std_logic;
signal \N__81205\ : std_logic;
signal \N__81204\ : std_logic;
signal \N__81203\ : std_logic;
signal \N__81196\ : std_logic;
signal \N__81195\ : std_logic;
signal \N__81194\ : std_logic;
signal \N__81187\ : std_logic;
signal \N__81186\ : std_logic;
signal \N__81185\ : std_logic;
signal \N__81178\ : std_logic;
signal \N__81177\ : std_logic;
signal \N__81176\ : std_logic;
signal \N__81169\ : std_logic;
signal \N__81168\ : std_logic;
signal \N__81167\ : std_logic;
signal \N__81160\ : std_logic;
signal \N__81159\ : std_logic;
signal \N__81158\ : std_logic;
signal \N__81151\ : std_logic;
signal \N__81150\ : std_logic;
signal \N__81149\ : std_logic;
signal \N__81142\ : std_logic;
signal \N__81141\ : std_logic;
signal \N__81140\ : std_logic;
signal \N__81133\ : std_logic;
signal \N__81132\ : std_logic;
signal \N__81131\ : std_logic;
signal \N__81114\ : std_logic;
signal \N__81111\ : std_logic;
signal \N__81108\ : std_logic;
signal \N__81105\ : std_logic;
signal \N__81104\ : std_logic;
signal \N__81103\ : std_logic;
signal \N__81100\ : std_logic;
signal \N__81097\ : std_logic;
signal \N__81094\ : std_logic;
signal \N__81091\ : std_logic;
signal \N__81086\ : std_logic;
signal \N__81081\ : std_logic;
signal \N__81078\ : std_logic;
signal \N__81075\ : std_logic;
signal \N__81072\ : std_logic;
signal \N__81071\ : std_logic;
signal \N__81068\ : std_logic;
signal \N__81065\ : std_logic;
signal \N__81062\ : std_logic;
signal \N__81059\ : std_logic;
signal \N__81058\ : std_logic;
signal \N__81057\ : std_logic;
signal \N__81054\ : std_logic;
signal \N__81051\ : std_logic;
signal \N__81048\ : std_logic;
signal \N__81045\ : std_logic;
signal \N__81042\ : std_logic;
signal \N__81039\ : std_logic;
signal \N__81036\ : std_logic;
signal \N__81033\ : std_logic;
signal \N__81032\ : std_logic;
signal \N__81031\ : std_logic;
signal \N__81028\ : std_logic;
signal \N__81025\ : std_logic;
signal \N__81020\ : std_logic;
signal \N__81015\ : std_logic;
signal \N__81006\ : std_logic;
signal \N__81003\ : std_logic;
signal \N__81002\ : std_logic;
signal \N__80999\ : std_logic;
signal \N__80996\ : std_logic;
signal \N__80991\ : std_logic;
signal \N__80988\ : std_logic;
signal \N__80987\ : std_logic;
signal \N__80986\ : std_logic;
signal \N__80983\ : std_logic;
signal \N__80982\ : std_logic;
signal \N__80979\ : std_logic;
signal \N__80976\ : std_logic;
signal \N__80975\ : std_logic;
signal \N__80974\ : std_logic;
signal \N__80973\ : std_logic;
signal \N__80970\ : std_logic;
signal \N__80967\ : std_logic;
signal \N__80966\ : std_logic;
signal \N__80963\ : std_logic;
signal \N__80960\ : std_logic;
signal \N__80957\ : std_logic;
signal \N__80952\ : std_logic;
signal \N__80951\ : std_logic;
signal \N__80948\ : std_logic;
signal \N__80945\ : std_logic;
signal \N__80944\ : std_logic;
signal \N__80943\ : std_logic;
signal \N__80942\ : std_logic;
signal \N__80941\ : std_logic;
signal \N__80940\ : std_logic;
signal \N__80937\ : std_logic;
signal \N__80928\ : std_logic;
signal \N__80925\ : std_logic;
signal \N__80924\ : std_logic;
signal \N__80923\ : std_logic;
signal \N__80922\ : std_logic;
signal \N__80921\ : std_logic;
signal \N__80920\ : std_logic;
signal \N__80919\ : std_logic;
signal \N__80918\ : std_logic;
signal \N__80913\ : std_logic;
signal \N__80908\ : std_logic;
signal \N__80905\ : std_logic;
signal \N__80900\ : std_logic;
signal \N__80899\ : std_logic;
signal \N__80894\ : std_logic;
signal \N__80889\ : std_logic;
signal \N__80888\ : std_logic;
signal \N__80885\ : std_logic;
signal \N__80882\ : std_logic;
signal \N__80875\ : std_logic;
signal \N__80872\ : std_logic;
signal \N__80871\ : std_logic;
signal \N__80868\ : std_logic;
signal \N__80867\ : std_logic;
signal \N__80864\ : std_logic;
signal \N__80859\ : std_logic;
signal \N__80856\ : std_logic;
signal \N__80853\ : std_logic;
signal \N__80850\ : std_logic;
signal \N__80847\ : std_logic;
signal \N__80844\ : std_logic;
signal \N__80843\ : std_logic;
signal \N__80840\ : std_logic;
signal \N__80837\ : std_logic;
signal \N__80834\ : std_logic;
signal \N__80831\ : std_logic;
signal \N__80828\ : std_logic;
signal \N__80825\ : std_logic;
signal \N__80820\ : std_logic;
signal \N__80813\ : std_logic;
signal \N__80810\ : std_logic;
signal \N__80807\ : std_logic;
signal \N__80804\ : std_logic;
signal \N__80799\ : std_logic;
signal \N__80796\ : std_logic;
signal \N__80793\ : std_logic;
signal \N__80790\ : std_logic;
signal \N__80787\ : std_logic;
signal \N__80784\ : std_logic;
signal \N__80781\ : std_logic;
signal \N__80776\ : std_logic;
signal \N__80769\ : std_logic;
signal \N__80764\ : std_logic;
signal \N__80757\ : std_logic;
signal \N__80748\ : std_logic;
signal \N__80747\ : std_logic;
signal \N__80746\ : std_logic;
signal \N__80743\ : std_logic;
signal \N__80742\ : std_logic;
signal \N__80741\ : std_logic;
signal \N__80740\ : std_logic;
signal \N__80739\ : std_logic;
signal \N__80738\ : std_logic;
signal \N__80737\ : std_logic;
signal \N__80736\ : std_logic;
signal \N__80735\ : std_logic;
signal \N__80734\ : std_logic;
signal \N__80733\ : std_logic;
signal \N__80730\ : std_logic;
signal \N__80729\ : std_logic;
signal \N__80726\ : std_logic;
signal \N__80723\ : std_logic;
signal \N__80720\ : std_logic;
signal \N__80719\ : std_logic;
signal \N__80718\ : std_logic;
signal \N__80715\ : std_logic;
signal \N__80712\ : std_logic;
signal \N__80711\ : std_logic;
signal \N__80708\ : std_logic;
signal \N__80707\ : std_logic;
signal \N__80704\ : std_logic;
signal \N__80703\ : std_logic;
signal \N__80700\ : std_logic;
signal \N__80697\ : std_logic;
signal \N__80696\ : std_logic;
signal \N__80693\ : std_logic;
signal \N__80688\ : std_logic;
signal \N__80685\ : std_logic;
signal \N__80682\ : std_logic;
signal \N__80679\ : std_logic;
signal \N__80674\ : std_logic;
signal \N__80673\ : std_logic;
signal \N__80672\ : std_logic;
signal \N__80671\ : std_logic;
signal \N__80668\ : std_logic;
signal \N__80665\ : std_logic;
signal \N__80662\ : std_logic;
signal \N__80659\ : std_logic;
signal \N__80656\ : std_logic;
signal \N__80655\ : std_logic;
signal \N__80650\ : std_logic;
signal \N__80647\ : std_logic;
signal \N__80644\ : std_logic;
signal \N__80641\ : std_logic;
signal \N__80638\ : std_logic;
signal \N__80635\ : std_logic;
signal \N__80632\ : std_logic;
signal \N__80627\ : std_logic;
signal \N__80624\ : std_logic;
signal \N__80619\ : std_logic;
signal \N__80618\ : std_logic;
signal \N__80617\ : std_logic;
signal \N__80616\ : std_logic;
signal \N__80615\ : std_logic;
signal \N__80612\ : std_logic;
signal \N__80609\ : std_logic;
signal \N__80606\ : std_logic;
signal \N__80605\ : std_logic;
signal \N__80602\ : std_logic;
signal \N__80595\ : std_logic;
signal \N__80592\ : std_logic;
signal \N__80589\ : std_logic;
signal \N__80586\ : std_logic;
signal \N__80581\ : std_logic;
signal \N__80576\ : std_logic;
signal \N__80575\ : std_logic;
signal \N__80568\ : std_logic;
signal \N__80565\ : std_logic;
signal \N__80562\ : std_logic;
signal \N__80557\ : std_logic;
signal \N__80554\ : std_logic;
signal \N__80549\ : std_logic;
signal \N__80546\ : std_logic;
signal \N__80543\ : std_logic;
signal \N__80540\ : std_logic;
signal \N__80535\ : std_logic;
signal \N__80532\ : std_logic;
signal \N__80527\ : std_logic;
signal \N__80524\ : std_logic;
signal \N__80521\ : std_logic;
signal \N__80518\ : std_logic;
signal \N__80515\ : std_logic;
signal \N__80510\ : std_logic;
signal \N__80509\ : std_logic;
signal \N__80508\ : std_logic;
signal \N__80505\ : std_logic;
signal \N__80502\ : std_logic;
signal \N__80497\ : std_logic;
signal \N__80492\ : std_logic;
signal \N__80487\ : std_logic;
signal \N__80484\ : std_logic;
signal \N__80481\ : std_logic;
signal \N__80478\ : std_logic;
signal \N__80471\ : std_logic;
signal \N__80466\ : std_logic;
signal \N__80463\ : std_logic;
signal \N__80458\ : std_logic;
signal \N__80453\ : std_logic;
signal \N__80444\ : std_logic;
signal \N__80433\ : std_logic;
signal \N__80432\ : std_logic;
signal \N__80431\ : std_logic;
signal \N__80430\ : std_logic;
signal \N__80429\ : std_logic;
signal \N__80428\ : std_logic;
signal \N__80427\ : std_logic;
signal \N__80426\ : std_logic;
signal \N__80425\ : std_logic;
signal \N__80424\ : std_logic;
signal \N__80423\ : std_logic;
signal \N__80422\ : std_logic;
signal \N__80421\ : std_logic;
signal \N__80420\ : std_logic;
signal \N__80419\ : std_logic;
signal \N__80418\ : std_logic;
signal \N__80417\ : std_logic;
signal \N__80416\ : std_logic;
signal \N__80415\ : std_logic;
signal \N__80414\ : std_logic;
signal \N__80413\ : std_logic;
signal \N__80412\ : std_logic;
signal \N__80407\ : std_logic;
signal \N__80404\ : std_logic;
signal \N__80403\ : std_logic;
signal \N__80402\ : std_logic;
signal \N__80401\ : std_logic;
signal \N__80400\ : std_logic;
signal \N__80399\ : std_logic;
signal \N__80398\ : std_logic;
signal \N__80397\ : std_logic;
signal \N__80396\ : std_logic;
signal \N__80395\ : std_logic;
signal \N__80392\ : std_logic;
signal \N__80389\ : std_logic;
signal \N__80386\ : std_logic;
signal \N__80385\ : std_logic;
signal \N__80382\ : std_logic;
signal \N__80379\ : std_logic;
signal \N__80376\ : std_logic;
signal \N__80373\ : std_logic;
signal \N__80368\ : std_logic;
signal \N__80365\ : std_logic;
signal \N__80360\ : std_logic;
signal \N__80355\ : std_logic;
signal \N__80344\ : std_logic;
signal \N__80341\ : std_logic;
signal \N__80338\ : std_logic;
signal \N__80329\ : std_logic;
signal \N__80328\ : std_logic;
signal \N__80325\ : std_logic;
signal \N__80324\ : std_logic;
signal \N__80323\ : std_logic;
signal \N__80322\ : std_logic;
signal \N__80321\ : std_logic;
signal \N__80320\ : std_logic;
signal \N__80319\ : std_logic;
signal \N__80318\ : std_logic;
signal \N__80315\ : std_logic;
signal \N__80312\ : std_logic;
signal \N__80307\ : std_logic;
signal \N__80304\ : std_logic;
signal \N__80299\ : std_logic;
signal \N__80296\ : std_logic;
signal \N__80293\ : std_logic;
signal \N__80288\ : std_logic;
signal \N__80283\ : std_logic;
signal \N__80276\ : std_logic;
signal \N__80267\ : std_logic;
signal \N__80266\ : std_logic;
signal \N__80265\ : std_logic;
signal \N__80264\ : std_logic;
signal \N__80263\ : std_logic;
signal \N__80262\ : std_logic;
signal \N__80261\ : std_logic;
signal \N__80260\ : std_logic;
signal \N__80259\ : std_logic;
signal \N__80256\ : std_logic;
signal \N__80253\ : std_logic;
signal \N__80250\ : std_logic;
signal \N__80241\ : std_logic;
signal \N__80236\ : std_logic;
signal \N__80233\ : std_logic;
signal \N__80230\ : std_logic;
signal \N__80227\ : std_logic;
signal \N__80224\ : std_logic;
signal \N__80221\ : std_logic;
signal \N__80218\ : std_logic;
signal \N__80213\ : std_logic;
signal \N__80206\ : std_logic;
signal \N__80203\ : std_logic;
signal \N__80200\ : std_logic;
signal \N__80197\ : std_logic;
signal \N__80186\ : std_logic;
signal \N__80183\ : std_logic;
signal \N__80180\ : std_logic;
signal \N__80171\ : std_logic;
signal \N__80162\ : std_logic;
signal \N__80155\ : std_logic;
signal \N__80136\ : std_logic;
signal \N__80135\ : std_logic;
signal \N__80132\ : std_logic;
signal \N__80131\ : std_logic;
signal \N__80128\ : std_logic;
signal \N__80125\ : std_logic;
signal \N__80122\ : std_logic;
signal \N__80119\ : std_logic;
signal \N__80116\ : std_logic;
signal \N__80113\ : std_logic;
signal \N__80110\ : std_logic;
signal \N__80107\ : std_logic;
signal \N__80100\ : std_logic;
signal \N__80099\ : std_logic;
signal \N__80098\ : std_logic;
signal \N__80097\ : std_logic;
signal \N__80096\ : std_logic;
signal \N__80095\ : std_logic;
signal \N__80094\ : std_logic;
signal \N__80093\ : std_logic;
signal \N__80090\ : std_logic;
signal \N__80087\ : std_logic;
signal \N__80084\ : std_logic;
signal \N__80081\ : std_logic;
signal \N__80080\ : std_logic;
signal \N__80079\ : std_logic;
signal \N__80076\ : std_logic;
signal \N__80073\ : std_logic;
signal \N__80070\ : std_logic;
signal \N__80067\ : std_logic;
signal \N__80064\ : std_logic;
signal \N__80061\ : std_logic;
signal \N__80060\ : std_logic;
signal \N__80055\ : std_logic;
signal \N__80052\ : std_logic;
signal \N__80051\ : std_logic;
signal \N__80048\ : std_logic;
signal \N__80045\ : std_logic;
signal \N__80044\ : std_logic;
signal \N__80041\ : std_logic;
signal \N__80036\ : std_logic;
signal \N__80033\ : std_logic;
signal \N__80032\ : std_logic;
signal \N__80031\ : std_logic;
signal \N__80030\ : std_logic;
signal \N__80029\ : std_logic;
signal \N__80026\ : std_logic;
signal \N__80023\ : std_logic;
signal \N__80020\ : std_logic;
signal \N__80017\ : std_logic;
signal \N__80016\ : std_logic;
signal \N__80013\ : std_logic;
signal \N__80010\ : std_logic;
signal \N__80009\ : std_logic;
signal \N__80008\ : std_logic;
signal \N__80007\ : std_logic;
signal \N__80004\ : std_logic;
signal \N__80001\ : std_logic;
signal \N__79998\ : std_logic;
signal \N__79995\ : std_logic;
signal \N__79992\ : std_logic;
signal \N__79989\ : std_logic;
signal \N__79988\ : std_logic;
signal \N__79987\ : std_logic;
signal \N__79986\ : std_logic;
signal \N__79985\ : std_logic;
signal \N__79984\ : std_logic;
signal \N__79983\ : std_logic;
signal \N__79980\ : std_logic;
signal \N__79975\ : std_logic;
signal \N__79972\ : std_logic;
signal \N__79967\ : std_logic;
signal \N__79964\ : std_logic;
signal \N__79961\ : std_logic;
signal \N__79958\ : std_logic;
signal \N__79955\ : std_logic;
signal \N__79954\ : std_logic;
signal \N__79953\ : std_logic;
signal \N__79952\ : std_logic;
signal \N__79949\ : std_logic;
signal \N__79948\ : std_logic;
signal \N__79947\ : std_logic;
signal \N__79944\ : std_logic;
signal \N__79941\ : std_logic;
signal \N__79938\ : std_logic;
signal \N__79929\ : std_logic;
signal \N__79922\ : std_logic;
signal \N__79919\ : std_logic;
signal \N__79914\ : std_logic;
signal \N__79911\ : std_logic;
signal \N__79908\ : std_logic;
signal \N__79901\ : std_logic;
signal \N__79892\ : std_logic;
signal \N__79889\ : std_logic;
signal \N__79886\ : std_logic;
signal \N__79883\ : std_logic;
signal \N__79878\ : std_logic;
signal \N__79875\ : std_logic;
signal \N__79868\ : std_logic;
signal \N__79865\ : std_logic;
signal \N__79860\ : std_logic;
signal \N__79857\ : std_logic;
signal \N__79848\ : std_logic;
signal \N__79845\ : std_logic;
signal \N__79842\ : std_logic;
signal \N__79833\ : std_logic;
signal \N__79830\ : std_logic;
signal \N__79827\ : std_logic;
signal \N__79824\ : std_logic;
signal \N__79821\ : std_logic;
signal \N__79814\ : std_logic;
signal \N__79811\ : std_logic;
signal \N__79800\ : std_logic;
signal \N__79797\ : std_logic;
signal \N__79796\ : std_logic;
signal \N__79793\ : std_logic;
signal \N__79792\ : std_logic;
signal \N__79791\ : std_logic;
signal \N__79788\ : std_logic;
signal \N__79787\ : std_logic;
signal \N__79786\ : std_logic;
signal \N__79785\ : std_logic;
signal \N__79784\ : std_logic;
signal \N__79781\ : std_logic;
signal \N__79778\ : std_logic;
signal \N__79777\ : std_logic;
signal \N__79776\ : std_logic;
signal \N__79769\ : std_logic;
signal \N__79766\ : std_logic;
signal \N__79763\ : std_logic;
signal \N__79760\ : std_logic;
signal \N__79759\ : std_logic;
signal \N__79758\ : std_logic;
signal \N__79757\ : std_logic;
signal \N__79756\ : std_logic;
signal \N__79751\ : std_logic;
signal \N__79746\ : std_logic;
signal \N__79743\ : std_logic;
signal \N__79740\ : std_logic;
signal \N__79737\ : std_logic;
signal \N__79734\ : std_logic;
signal \N__79729\ : std_logic;
signal \N__79728\ : std_logic;
signal \N__79727\ : std_logic;
signal \N__79724\ : std_logic;
signal \N__79721\ : std_logic;
signal \N__79718\ : std_logic;
signal \N__79709\ : std_logic;
signal \N__79704\ : std_logic;
signal \N__79703\ : std_logic;
signal \N__79702\ : std_logic;
signal \N__79699\ : std_logic;
signal \N__79698\ : std_logic;
signal \N__79695\ : std_logic;
signal \N__79692\ : std_logic;
signal \N__79689\ : std_logic;
signal \N__79686\ : std_logic;
signal \N__79681\ : std_logic;
signal \N__79678\ : std_logic;
signal \N__79677\ : std_logic;
signal \N__79674\ : std_logic;
signal \N__79671\ : std_logic;
signal \N__79668\ : std_logic;
signal \N__79665\ : std_logic;
signal \N__79662\ : std_logic;
signal \N__79653\ : std_logic;
signal \N__79650\ : std_logic;
signal \N__79649\ : std_logic;
signal \N__79648\ : std_logic;
signal \N__79647\ : std_logic;
signal \N__79646\ : std_logic;
signal \N__79641\ : std_logic;
signal \N__79632\ : std_logic;
signal \N__79629\ : std_logic;
signal \N__79628\ : std_logic;
signal \N__79627\ : std_logic;
signal \N__79626\ : std_logic;
signal \N__79623\ : std_logic;
signal \N__79622\ : std_logic;
signal \N__79619\ : std_logic;
signal \N__79616\ : std_logic;
signal \N__79613\ : std_logic;
signal \N__79608\ : std_logic;
signal \N__79605\ : std_logic;
signal \N__79602\ : std_logic;
signal \N__79599\ : std_logic;
signal \N__79596\ : std_logic;
signal \N__79593\ : std_logic;
signal \N__79590\ : std_logic;
signal \N__79589\ : std_logic;
signal \N__79588\ : std_logic;
signal \N__79587\ : std_logic;
signal \N__79582\ : std_logic;
signal \N__79579\ : std_logic;
signal \N__79576\ : std_logic;
signal \N__79571\ : std_logic;
signal \N__79568\ : std_logic;
signal \N__79565\ : std_logic;
signal \N__79560\ : std_logic;
signal \N__79557\ : std_logic;
signal \N__79554\ : std_logic;
signal \N__79551\ : std_logic;
signal \N__79548\ : std_logic;
signal \N__79543\ : std_logic;
signal \N__79542\ : std_logic;
signal \N__79537\ : std_logic;
signal \N__79532\ : std_logic;
signal \N__79527\ : std_logic;
signal \N__79522\ : std_logic;
signal \N__79519\ : std_logic;
signal \N__79516\ : std_logic;
signal \N__79513\ : std_logic;
signal \N__79510\ : std_logic;
signal \N__79505\ : std_logic;
signal \N__79502\ : std_logic;
signal \N__79491\ : std_logic;
signal \N__79490\ : std_logic;
signal \N__79489\ : std_logic;
signal \N__79488\ : std_logic;
signal \N__79485\ : std_logic;
signal \N__79484\ : std_logic;
signal \N__79483\ : std_logic;
signal \N__79482\ : std_logic;
signal \N__79481\ : std_logic;
signal \N__79478\ : std_logic;
signal \N__79477\ : std_logic;
signal \N__79476\ : std_logic;
signal \N__79473\ : std_logic;
signal \N__79472\ : std_logic;
signal \N__79471\ : std_logic;
signal \N__79468\ : std_logic;
signal \N__79465\ : std_logic;
signal \N__79464\ : std_logic;
signal \N__79463\ : std_logic;
signal \N__79458\ : std_logic;
signal \N__79457\ : std_logic;
signal \N__79456\ : std_logic;
signal \N__79453\ : std_logic;
signal \N__79450\ : std_logic;
signal \N__79447\ : std_logic;
signal \N__79444\ : std_logic;
signal \N__79443\ : std_logic;
signal \N__79442\ : std_logic;
signal \N__79441\ : std_logic;
signal \N__79440\ : std_logic;
signal \N__79439\ : std_logic;
signal \N__79436\ : std_logic;
signal \N__79433\ : std_logic;
signal \N__79428\ : std_logic;
signal \N__79425\ : std_logic;
signal \N__79422\ : std_logic;
signal \N__79421\ : std_logic;
signal \N__79420\ : std_logic;
signal \N__79415\ : std_logic;
signal \N__79412\ : std_logic;
signal \N__79407\ : std_logic;
signal \N__79404\ : std_logic;
signal \N__79399\ : std_logic;
signal \N__79398\ : std_logic;
signal \N__79397\ : std_logic;
signal \N__79396\ : std_logic;
signal \N__79393\ : std_logic;
signal \N__79388\ : std_logic;
signal \N__79385\ : std_logic;
signal \N__79380\ : std_logic;
signal \N__79373\ : std_logic;
signal \N__79370\ : std_logic;
signal \N__79367\ : std_logic;
signal \N__79366\ : std_logic;
signal \N__79365\ : std_logic;
signal \N__79364\ : std_logic;
signal \N__79363\ : std_logic;
signal \N__79362\ : std_logic;
signal \N__79361\ : std_logic;
signal \N__79360\ : std_logic;
signal \N__79359\ : std_logic;
signal \N__79358\ : std_logic;
signal \N__79357\ : std_logic;
signal \N__79356\ : std_logic;
signal \N__79355\ : std_logic;
signal \N__79354\ : std_logic;
signal \N__79351\ : std_logic;
signal \N__79348\ : std_logic;
signal \N__79345\ : std_logic;
signal \N__79342\ : std_logic;
signal \N__79337\ : std_logic;
signal \N__79334\ : std_logic;
signal \N__79327\ : std_logic;
signal \N__79324\ : std_logic;
signal \N__79321\ : std_logic;
signal \N__79316\ : std_logic;
signal \N__79311\ : std_logic;
signal \N__79308\ : std_logic;
signal \N__79305\ : std_logic;
signal \N__79300\ : std_logic;
signal \N__79295\ : std_logic;
signal \N__79288\ : std_logic;
signal \N__79277\ : std_logic;
signal \N__79274\ : std_logic;
signal \N__79269\ : std_logic;
signal \N__79266\ : std_logic;
signal \N__79261\ : std_logic;
signal \N__79248\ : std_logic;
signal \N__79227\ : std_logic;
signal \N__79226\ : std_logic;
signal \N__79223\ : std_logic;
signal \N__79220\ : std_logic;
signal \N__79217\ : std_logic;
signal \N__79214\ : std_logic;
signal \N__79209\ : std_logic;
signal \N__79206\ : std_logic;
signal \N__79205\ : std_logic;
signal \N__79204\ : std_logic;
signal \N__79203\ : std_logic;
signal \N__79200\ : std_logic;
signal \N__79197\ : std_logic;
signal \N__79194\ : std_logic;
signal \N__79193\ : std_logic;
signal \N__79192\ : std_logic;
signal \N__79191\ : std_logic;
signal \N__79190\ : std_logic;
signal \N__79189\ : std_logic;
signal \N__79186\ : std_logic;
signal \N__79185\ : std_logic;
signal \N__79184\ : std_logic;
signal \N__79183\ : std_logic;
signal \N__79182\ : std_logic;
signal \N__79177\ : std_logic;
signal \N__79174\ : std_logic;
signal \N__79173\ : std_logic;
signal \N__79172\ : std_logic;
signal \N__79169\ : std_logic;
signal \N__79168\ : std_logic;
signal \N__79167\ : std_logic;
signal \N__79164\ : std_logic;
signal \N__79161\ : std_logic;
signal \N__79158\ : std_logic;
signal \N__79155\ : std_logic;
signal \N__79152\ : std_logic;
signal \N__79149\ : std_logic;
signal \N__79148\ : std_logic;
signal \N__79145\ : std_logic;
signal \N__79142\ : std_logic;
signal \N__79141\ : std_logic;
signal \N__79140\ : std_logic;
signal \N__79137\ : std_logic;
signal \N__79132\ : std_logic;
signal \N__79129\ : std_logic;
signal \N__79126\ : std_logic;
signal \N__79125\ : std_logic;
signal \N__79120\ : std_logic;
signal \N__79117\ : std_logic;
signal \N__79114\ : std_logic;
signal \N__79111\ : std_logic;
signal \N__79110\ : std_logic;
signal \N__79109\ : std_logic;
signal \N__79108\ : std_logic;
signal \N__79107\ : std_logic;
signal \N__79106\ : std_logic;
signal \N__79101\ : std_logic;
signal \N__79096\ : std_logic;
signal \N__79093\ : std_logic;
signal \N__79088\ : std_logic;
signal \N__79085\ : std_logic;
signal \N__79084\ : std_logic;
signal \N__79083\ : std_logic;
signal \N__79078\ : std_logic;
signal \N__79075\ : std_logic;
signal \N__79072\ : std_logic;
signal \N__79069\ : std_logic;
signal \N__79066\ : std_logic;
signal \N__79063\ : std_logic;
signal \N__79060\ : std_logic;
signal \N__79055\ : std_logic;
signal \N__79052\ : std_logic;
signal \N__79051\ : std_logic;
signal \N__79046\ : std_logic;
signal \N__79043\ : std_logic;
signal \N__79040\ : std_logic;
signal \N__79037\ : std_logic;
signal \N__79034\ : std_logic;
signal \N__79029\ : std_logic;
signal \N__79022\ : std_logic;
signal \N__79019\ : std_logic;
signal \N__79016\ : std_logic;
signal \N__79009\ : std_logic;
signal \N__79006\ : std_logic;
signal \N__79001\ : std_logic;
signal \N__78998\ : std_logic;
signal \N__78995\ : std_logic;
signal \N__78994\ : std_logic;
signal \N__78985\ : std_logic;
signal \N__78980\ : std_logic;
signal \N__78979\ : std_logic;
signal \N__78978\ : std_logic;
signal \N__78975\ : std_logic;
signal \N__78970\ : std_logic;
signal \N__78963\ : std_logic;
signal \N__78960\ : std_logic;
signal \N__78955\ : std_logic;
signal \N__78952\ : std_logic;
signal \N__78949\ : std_logic;
signal \N__78946\ : std_logic;
signal \N__78943\ : std_logic;
signal \N__78938\ : std_logic;
signal \N__78933\ : std_logic;
signal \N__78926\ : std_logic;
signal \N__78915\ : std_logic;
signal \N__78912\ : std_logic;
signal \N__78911\ : std_logic;
signal \N__78908\ : std_logic;
signal \N__78905\ : std_logic;
signal \N__78904\ : std_logic;
signal \N__78901\ : std_logic;
signal \N__78898\ : std_logic;
signal \N__78897\ : std_logic;
signal \N__78896\ : std_logic;
signal \N__78895\ : std_logic;
signal \N__78892\ : std_logic;
signal \N__78891\ : std_logic;
signal \N__78890\ : std_logic;
signal \N__78887\ : std_logic;
signal \N__78884\ : std_logic;
signal \N__78881\ : std_logic;
signal \N__78876\ : std_logic;
signal \N__78873\ : std_logic;
signal \N__78870\ : std_logic;
signal \N__78867\ : std_logic;
signal \N__78852\ : std_logic;
signal \N__78849\ : std_logic;
signal \N__78846\ : std_logic;
signal \N__78843\ : std_logic;
signal \N__78842\ : std_logic;
signal \N__78841\ : std_logic;
signal \N__78838\ : std_logic;
signal \N__78833\ : std_logic;
signal \N__78830\ : std_logic;
signal \N__78825\ : std_logic;
signal \N__78824\ : std_logic;
signal \N__78823\ : std_logic;
signal \N__78822\ : std_logic;
signal \N__78821\ : std_logic;
signal \N__78820\ : std_logic;
signal \N__78819\ : std_logic;
signal \N__78818\ : std_logic;
signal \N__78817\ : std_logic;
signal \N__78816\ : std_logic;
signal \N__78815\ : std_logic;
signal \N__78814\ : std_logic;
signal \N__78813\ : std_logic;
signal \N__78812\ : std_logic;
signal \N__78811\ : std_logic;
signal \N__78810\ : std_logic;
signal \N__78809\ : std_logic;
signal \N__78808\ : std_logic;
signal \N__78807\ : std_logic;
signal \N__78806\ : std_logic;
signal \N__78805\ : std_logic;
signal \N__78804\ : std_logic;
signal \N__78803\ : std_logic;
signal \N__78802\ : std_logic;
signal \N__78801\ : std_logic;
signal \N__78800\ : std_logic;
signal \N__78799\ : std_logic;
signal \N__78798\ : std_logic;
signal \N__78797\ : std_logic;
signal \N__78796\ : std_logic;
signal \N__78795\ : std_logic;
signal \N__78794\ : std_logic;
signal \N__78793\ : std_logic;
signal \N__78792\ : std_logic;
signal \N__78791\ : std_logic;
signal \N__78790\ : std_logic;
signal \N__78789\ : std_logic;
signal \N__78788\ : std_logic;
signal \N__78787\ : std_logic;
signal \N__78786\ : std_logic;
signal \N__78785\ : std_logic;
signal \N__78784\ : std_logic;
signal \N__78783\ : std_logic;
signal \N__78782\ : std_logic;
signal \N__78781\ : std_logic;
signal \N__78780\ : std_logic;
signal \N__78779\ : std_logic;
signal \N__78778\ : std_logic;
signal \N__78777\ : std_logic;
signal \N__78776\ : std_logic;
signal \N__78775\ : std_logic;
signal \N__78774\ : std_logic;
signal \N__78773\ : std_logic;
signal \N__78772\ : std_logic;
signal \N__78771\ : std_logic;
signal \N__78770\ : std_logic;
signal \N__78769\ : std_logic;
signal \N__78768\ : std_logic;
signal \N__78767\ : std_logic;
signal \N__78766\ : std_logic;
signal \N__78765\ : std_logic;
signal \N__78764\ : std_logic;
signal \N__78763\ : std_logic;
signal \N__78762\ : std_logic;
signal \N__78761\ : std_logic;
signal \N__78760\ : std_logic;
signal \N__78759\ : std_logic;
signal \N__78758\ : std_logic;
signal \N__78757\ : std_logic;
signal \N__78756\ : std_logic;
signal \N__78755\ : std_logic;
signal \N__78754\ : std_logic;
signal \N__78753\ : std_logic;
signal \N__78752\ : std_logic;
signal \N__78751\ : std_logic;
signal \N__78750\ : std_logic;
signal \N__78749\ : std_logic;
signal \N__78748\ : std_logic;
signal \N__78747\ : std_logic;
signal \N__78746\ : std_logic;
signal \N__78745\ : std_logic;
signal \N__78744\ : std_logic;
signal \N__78743\ : std_logic;
signal \N__78742\ : std_logic;
signal \N__78741\ : std_logic;
signal \N__78740\ : std_logic;
signal \N__78739\ : std_logic;
signal \N__78738\ : std_logic;
signal \N__78737\ : std_logic;
signal \N__78736\ : std_logic;
signal \N__78735\ : std_logic;
signal \N__78734\ : std_logic;
signal \N__78733\ : std_logic;
signal \N__78732\ : std_logic;
signal \N__78731\ : std_logic;
signal \N__78730\ : std_logic;
signal \N__78729\ : std_logic;
signal \N__78728\ : std_logic;
signal \N__78727\ : std_logic;
signal \N__78726\ : std_logic;
signal \N__78725\ : std_logic;
signal \N__78724\ : std_logic;
signal \N__78723\ : std_logic;
signal \N__78722\ : std_logic;
signal \N__78721\ : std_logic;
signal \N__78720\ : std_logic;
signal \N__78719\ : std_logic;
signal \N__78718\ : std_logic;
signal \N__78717\ : std_logic;
signal \N__78716\ : std_logic;
signal \N__78715\ : std_logic;
signal \N__78714\ : std_logic;
signal \N__78713\ : std_logic;
signal \N__78712\ : std_logic;
signal \N__78711\ : std_logic;
signal \N__78710\ : std_logic;
signal \N__78709\ : std_logic;
signal \N__78708\ : std_logic;
signal \N__78707\ : std_logic;
signal \N__78706\ : std_logic;
signal \N__78705\ : std_logic;
signal \N__78704\ : std_logic;
signal \N__78703\ : std_logic;
signal \N__78702\ : std_logic;
signal \N__78701\ : std_logic;
signal \N__78700\ : std_logic;
signal \N__78699\ : std_logic;
signal \N__78698\ : std_logic;
signal \N__78697\ : std_logic;
signal \N__78696\ : std_logic;
signal \N__78695\ : std_logic;
signal \N__78694\ : std_logic;
signal \N__78693\ : std_logic;
signal \N__78692\ : std_logic;
signal \N__78691\ : std_logic;
signal \N__78690\ : std_logic;
signal \N__78689\ : std_logic;
signal \N__78688\ : std_logic;
signal \N__78687\ : std_logic;
signal \N__78686\ : std_logic;
signal \N__78685\ : std_logic;
signal \N__78684\ : std_logic;
signal \N__78683\ : std_logic;
signal \N__78682\ : std_logic;
signal \N__78681\ : std_logic;
signal \N__78680\ : std_logic;
signal \N__78679\ : std_logic;
signal \N__78678\ : std_logic;
signal \N__78677\ : std_logic;
signal \N__78676\ : std_logic;
signal \N__78675\ : std_logic;
signal \N__78674\ : std_logic;
signal \N__78673\ : std_logic;
signal \N__78672\ : std_logic;
signal \N__78671\ : std_logic;
signal \N__78670\ : std_logic;
signal \N__78669\ : std_logic;
signal \N__78668\ : std_logic;
signal \N__78667\ : std_logic;
signal \N__78666\ : std_logic;
signal \N__78665\ : std_logic;
signal \N__78664\ : std_logic;
signal \N__78663\ : std_logic;
signal \N__78662\ : std_logic;
signal \N__78661\ : std_logic;
signal \N__78660\ : std_logic;
signal \N__78659\ : std_logic;
signal \N__78658\ : std_logic;
signal \N__78657\ : std_logic;
signal \N__78656\ : std_logic;
signal \N__78655\ : std_logic;
signal \N__78654\ : std_logic;
signal \N__78653\ : std_logic;
signal \N__78652\ : std_logic;
signal \N__78651\ : std_logic;
signal \N__78650\ : std_logic;
signal \N__78649\ : std_logic;
signal \N__78648\ : std_logic;
signal \N__78647\ : std_logic;
signal \N__78646\ : std_logic;
signal \N__78645\ : std_logic;
signal \N__78644\ : std_logic;
signal \N__78643\ : std_logic;
signal \N__78642\ : std_logic;
signal \N__78641\ : std_logic;
signal \N__78640\ : std_logic;
signal \N__78639\ : std_logic;
signal \N__78638\ : std_logic;
signal \N__78637\ : std_logic;
signal \N__78636\ : std_logic;
signal \N__78635\ : std_logic;
signal \N__78634\ : std_logic;
signal \N__78633\ : std_logic;
signal \N__78632\ : std_logic;
signal \N__78631\ : std_logic;
signal \N__78630\ : std_logic;
signal \N__78629\ : std_logic;
signal \N__78628\ : std_logic;
signal \N__78627\ : std_logic;
signal \N__78626\ : std_logic;
signal \N__78625\ : std_logic;
signal \N__78624\ : std_logic;
signal \N__78623\ : std_logic;
signal \N__78622\ : std_logic;
signal \N__78621\ : std_logic;
signal \N__78620\ : std_logic;
signal \N__78619\ : std_logic;
signal \N__78618\ : std_logic;
signal \N__78617\ : std_logic;
signal \N__78616\ : std_logic;
signal \N__78615\ : std_logic;
signal \N__78614\ : std_logic;
signal \N__78613\ : std_logic;
signal \N__78612\ : std_logic;
signal \N__78611\ : std_logic;
signal \N__78610\ : std_logic;
signal \N__78609\ : std_logic;
signal \N__78608\ : std_logic;
signal \N__78607\ : std_logic;
signal \N__78606\ : std_logic;
signal \N__78605\ : std_logic;
signal \N__78604\ : std_logic;
signal \N__78603\ : std_logic;
signal \N__78602\ : std_logic;
signal \N__78601\ : std_logic;
signal \N__78600\ : std_logic;
signal \N__78599\ : std_logic;
signal \N__78598\ : std_logic;
signal \N__78597\ : std_logic;
signal \N__78596\ : std_logic;
signal \N__78595\ : std_logic;
signal \N__78594\ : std_logic;
signal \N__78593\ : std_logic;
signal \N__78592\ : std_logic;
signal \N__78591\ : std_logic;
signal \N__78590\ : std_logic;
signal \N__78589\ : std_logic;
signal \N__78588\ : std_logic;
signal \N__78587\ : std_logic;
signal \N__78586\ : std_logic;
signal \N__78585\ : std_logic;
signal \N__78584\ : std_logic;
signal \N__78583\ : std_logic;
signal \N__78582\ : std_logic;
signal \N__78581\ : std_logic;
signal \N__78580\ : std_logic;
signal \N__78579\ : std_logic;
signal \N__78578\ : std_logic;
signal \N__78577\ : std_logic;
signal \N__78576\ : std_logic;
signal \N__78575\ : std_logic;
signal \N__78574\ : std_logic;
signal \N__78573\ : std_logic;
signal \N__78572\ : std_logic;
signal \N__78571\ : std_logic;
signal \N__78570\ : std_logic;
signal \N__78569\ : std_logic;
signal \N__78568\ : std_logic;
signal \N__78567\ : std_logic;
signal \N__78566\ : std_logic;
signal \N__78565\ : std_logic;
signal \N__78564\ : std_logic;
signal \N__78563\ : std_logic;
signal \N__78562\ : std_logic;
signal \N__78033\ : std_logic;
signal \N__78030\ : std_logic;
signal \N__78027\ : std_logic;
signal \N__78026\ : std_logic;
signal \N__78025\ : std_logic;
signal \N__78024\ : std_logic;
signal \N__78021\ : std_logic;
signal \N__78020\ : std_logic;
signal \N__78019\ : std_logic;
signal \N__78018\ : std_logic;
signal \N__78017\ : std_logic;
signal \N__78014\ : std_logic;
signal \N__78009\ : std_logic;
signal \N__78006\ : std_logic;
signal \N__78003\ : std_logic;
signal \N__77998\ : std_logic;
signal \N__77995\ : std_logic;
signal \N__77992\ : std_logic;
signal \N__77987\ : std_logic;
signal \N__77982\ : std_logic;
signal \N__77979\ : std_logic;
signal \N__77976\ : std_logic;
signal \N__77971\ : std_logic;
signal \N__77966\ : std_logic;
signal \N__77963\ : std_logic;
signal \N__77958\ : std_logic;
signal \N__77957\ : std_logic;
signal \N__77956\ : std_logic;
signal \N__77955\ : std_logic;
signal \N__77954\ : std_logic;
signal \N__77951\ : std_logic;
signal \N__77948\ : std_logic;
signal \N__77945\ : std_logic;
signal \N__77942\ : std_logic;
signal \N__77939\ : std_logic;
signal \N__77938\ : std_logic;
signal \N__77933\ : std_logic;
signal \N__77928\ : std_logic;
signal \N__77925\ : std_logic;
signal \N__77922\ : std_logic;
signal \N__77919\ : std_logic;
signal \N__77914\ : std_logic;
signal \N__77911\ : std_logic;
signal \N__77906\ : std_logic;
signal \N__77903\ : std_logic;
signal \N__77898\ : std_logic;
signal \N__77895\ : std_logic;
signal \N__77892\ : std_logic;
signal \N__77889\ : std_logic;
signal \N__77886\ : std_logic;
signal \N__77883\ : std_logic;
signal \N__77880\ : std_logic;
signal \N__77879\ : std_logic;
signal \N__77876\ : std_logic;
signal \N__77873\ : std_logic;
signal \N__77872\ : std_logic;
signal \N__77869\ : std_logic;
signal \N__77866\ : std_logic;
signal \N__77863\ : std_logic;
signal \N__77858\ : std_logic;
signal \N__77857\ : std_logic;
signal \N__77856\ : std_logic;
signal \N__77853\ : std_logic;
signal \N__77850\ : std_logic;
signal \N__77847\ : std_logic;
signal \N__77846\ : std_logic;
signal \N__77845\ : std_logic;
signal \N__77844\ : std_logic;
signal \N__77841\ : std_logic;
signal \N__77838\ : std_logic;
signal \N__77833\ : std_logic;
signal \N__77826\ : std_logic;
signal \N__77817\ : std_logic;
signal \N__77816\ : std_logic;
signal \N__77813\ : std_logic;
signal \N__77812\ : std_logic;
signal \N__77811\ : std_logic;
signal \N__77810\ : std_logic;
signal \N__77807\ : std_logic;
signal \N__77804\ : std_logic;
signal \N__77799\ : std_logic;
signal \N__77796\ : std_logic;
signal \N__77793\ : std_logic;
signal \N__77792\ : std_logic;
signal \N__77789\ : std_logic;
signal \N__77784\ : std_logic;
signal \N__77781\ : std_logic;
signal \N__77778\ : std_logic;
signal \N__77777\ : std_logic;
signal \N__77776\ : std_logic;
signal \N__77771\ : std_logic;
signal \N__77766\ : std_logic;
signal \N__77761\ : std_logic;
signal \N__77754\ : std_logic;
signal \N__77751\ : std_logic;
signal \N__77748\ : std_logic;
signal \N__77745\ : std_logic;
signal \N__77742\ : std_logic;
signal \N__77739\ : std_logic;
signal \N__77736\ : std_logic;
signal \N__77733\ : std_logic;
signal \N__77730\ : std_logic;
signal \N__77727\ : std_logic;
signal \N__77726\ : std_logic;
signal \N__77723\ : std_logic;
signal \N__77720\ : std_logic;
signal \N__77715\ : std_logic;
signal \N__77712\ : std_logic;
signal \N__77709\ : std_logic;
signal \N__77706\ : std_logic;
signal \N__77705\ : std_logic;
signal \N__77702\ : std_logic;
signal \N__77699\ : std_logic;
signal \N__77696\ : std_logic;
signal \N__77693\ : std_logic;
signal \N__77688\ : std_logic;
signal \N__77687\ : std_logic;
signal \N__77684\ : std_logic;
signal \N__77681\ : std_logic;
signal \N__77678\ : std_logic;
signal \N__77675\ : std_logic;
signal \N__77674\ : std_logic;
signal \N__77673\ : std_logic;
signal \N__77668\ : std_logic;
signal \N__77663\ : std_logic;
signal \N__77658\ : std_logic;
signal \N__77655\ : std_logic;
signal \N__77654\ : std_logic;
signal \N__77651\ : std_logic;
signal \N__77650\ : std_logic;
signal \N__77649\ : std_logic;
signal \N__77646\ : std_logic;
signal \N__77643\ : std_logic;
signal \N__77640\ : std_logic;
signal \N__77639\ : std_logic;
signal \N__77638\ : std_logic;
signal \N__77635\ : std_logic;
signal \N__77632\ : std_logic;
signal \N__77629\ : std_logic;
signal \N__77626\ : std_logic;
signal \N__77623\ : std_logic;
signal \N__77620\ : std_logic;
signal \N__77617\ : std_logic;
signal \N__77614\ : std_logic;
signal \N__77611\ : std_logic;
signal \N__77608\ : std_logic;
signal \N__77605\ : std_logic;
signal \N__77602\ : std_logic;
signal \N__77593\ : std_logic;
signal \N__77590\ : std_logic;
signal \N__77583\ : std_logic;
signal \N__77580\ : std_logic;
signal \N__77579\ : std_logic;
signal \N__77578\ : std_logic;
signal \N__77575\ : std_logic;
signal \N__77574\ : std_logic;
signal \N__77573\ : std_logic;
signal \N__77570\ : std_logic;
signal \N__77569\ : std_logic;
signal \N__77566\ : std_logic;
signal \N__77563\ : std_logic;
signal \N__77560\ : std_logic;
signal \N__77557\ : std_logic;
signal \N__77554\ : std_logic;
signal \N__77551\ : std_logic;
signal \N__77546\ : std_logic;
signal \N__77543\ : std_logic;
signal \N__77538\ : std_logic;
signal \N__77535\ : std_logic;
signal \N__77532\ : std_logic;
signal \N__77529\ : std_logic;
signal \N__77526\ : std_logic;
signal \N__77517\ : std_logic;
signal \N__77514\ : std_logic;
signal \N__77511\ : std_logic;
signal \N__77508\ : std_logic;
signal \N__77505\ : std_logic;
signal \N__77502\ : std_logic;
signal \N__77501\ : std_logic;
signal \N__77498\ : std_logic;
signal \N__77495\ : std_logic;
signal \N__77490\ : std_logic;
signal \N__77489\ : std_logic;
signal \N__77486\ : std_logic;
signal \N__77483\ : std_logic;
signal \N__77480\ : std_logic;
signal \N__77477\ : std_logic;
signal \N__77474\ : std_logic;
signal \N__77471\ : std_logic;
signal \N__77466\ : std_logic;
signal \N__77463\ : std_logic;
signal \N__77460\ : std_logic;
signal \N__77457\ : std_logic;
signal \N__77454\ : std_logic;
signal \N__77453\ : std_logic;
signal \N__77450\ : std_logic;
signal \N__77447\ : std_logic;
signal \N__77446\ : std_logic;
signal \N__77441\ : std_logic;
signal \N__77440\ : std_logic;
signal \N__77437\ : std_logic;
signal \N__77434\ : std_logic;
signal \N__77431\ : std_logic;
signal \N__77428\ : std_logic;
signal \N__77421\ : std_logic;
signal \N__77418\ : std_logic;
signal \N__77417\ : std_logic;
signal \N__77414\ : std_logic;
signal \N__77411\ : std_logic;
signal \N__77406\ : std_logic;
signal \N__77405\ : std_logic;
signal \N__77402\ : std_logic;
signal \N__77399\ : std_logic;
signal \N__77394\ : std_logic;
signal \N__77393\ : std_logic;
signal \N__77392\ : std_logic;
signal \N__77391\ : std_logic;
signal \N__77388\ : std_logic;
signal \N__77383\ : std_logic;
signal \N__77380\ : std_logic;
signal \N__77377\ : std_logic;
signal \N__77376\ : std_logic;
signal \N__77373\ : std_logic;
signal \N__77368\ : std_logic;
signal \N__77365\ : std_logic;
signal \N__77362\ : std_logic;
signal \N__77355\ : std_logic;
signal \N__77352\ : std_logic;
signal \N__77351\ : std_logic;
signal \N__77348\ : std_logic;
signal \N__77345\ : std_logic;
signal \N__77342\ : std_logic;
signal \N__77341\ : std_logic;
signal \N__77336\ : std_logic;
signal \N__77333\ : std_logic;
signal \N__77332\ : std_logic;
signal \N__77329\ : std_logic;
signal \N__77326\ : std_logic;
signal \N__77323\ : std_logic;
signal \N__77318\ : std_logic;
signal \N__77315\ : std_logic;
signal \N__77312\ : std_logic;
signal \N__77307\ : std_logic;
signal \N__77304\ : std_logic;
signal \N__77301\ : std_logic;
signal \N__77298\ : std_logic;
signal \N__77295\ : std_logic;
signal \N__77292\ : std_logic;
signal \N__77291\ : std_logic;
signal \N__77288\ : std_logic;
signal \N__77287\ : std_logic;
signal \N__77284\ : std_logic;
signal \N__77281\ : std_logic;
signal \N__77280\ : std_logic;
signal \N__77277\ : std_logic;
signal \N__77274\ : std_logic;
signal \N__77273\ : std_logic;
signal \N__77270\ : std_logic;
signal \N__77267\ : std_logic;
signal \N__77266\ : std_logic;
signal \N__77261\ : std_logic;
signal \N__77258\ : std_logic;
signal \N__77255\ : std_logic;
signal \N__77252\ : std_logic;
signal \N__77249\ : std_logic;
signal \N__77246\ : std_logic;
signal \N__77243\ : std_logic;
signal \N__77238\ : std_logic;
signal \N__77229\ : std_logic;
signal \N__77226\ : std_logic;
signal \N__77223\ : std_logic;
signal \N__77220\ : std_logic;
signal \N__77217\ : std_logic;
signal \N__77216\ : std_logic;
signal \N__77213\ : std_logic;
signal \N__77210\ : std_logic;
signal \N__77209\ : std_logic;
signal \N__77204\ : std_logic;
signal \N__77201\ : std_logic;
signal \N__77198\ : std_logic;
signal \N__77195\ : std_logic;
signal \N__77190\ : std_logic;
signal \N__77189\ : std_logic;
signal \N__77188\ : std_logic;
signal \N__77187\ : std_logic;
signal \N__77184\ : std_logic;
signal \N__77181\ : std_logic;
signal \N__77180\ : std_logic;
signal \N__77177\ : std_logic;
signal \N__77174\ : std_logic;
signal \N__77171\ : std_logic;
signal \N__77168\ : std_logic;
signal \N__77165\ : std_logic;
signal \N__77162\ : std_logic;
signal \N__77151\ : std_logic;
signal \N__77150\ : std_logic;
signal \N__77147\ : std_logic;
signal \N__77144\ : std_logic;
signal \N__77141\ : std_logic;
signal \N__77138\ : std_logic;
signal \N__77133\ : std_logic;
signal \N__77132\ : std_logic;
signal \N__77131\ : std_logic;
signal \N__77130\ : std_logic;
signal \N__77129\ : std_logic;
signal \N__77128\ : std_logic;
signal \N__77125\ : std_logic;
signal \N__77124\ : std_logic;
signal \N__77123\ : std_logic;
signal \N__77122\ : std_logic;
signal \N__77121\ : std_logic;
signal \N__77118\ : std_logic;
signal \N__77115\ : std_logic;
signal \N__77112\ : std_logic;
signal \N__77111\ : std_logic;
signal \N__77110\ : std_logic;
signal \N__77107\ : std_logic;
signal \N__77106\ : std_logic;
signal \N__77103\ : std_logic;
signal \N__77102\ : std_logic;
signal \N__77101\ : std_logic;
signal \N__77100\ : std_logic;
signal \N__77099\ : std_logic;
signal \N__77098\ : std_logic;
signal \N__77093\ : std_logic;
signal \N__77092\ : std_logic;
signal \N__77091\ : std_logic;
signal \N__77090\ : std_logic;
signal \N__77087\ : std_logic;
signal \N__77084\ : std_logic;
signal \N__77081\ : std_logic;
signal \N__77078\ : std_logic;
signal \N__77075\ : std_logic;
signal \N__77072\ : std_logic;
signal \N__77069\ : std_logic;
signal \N__77066\ : std_logic;
signal \N__77065\ : std_logic;
signal \N__77062\ : std_logic;
signal \N__77059\ : std_logic;
signal \N__77058\ : std_logic;
signal \N__77055\ : std_logic;
signal \N__77052\ : std_logic;
signal \N__77049\ : std_logic;
signal \N__77046\ : std_logic;
signal \N__77045\ : std_logic;
signal \N__77044\ : std_logic;
signal \N__77041\ : std_logic;
signal \N__77038\ : std_logic;
signal \N__77035\ : std_logic;
signal \N__77028\ : std_logic;
signal \N__77023\ : std_logic;
signal \N__77020\ : std_logic;
signal \N__77017\ : std_logic;
signal \N__77012\ : std_logic;
signal \N__77009\ : std_logic;
signal \N__77006\ : std_logic;
signal \N__77003\ : std_logic;
signal \N__76998\ : std_logic;
signal \N__76997\ : std_logic;
signal \N__76994\ : std_logic;
signal \N__76985\ : std_logic;
signal \N__76982\ : std_logic;
signal \N__76979\ : std_logic;
signal \N__76974\ : std_logic;
signal \N__76963\ : std_logic;
signal \N__76958\ : std_logic;
signal \N__76955\ : std_logic;
signal \N__76954\ : std_logic;
signal \N__76949\ : std_logic;
signal \N__76946\ : std_logic;
signal \N__76945\ : std_logic;
signal \N__76944\ : std_logic;
signal \N__76941\ : std_logic;
signal \N__76936\ : std_logic;
signal \N__76933\ : std_logic;
signal \N__76926\ : std_logic;
signal \N__76923\ : std_logic;
signal \N__76920\ : std_logic;
signal \N__76917\ : std_logic;
signal \N__76916\ : std_logic;
signal \N__76913\ : std_logic;
signal \N__76912\ : std_logic;
signal \N__76909\ : std_logic;
signal \N__76906\ : std_logic;
signal \N__76903\ : std_logic;
signal \N__76900\ : std_logic;
signal \N__76895\ : std_logic;
signal \N__76892\ : std_logic;
signal \N__76887\ : std_logic;
signal \N__76884\ : std_logic;
signal \N__76883\ : std_logic;
signal \N__76880\ : std_logic;
signal \N__76877\ : std_logic;
signal \N__76874\ : std_logic;
signal \N__76865\ : std_logic;
signal \N__76860\ : std_logic;
signal \N__76855\ : std_logic;
signal \N__76852\ : std_logic;
signal \N__76845\ : std_logic;
signal \N__76842\ : std_logic;
signal \N__76833\ : std_logic;
signal \N__76832\ : std_logic;
signal \N__76829\ : std_logic;
signal \N__76828\ : std_logic;
signal \N__76825\ : std_logic;
signal \N__76822\ : std_logic;
signal \N__76819\ : std_logic;
signal \N__76816\ : std_logic;
signal \N__76815\ : std_logic;
signal \N__76810\ : std_logic;
signal \N__76807\ : std_logic;
signal \N__76804\ : std_logic;
signal \N__76801\ : std_logic;
signal \N__76798\ : std_logic;
signal \N__76797\ : std_logic;
signal \N__76794\ : std_logic;
signal \N__76791\ : std_logic;
signal \N__76788\ : std_logic;
signal \N__76785\ : std_logic;
signal \N__76776\ : std_logic;
signal \N__76773\ : std_logic;
signal \N__76770\ : std_logic;
signal \N__76767\ : std_logic;
signal \N__76764\ : std_logic;
signal \N__76761\ : std_logic;
signal \N__76758\ : std_logic;
signal \N__76755\ : std_logic;
signal \N__76752\ : std_logic;
signal \N__76749\ : std_logic;
signal \N__76746\ : std_logic;
signal \N__76743\ : std_logic;
signal \N__76742\ : std_logic;
signal \N__76741\ : std_logic;
signal \N__76738\ : std_logic;
signal \N__76735\ : std_logic;
signal \N__76732\ : std_logic;
signal \N__76727\ : std_logic;
signal \N__76726\ : std_logic;
signal \N__76723\ : std_logic;
signal \N__76720\ : std_logic;
signal \N__76717\ : std_logic;
signal \N__76710\ : std_logic;
signal \N__76707\ : std_logic;
signal \N__76704\ : std_logic;
signal \N__76701\ : std_logic;
signal \N__76698\ : std_logic;
signal \N__76695\ : std_logic;
signal \N__76694\ : std_logic;
signal \N__76693\ : std_logic;
signal \N__76688\ : std_logic;
signal \N__76687\ : std_logic;
signal \N__76684\ : std_logic;
signal \N__76683\ : std_logic;
signal \N__76682\ : std_logic;
signal \N__76679\ : std_logic;
signal \N__76676\ : std_logic;
signal \N__76675\ : std_logic;
signal \N__76674\ : std_logic;
signal \N__76671\ : std_logic;
signal \N__76668\ : std_logic;
signal \N__76665\ : std_logic;
signal \N__76660\ : std_logic;
signal \N__76657\ : std_logic;
signal \N__76656\ : std_logic;
signal \N__76655\ : std_logic;
signal \N__76654\ : std_logic;
signal \N__76653\ : std_logic;
signal \N__76652\ : std_logic;
signal \N__76649\ : std_logic;
signal \N__76644\ : std_logic;
signal \N__76641\ : std_logic;
signal \N__76636\ : std_logic;
signal \N__76631\ : std_logic;
signal \N__76630\ : std_logic;
signal \N__76629\ : std_logic;
signal \N__76626\ : std_logic;
signal \N__76625\ : std_logic;
signal \N__76624\ : std_logic;
signal \N__76623\ : std_logic;
signal \N__76622\ : std_logic;
signal \N__76617\ : std_logic;
signal \N__76614\ : std_logic;
signal \N__76613\ : std_logic;
signal \N__76612\ : std_logic;
signal \N__76611\ : std_logic;
signal \N__76610\ : std_logic;
signal \N__76607\ : std_logic;
signal \N__76600\ : std_logic;
signal \N__76599\ : std_logic;
signal \N__76596\ : std_logic;
signal \N__76595\ : std_logic;
signal \N__76592\ : std_logic;
signal \N__76589\ : std_logic;
signal \N__76586\ : std_logic;
signal \N__76583\ : std_logic;
signal \N__76582\ : std_logic;
signal \N__76579\ : std_logic;
signal \N__76576\ : std_logic;
signal \N__76573\ : std_logic;
signal \N__76570\ : std_logic;
signal \N__76567\ : std_logic;
signal \N__76564\ : std_logic;
signal \N__76559\ : std_logic;
signal \N__76554\ : std_logic;
signal \N__76551\ : std_logic;
signal \N__76550\ : std_logic;
signal \N__76549\ : std_logic;
signal \N__76548\ : std_logic;
signal \N__76545\ : std_logic;
signal \N__76542\ : std_logic;
signal \N__76539\ : std_logic;
signal \N__76536\ : std_logic;
signal \N__76531\ : std_logic;
signal \N__76530\ : std_logic;
signal \N__76529\ : std_logic;
signal \N__76526\ : std_logic;
signal \N__76525\ : std_logic;
signal \N__76520\ : std_logic;
signal \N__76513\ : std_logic;
signal \N__76510\ : std_logic;
signal \N__76505\ : std_logic;
signal \N__76502\ : std_logic;
signal \N__76499\ : std_logic;
signal \N__76496\ : std_logic;
signal \N__76493\ : std_logic;
signal \N__76484\ : std_logic;
signal \N__76481\ : std_logic;
signal \N__76478\ : std_logic;
signal \N__76475\ : std_logic;
signal \N__76472\ : std_logic;
signal \N__76469\ : std_logic;
signal \N__76464\ : std_logic;
signal \N__76459\ : std_logic;
signal \N__76456\ : std_logic;
signal \N__76449\ : std_logic;
signal \N__76446\ : std_logic;
signal \N__76443\ : std_logic;
signal \N__76434\ : std_logic;
signal \N__76429\ : std_logic;
signal \N__76426\ : std_logic;
signal \N__76423\ : std_logic;
signal \N__76420\ : std_logic;
signal \N__76417\ : std_logic;
signal \N__76414\ : std_logic;
signal \N__76411\ : std_logic;
signal \N__76398\ : std_logic;
signal \N__76395\ : std_logic;
signal \N__76394\ : std_logic;
signal \N__76393\ : std_logic;
signal \N__76390\ : std_logic;
signal \N__76389\ : std_logic;
signal \N__76386\ : std_logic;
signal \N__76385\ : std_logic;
signal \N__76384\ : std_logic;
signal \N__76383\ : std_logic;
signal \N__76382\ : std_logic;
signal \N__76379\ : std_logic;
signal \N__76378\ : std_logic;
signal \N__76375\ : std_logic;
signal \N__76372\ : std_logic;
signal \N__76369\ : std_logic;
signal \N__76366\ : std_logic;
signal \N__76365\ : std_logic;
signal \N__76362\ : std_logic;
signal \N__76359\ : std_logic;
signal \N__76356\ : std_logic;
signal \N__76355\ : std_logic;
signal \N__76354\ : std_logic;
signal \N__76351\ : std_logic;
signal \N__76348\ : std_logic;
signal \N__76343\ : std_logic;
signal \N__76338\ : std_logic;
signal \N__76335\ : std_logic;
signal \N__76332\ : std_logic;
signal \N__76329\ : std_logic;
signal \N__76326\ : std_logic;
signal \N__76325\ : std_logic;
signal \N__76324\ : std_logic;
signal \N__76321\ : std_logic;
signal \N__76318\ : std_logic;
signal \N__76317\ : std_logic;
signal \N__76316\ : std_logic;
signal \N__76315\ : std_logic;
signal \N__76310\ : std_logic;
signal \N__76305\ : std_logic;
signal \N__76302\ : std_logic;
signal \N__76295\ : std_logic;
signal \N__76294\ : std_logic;
signal \N__76293\ : std_logic;
signal \N__76290\ : std_logic;
signal \N__76289\ : std_logic;
signal \N__76286\ : std_logic;
signal \N__76285\ : std_logic;
signal \N__76282\ : std_logic;
signal \N__76279\ : std_logic;
signal \N__76276\ : std_logic;
signal \N__76275\ : std_logic;
signal \N__76274\ : std_logic;
signal \N__76271\ : std_logic;
signal \N__76268\ : std_logic;
signal \N__76265\ : std_logic;
signal \N__76260\ : std_logic;
signal \N__76257\ : std_logic;
signal \N__76254\ : std_logic;
signal \N__76251\ : std_logic;
signal \N__76248\ : std_logic;
signal \N__76245\ : std_logic;
signal \N__76242\ : std_logic;
signal \N__76239\ : std_logic;
signal \N__76232\ : std_logic;
signal \N__76229\ : std_logic;
signal \N__76228\ : std_logic;
signal \N__76227\ : std_logic;
signal \N__76224\ : std_logic;
signal \N__76221\ : std_logic;
signal \N__76218\ : std_logic;
signal \N__76215\ : std_logic;
signal \N__76212\ : std_logic;
signal \N__76209\ : std_logic;
signal \N__76206\ : std_logic;
signal \N__76199\ : std_logic;
signal \N__76194\ : std_logic;
signal \N__76191\ : std_logic;
signal \N__76188\ : std_logic;
signal \N__76183\ : std_logic;
signal \N__76180\ : std_logic;
signal \N__76175\ : std_logic;
signal \N__76172\ : std_logic;
signal \N__76167\ : std_logic;
signal \N__76164\ : std_logic;
signal \N__76161\ : std_logic;
signal \N__76158\ : std_logic;
signal \N__76155\ : std_logic;
signal \N__76154\ : std_logic;
signal \N__76153\ : std_logic;
signal \N__76152\ : std_logic;
signal \N__76151\ : std_logic;
signal \N__76150\ : std_logic;
signal \N__76149\ : std_logic;
signal \N__76148\ : std_logic;
signal \N__76135\ : std_logic;
signal \N__76130\ : std_logic;
signal \N__76125\ : std_logic;
signal \N__76122\ : std_logic;
signal \N__76117\ : std_logic;
signal \N__76112\ : std_logic;
signal \N__76107\ : std_logic;
signal \N__76104\ : std_logic;
signal \N__76099\ : std_logic;
signal \N__76086\ : std_logic;
signal \N__76083\ : std_logic;
signal \N__76082\ : std_logic;
signal \N__76079\ : std_logic;
signal \N__76076\ : std_logic;
signal \N__76071\ : std_logic;
signal \N__76070\ : std_logic;
signal \N__76067\ : std_logic;
signal \N__76064\ : std_logic;
signal \N__76061\ : std_logic;
signal \N__76058\ : std_logic;
signal \N__76053\ : std_logic;
signal \N__76052\ : std_logic;
signal \N__76049\ : std_logic;
signal \N__76048\ : std_logic;
signal \N__76047\ : std_logic;
signal \N__76044\ : std_logic;
signal \N__76041\ : std_logic;
signal \N__76038\ : std_logic;
signal \N__76037\ : std_logic;
signal \N__76036\ : std_logic;
signal \N__76033\ : std_logic;
signal \N__76030\ : std_logic;
signal \N__76027\ : std_logic;
signal \N__76022\ : std_logic;
signal \N__76019\ : std_logic;
signal \N__76016\ : std_logic;
signal \N__76013\ : std_logic;
signal \N__76008\ : std_logic;
signal \N__76005\ : std_logic;
signal \N__75996\ : std_logic;
signal \N__75993\ : std_logic;
signal \N__75990\ : std_logic;
signal \N__75989\ : std_logic;
signal \N__75986\ : std_logic;
signal \N__75983\ : std_logic;
signal \N__75980\ : std_logic;
signal \N__75977\ : std_logic;
signal \N__75974\ : std_logic;
signal \N__75969\ : std_logic;
signal \N__75966\ : std_logic;
signal \N__75963\ : std_logic;
signal \N__75962\ : std_logic;
signal \N__75959\ : std_logic;
signal \N__75956\ : std_logic;
signal \N__75951\ : std_logic;
signal \N__75948\ : std_logic;
signal \N__75947\ : std_logic;
signal \N__75946\ : std_logic;
signal \N__75943\ : std_logic;
signal \N__75940\ : std_logic;
signal \N__75939\ : std_logic;
signal \N__75938\ : std_logic;
signal \N__75935\ : std_logic;
signal \N__75932\ : std_logic;
signal \N__75929\ : std_logic;
signal \N__75926\ : std_logic;
signal \N__75923\ : std_logic;
signal \N__75920\ : std_logic;
signal \N__75913\ : std_logic;
signal \N__75910\ : std_logic;
signal \N__75909\ : std_logic;
signal \N__75906\ : std_logic;
signal \N__75903\ : std_logic;
signal \N__75900\ : std_logic;
signal \N__75897\ : std_logic;
signal \N__75894\ : std_logic;
signal \N__75891\ : std_logic;
signal \N__75888\ : std_logic;
signal \N__75883\ : std_logic;
signal \N__75880\ : std_logic;
signal \N__75873\ : std_logic;
signal \N__75870\ : std_logic;
signal \N__75867\ : std_logic;
signal \N__75864\ : std_logic;
signal \N__75861\ : std_logic;
signal \N__75858\ : std_logic;
signal \N__75857\ : std_logic;
signal \N__75854\ : std_logic;
signal \N__75851\ : std_logic;
signal \N__75848\ : std_logic;
signal \N__75847\ : std_logic;
signal \N__75844\ : std_logic;
signal \N__75841\ : std_logic;
signal \N__75838\ : std_logic;
signal \N__75831\ : std_logic;
signal \N__75830\ : std_logic;
signal \N__75827\ : std_logic;
signal \N__75824\ : std_logic;
signal \N__75823\ : std_logic;
signal \N__75820\ : std_logic;
signal \N__75815\ : std_logic;
signal \N__75810\ : std_logic;
signal \N__75807\ : std_logic;
signal \N__75804\ : std_logic;
signal \N__75801\ : std_logic;
signal \N__75798\ : std_logic;
signal \N__75795\ : std_logic;
signal \N__75792\ : std_logic;
signal \N__75789\ : std_logic;
signal \N__75786\ : std_logic;
signal \N__75785\ : std_logic;
signal \N__75784\ : std_logic;
signal \N__75779\ : std_logic;
signal \N__75778\ : std_logic;
signal \N__75775\ : std_logic;
signal \N__75772\ : std_logic;
signal \N__75769\ : std_logic;
signal \N__75766\ : std_logic;
signal \N__75765\ : std_logic;
signal \N__75762\ : std_logic;
signal \N__75757\ : std_logic;
signal \N__75754\ : std_logic;
signal \N__75751\ : std_logic;
signal \N__75748\ : std_logic;
signal \N__75745\ : std_logic;
signal \N__75742\ : std_logic;
signal \N__75739\ : std_logic;
signal \N__75732\ : std_logic;
signal \N__75731\ : std_logic;
signal \N__75730\ : std_logic;
signal \N__75729\ : std_logic;
signal \N__75726\ : std_logic;
signal \N__75719\ : std_logic;
signal \N__75716\ : std_logic;
signal \N__75713\ : std_logic;
signal \N__75708\ : std_logic;
signal \N__75705\ : std_logic;
signal \N__75702\ : std_logic;
signal \N__75701\ : std_logic;
signal \N__75700\ : std_logic;
signal \N__75697\ : std_logic;
signal \N__75694\ : std_logic;
signal \N__75691\ : std_logic;
signal \N__75688\ : std_logic;
signal \N__75685\ : std_logic;
signal \N__75682\ : std_logic;
signal \N__75679\ : std_logic;
signal \N__75678\ : std_logic;
signal \N__75675\ : std_logic;
signal \N__75672\ : std_logic;
signal \N__75669\ : std_logic;
signal \N__75666\ : std_logic;
signal \N__75663\ : std_logic;
signal \N__75660\ : std_logic;
signal \N__75657\ : std_logic;
signal \N__75654\ : std_logic;
signal \N__75649\ : std_logic;
signal \N__75646\ : std_logic;
signal \N__75641\ : std_logic;
signal \N__75636\ : std_logic;
signal \N__75633\ : std_logic;
signal \N__75630\ : std_logic;
signal \N__75627\ : std_logic;
signal \N__75624\ : std_logic;
signal \N__75621\ : std_logic;
signal \N__75620\ : std_logic;
signal \N__75615\ : std_logic;
signal \N__75614\ : std_logic;
signal \N__75613\ : std_logic;
signal \N__75612\ : std_logic;
signal \N__75611\ : std_logic;
signal \N__75608\ : std_logic;
signal \N__75605\ : std_logic;
signal \N__75600\ : std_logic;
signal \N__75597\ : std_logic;
signal \N__75590\ : std_logic;
signal \N__75587\ : std_logic;
signal \N__75584\ : std_logic;
signal \N__75579\ : std_logic;
signal \N__75576\ : std_logic;
signal \N__75573\ : std_logic;
signal \N__75570\ : std_logic;
signal \N__75567\ : std_logic;
signal \N__75566\ : std_logic;
signal \N__75563\ : std_logic;
signal \N__75562\ : std_logic;
signal \N__75559\ : std_logic;
signal \N__75558\ : std_logic;
signal \N__75555\ : std_logic;
signal \N__75554\ : std_logic;
signal \N__75553\ : std_logic;
signal \N__75550\ : std_logic;
signal \N__75549\ : std_logic;
signal \N__75548\ : std_logic;
signal \N__75545\ : std_logic;
signal \N__75542\ : std_logic;
signal \N__75539\ : std_logic;
signal \N__75536\ : std_logic;
signal \N__75533\ : std_logic;
signal \N__75528\ : std_logic;
signal \N__75525\ : std_logic;
signal \N__75522\ : std_logic;
signal \N__75507\ : std_logic;
signal \N__75506\ : std_logic;
signal \N__75501\ : std_logic;
signal \N__75500\ : std_logic;
signal \N__75499\ : std_logic;
signal \N__75498\ : std_logic;
signal \N__75495\ : std_logic;
signal \N__75494\ : std_logic;
signal \N__75493\ : std_logic;
signal \N__75492\ : std_logic;
signal \N__75489\ : std_logic;
signal \N__75484\ : std_logic;
signal \N__75481\ : std_logic;
signal \N__75476\ : std_logic;
signal \N__75473\ : std_logic;
signal \N__75470\ : std_logic;
signal \N__75467\ : std_logic;
signal \N__75464\ : std_logic;
signal \N__75461\ : std_logic;
signal \N__75458\ : std_logic;
signal \N__75455\ : std_logic;
signal \N__75452\ : std_logic;
signal \N__75449\ : std_logic;
signal \N__75442\ : std_logic;
signal \N__75439\ : std_logic;
signal \N__75436\ : std_logic;
signal \N__75433\ : std_logic;
signal \N__75426\ : std_logic;
signal \N__75423\ : std_logic;
signal \N__75422\ : std_logic;
signal \N__75421\ : std_logic;
signal \N__75420\ : std_logic;
signal \N__75417\ : std_logic;
signal \N__75416\ : std_logic;
signal \N__75415\ : std_logic;
signal \N__75408\ : std_logic;
signal \N__75407\ : std_logic;
signal \N__75406\ : std_logic;
signal \N__75403\ : std_logic;
signal \N__75400\ : std_logic;
signal \N__75399\ : std_logic;
signal \N__75398\ : std_logic;
signal \N__75397\ : std_logic;
signal \N__75394\ : std_logic;
signal \N__75393\ : std_logic;
signal \N__75390\ : std_logic;
signal \N__75385\ : std_logic;
signal \N__75380\ : std_logic;
signal \N__75375\ : std_logic;
signal \N__75374\ : std_logic;
signal \N__75373\ : std_logic;
signal \N__75370\ : std_logic;
signal \N__75367\ : std_logic;
signal \N__75364\ : std_logic;
signal \N__75359\ : std_logic;
signal \N__75356\ : std_logic;
signal \N__75353\ : std_logic;
signal \N__75350\ : std_logic;
signal \N__75347\ : std_logic;
signal \N__75344\ : std_logic;
signal \N__75341\ : std_logic;
signal \N__75338\ : std_logic;
signal \N__75337\ : std_logic;
signal \N__75334\ : std_logic;
signal \N__75331\ : std_logic;
signal \N__75328\ : std_logic;
signal \N__75327\ : std_logic;
signal \N__75326\ : std_logic;
signal \N__75321\ : std_logic;
signal \N__75318\ : std_logic;
signal \N__75313\ : std_logic;
signal \N__75310\ : std_logic;
signal \N__75307\ : std_logic;
signal \N__75302\ : std_logic;
signal \N__75301\ : std_logic;
signal \N__75298\ : std_logic;
signal \N__75295\ : std_logic;
signal \N__75290\ : std_logic;
signal \N__75287\ : std_logic;
signal \N__75280\ : std_logic;
signal \N__75277\ : std_logic;
signal \N__75274\ : std_logic;
signal \N__75261\ : std_logic;
signal \N__75258\ : std_logic;
signal \N__75257\ : std_logic;
signal \N__75256\ : std_logic;
signal \N__75255\ : std_logic;
signal \N__75254\ : std_logic;
signal \N__75253\ : std_logic;
signal \N__75252\ : std_logic;
signal \N__75251\ : std_logic;
signal \N__75250\ : std_logic;
signal \N__75249\ : std_logic;
signal \N__75248\ : std_logic;
signal \N__75245\ : std_logic;
signal \N__75244\ : std_logic;
signal \N__75243\ : std_logic;
signal \N__75242\ : std_logic;
signal \N__75239\ : std_logic;
signal \N__75236\ : std_logic;
signal \N__75233\ : std_logic;
signal \N__75230\ : std_logic;
signal \N__75229\ : std_logic;
signal \N__75228\ : std_logic;
signal \N__75225\ : std_logic;
signal \N__75224\ : std_logic;
signal \N__75219\ : std_logic;
signal \N__75216\ : std_logic;
signal \N__75211\ : std_logic;
signal \N__75208\ : std_logic;
signal \N__75205\ : std_logic;
signal \N__75202\ : std_logic;
signal \N__75199\ : std_logic;
signal \N__75196\ : std_logic;
signal \N__75195\ : std_logic;
signal \N__75190\ : std_logic;
signal \N__75187\ : std_logic;
signal \N__75186\ : std_logic;
signal \N__75185\ : std_logic;
signal \N__75182\ : std_logic;
signal \N__75179\ : std_logic;
signal \N__75178\ : std_logic;
signal \N__75177\ : std_logic;
signal \N__75174\ : std_logic;
signal \N__75171\ : std_logic;
signal \N__75166\ : std_logic;
signal \N__75163\ : std_logic;
signal \N__75160\ : std_logic;
signal \N__75153\ : std_logic;
signal \N__75150\ : std_logic;
signal \N__75147\ : std_logic;
signal \N__75142\ : std_logic;
signal \N__75139\ : std_logic;
signal \N__75138\ : std_logic;
signal \N__75137\ : std_logic;
signal \N__75134\ : std_logic;
signal \N__75131\ : std_logic;
signal \N__75128\ : std_logic;
signal \N__75125\ : std_logic;
signal \N__75122\ : std_logic;
signal \N__75117\ : std_logic;
signal \N__75114\ : std_logic;
signal \N__75113\ : std_logic;
signal \N__75112\ : std_logic;
signal \N__75111\ : std_logic;
signal \N__75110\ : std_logic;
signal \N__75103\ : std_logic;
signal \N__75098\ : std_logic;
signal \N__75093\ : std_logic;
signal \N__75088\ : std_logic;
signal \N__75085\ : std_logic;
signal \N__75080\ : std_logic;
signal \N__75077\ : std_logic;
signal \N__75074\ : std_logic;
signal \N__75071\ : std_logic;
signal \N__75068\ : std_logic;
signal \N__75065\ : std_logic;
signal \N__75062\ : std_logic;
signal \N__75057\ : std_logic;
signal \N__75054\ : std_logic;
signal \N__75051\ : std_logic;
signal \N__75048\ : std_logic;
signal \N__75047\ : std_logic;
signal \N__75046\ : std_logic;
signal \N__75041\ : std_logic;
signal \N__75034\ : std_logic;
signal \N__75029\ : std_logic;
signal \N__75028\ : std_logic;
signal \N__75027\ : std_logic;
signal \N__75022\ : std_logic;
signal \N__75019\ : std_logic;
signal \N__75012\ : std_logic;
signal \N__75007\ : std_logic;
signal \N__75002\ : std_logic;
signal \N__74999\ : std_logic;
signal \N__74996\ : std_logic;
signal \N__74993\ : std_logic;
signal \N__74990\ : std_logic;
signal \N__74987\ : std_logic;
signal \N__74984\ : std_logic;
signal \N__74977\ : std_logic;
signal \N__74964\ : std_logic;
signal \N__74963\ : std_logic;
signal \N__74962\ : std_logic;
signal \N__74961\ : std_logic;
signal \N__74958\ : std_logic;
signal \N__74955\ : std_logic;
signal \N__74952\ : std_logic;
signal \N__74949\ : std_logic;
signal \N__74946\ : std_logic;
signal \N__74943\ : std_logic;
signal \N__74940\ : std_logic;
signal \N__74937\ : std_logic;
signal \N__74934\ : std_logic;
signal \N__74933\ : std_logic;
signal \N__74930\ : std_logic;
signal \N__74927\ : std_logic;
signal \N__74922\ : std_logic;
signal \N__74919\ : std_logic;
signal \N__74914\ : std_logic;
signal \N__74911\ : std_logic;
signal \N__74904\ : std_logic;
signal \N__74903\ : std_logic;
signal \N__74900\ : std_logic;
signal \N__74897\ : std_logic;
signal \N__74894\ : std_logic;
signal \N__74893\ : std_logic;
signal \N__74890\ : std_logic;
signal \N__74887\ : std_logic;
signal \N__74884\ : std_logic;
signal \N__74881\ : std_logic;
signal \N__74874\ : std_logic;
signal \N__74871\ : std_logic;
signal \N__74870\ : std_logic;
signal \N__74867\ : std_logic;
signal \N__74866\ : std_logic;
signal \N__74863\ : std_logic;
signal \N__74860\ : std_logic;
signal \N__74857\ : std_logic;
signal \N__74854\ : std_logic;
signal \N__74851\ : std_logic;
signal \N__74848\ : std_logic;
signal \N__74841\ : std_logic;
signal \N__74838\ : std_logic;
signal \N__74837\ : std_logic;
signal \N__74834\ : std_logic;
signal \N__74831\ : std_logic;
signal \N__74828\ : std_logic;
signal \N__74825\ : std_logic;
signal \N__74822\ : std_logic;
signal \N__74817\ : std_logic;
signal \N__74816\ : std_logic;
signal \N__74815\ : std_logic;
signal \N__74812\ : std_logic;
signal \N__74811\ : std_logic;
signal \N__74808\ : std_logic;
signal \N__74805\ : std_logic;
signal \N__74802\ : std_logic;
signal \N__74799\ : std_logic;
signal \N__74794\ : std_logic;
signal \N__74789\ : std_logic;
signal \N__74786\ : std_logic;
signal \N__74783\ : std_logic;
signal \N__74778\ : std_logic;
signal \N__74775\ : std_logic;
signal \N__74774\ : std_logic;
signal \N__74773\ : std_logic;
signal \N__74772\ : std_logic;
signal \N__74769\ : std_logic;
signal \N__74768\ : std_logic;
signal \N__74765\ : std_logic;
signal \N__74760\ : std_logic;
signal \N__74757\ : std_logic;
signal \N__74752\ : std_logic;
signal \N__74745\ : std_logic;
signal \N__74742\ : std_logic;
signal \N__74739\ : std_logic;
signal \N__74736\ : std_logic;
signal \N__74733\ : std_logic;
signal \N__74730\ : std_logic;
signal \N__74727\ : std_logic;
signal \N__74724\ : std_logic;
signal \N__74721\ : std_logic;
signal \N__74718\ : std_logic;
signal \N__74715\ : std_logic;
signal \N__74714\ : std_logic;
signal \N__74713\ : std_logic;
signal \N__74712\ : std_logic;
signal \N__74709\ : std_logic;
signal \N__74704\ : std_logic;
signal \N__74701\ : std_logic;
signal \N__74698\ : std_logic;
signal \N__74695\ : std_logic;
signal \N__74692\ : std_logic;
signal \N__74689\ : std_logic;
signal \N__74686\ : std_logic;
signal \N__74679\ : std_logic;
signal \N__74678\ : std_logic;
signal \N__74675\ : std_logic;
signal \N__74674\ : std_logic;
signal \N__74673\ : std_logic;
signal \N__74670\ : std_logic;
signal \N__74667\ : std_logic;
signal \N__74666\ : std_logic;
signal \N__74663\ : std_logic;
signal \N__74660\ : std_logic;
signal \N__74659\ : std_logic;
signal \N__74658\ : std_logic;
signal \N__74655\ : std_logic;
signal \N__74652\ : std_logic;
signal \N__74647\ : std_logic;
signal \N__74644\ : std_logic;
signal \N__74643\ : std_logic;
signal \N__74642\ : std_logic;
signal \N__74637\ : std_logic;
signal \N__74636\ : std_logic;
signal \N__74633\ : std_logic;
signal \N__74632\ : std_logic;
signal \N__74631\ : std_logic;
signal \N__74626\ : std_logic;
signal \N__74625\ : std_logic;
signal \N__74622\ : std_logic;
signal \N__74619\ : std_logic;
signal \N__74616\ : std_logic;
signal \N__74613\ : std_logic;
signal \N__74610\ : std_logic;
signal \N__74607\ : std_logic;
signal \N__74604\ : std_logic;
signal \N__74601\ : std_logic;
signal \N__74598\ : std_logic;
signal \N__74595\ : std_logic;
signal \N__74592\ : std_logic;
signal \N__74589\ : std_logic;
signal \N__74586\ : std_logic;
signal \N__74581\ : std_logic;
signal \N__74578\ : std_logic;
signal \N__74573\ : std_logic;
signal \N__74570\ : std_logic;
signal \N__74563\ : std_logic;
signal \N__74562\ : std_logic;
signal \N__74559\ : std_logic;
signal \N__74556\ : std_logic;
signal \N__74553\ : std_logic;
signal \N__74548\ : std_logic;
signal \N__74545\ : std_logic;
signal \N__74542\ : std_logic;
signal \N__74529\ : std_logic;
signal \N__74526\ : std_logic;
signal \N__74525\ : std_logic;
signal \N__74524\ : std_logic;
signal \N__74521\ : std_logic;
signal \N__74520\ : std_logic;
signal \N__74517\ : std_logic;
signal \N__74514\ : std_logic;
signal \N__74511\ : std_logic;
signal \N__74508\ : std_logic;
signal \N__74507\ : std_logic;
signal \N__74504\ : std_logic;
signal \N__74501\ : std_logic;
signal \N__74500\ : std_logic;
signal \N__74499\ : std_logic;
signal \N__74498\ : std_logic;
signal \N__74493\ : std_logic;
signal \N__74490\ : std_logic;
signal \N__74487\ : std_logic;
signal \N__74484\ : std_logic;
signal \N__74481\ : std_logic;
signal \N__74480\ : std_logic;
signal \N__74477\ : std_logic;
signal \N__74474\ : std_logic;
signal \N__74471\ : std_logic;
signal \N__74470\ : std_logic;
signal \N__74469\ : std_logic;
signal \N__74466\ : std_logic;
signal \N__74459\ : std_logic;
signal \N__74456\ : std_logic;
signal \N__74453\ : std_logic;
signal \N__74448\ : std_logic;
signal \N__74447\ : std_logic;
signal \N__74442\ : std_logic;
signal \N__74441\ : std_logic;
signal \N__74436\ : std_logic;
signal \N__74429\ : std_logic;
signal \N__74426\ : std_logic;
signal \N__74423\ : std_logic;
signal \N__74420\ : std_logic;
signal \N__74417\ : std_logic;
signal \N__74414\ : std_logic;
signal \N__74407\ : std_logic;
signal \N__74406\ : std_logic;
signal \N__74403\ : std_logic;
signal \N__74398\ : std_logic;
signal \N__74395\ : std_logic;
signal \N__74388\ : std_logic;
signal \N__74387\ : std_logic;
signal \N__74386\ : std_logic;
signal \N__74383\ : std_logic;
signal \N__74382\ : std_logic;
signal \N__74381\ : std_logic;
signal \N__74378\ : std_logic;
signal \N__74375\ : std_logic;
signal \N__74372\ : std_logic;
signal \N__74369\ : std_logic;
signal \N__74366\ : std_logic;
signal \N__74365\ : std_logic;
signal \N__74362\ : std_logic;
signal \N__74359\ : std_logic;
signal \N__74358\ : std_logic;
signal \N__74355\ : std_logic;
signal \N__74352\ : std_logic;
signal \N__74349\ : std_logic;
signal \N__74348\ : std_logic;
signal \N__74345\ : std_logic;
signal \N__74344\ : std_logic;
signal \N__74341\ : std_logic;
signal \N__74338\ : std_logic;
signal \N__74335\ : std_logic;
signal \N__74332\ : std_logic;
signal \N__74329\ : std_logic;
signal \N__74326\ : std_logic;
signal \N__74323\ : std_logic;
signal \N__74320\ : std_logic;
signal \N__74317\ : std_logic;
signal \N__74312\ : std_logic;
signal \N__74309\ : std_logic;
signal \N__74306\ : std_logic;
signal \N__74303\ : std_logic;
signal \N__74302\ : std_logic;
signal \N__74297\ : std_logic;
signal \N__74292\ : std_logic;
signal \N__74289\ : std_logic;
signal \N__74288\ : std_logic;
signal \N__74285\ : std_logic;
signal \N__74280\ : std_logic;
signal \N__74279\ : std_logic;
signal \N__74276\ : std_logic;
signal \N__74273\ : std_logic;
signal \N__74270\ : std_logic;
signal \N__74267\ : std_logic;
signal \N__74264\ : std_logic;
signal \N__74259\ : std_logic;
signal \N__74256\ : std_logic;
signal \N__74247\ : std_logic;
signal \N__74242\ : std_logic;
signal \N__74239\ : std_logic;
signal \N__74238\ : std_logic;
signal \N__74235\ : std_logic;
signal \N__74230\ : std_logic;
signal \N__74227\ : std_logic;
signal \N__74220\ : std_logic;
signal \N__74217\ : std_logic;
signal \N__74216\ : std_logic;
signal \N__74213\ : std_logic;
signal \N__74210\ : std_logic;
signal \N__74209\ : std_logic;
signal \N__74208\ : std_logic;
signal \N__74207\ : std_logic;
signal \N__74206\ : std_logic;
signal \N__74205\ : std_logic;
signal \N__74204\ : std_logic;
signal \N__74203\ : std_logic;
signal \N__74202\ : std_logic;
signal \N__74197\ : std_logic;
signal \N__74194\ : std_logic;
signal \N__74189\ : std_logic;
signal \N__74188\ : std_logic;
signal \N__74187\ : std_logic;
signal \N__74184\ : std_logic;
signal \N__74181\ : std_logic;
signal \N__74180\ : std_logic;
signal \N__74179\ : std_logic;
signal \N__74178\ : std_logic;
signal \N__74171\ : std_logic;
signal \N__74166\ : std_logic;
signal \N__74163\ : std_logic;
signal \N__74158\ : std_logic;
signal \N__74157\ : std_logic;
signal \N__74156\ : std_logic;
signal \N__74151\ : std_logic;
signal \N__74150\ : std_logic;
signal \N__74147\ : std_logic;
signal \N__74146\ : std_logic;
signal \N__74145\ : std_logic;
signal \N__74142\ : std_logic;
signal \N__74139\ : std_logic;
signal \N__74136\ : std_logic;
signal \N__74135\ : std_logic;
signal \N__74132\ : std_logic;
signal \N__74127\ : std_logic;
signal \N__74124\ : std_logic;
signal \N__74121\ : std_logic;
signal \N__74118\ : std_logic;
signal \N__74117\ : std_logic;
signal \N__74116\ : std_logic;
signal \N__74115\ : std_logic;
signal \N__74112\ : std_logic;
signal \N__74111\ : std_logic;
signal \N__74108\ : std_logic;
signal \N__74105\ : std_logic;
signal \N__74104\ : std_logic;
signal \N__74101\ : std_logic;
signal \N__74098\ : std_logic;
signal \N__74095\ : std_logic;
signal \N__74092\ : std_logic;
signal \N__74089\ : std_logic;
signal \N__74086\ : std_logic;
signal \N__74081\ : std_logic;
signal \N__74076\ : std_logic;
signal \N__74073\ : std_logic;
signal \N__74070\ : std_logic;
signal \N__74069\ : std_logic;
signal \N__74068\ : std_logic;
signal \N__74067\ : std_logic;
signal \N__74066\ : std_logic;
signal \N__74063\ : std_logic;
signal \N__74060\ : std_logic;
signal \N__74057\ : std_logic;
signal \N__74052\ : std_logic;
signal \N__74051\ : std_logic;
signal \N__74048\ : std_logic;
signal \N__74045\ : std_logic;
signal \N__74040\ : std_logic;
signal \N__74035\ : std_logic;
signal \N__74030\ : std_logic;
signal \N__74025\ : std_logic;
signal \N__74022\ : std_logic;
signal \N__74021\ : std_logic;
signal \N__74018\ : std_logic;
signal \N__74015\ : std_logic;
signal \N__74010\ : std_logic;
signal \N__74003\ : std_logic;
signal \N__74000\ : std_logic;
signal \N__73997\ : std_logic;
signal \N__73990\ : std_logic;
signal \N__73981\ : std_logic;
signal \N__73978\ : std_logic;
signal \N__73975\ : std_logic;
signal \N__73972\ : std_logic;
signal \N__73967\ : std_logic;
signal \N__73964\ : std_logic;
signal \N__73957\ : std_logic;
signal \N__73944\ : std_logic;
signal \N__73943\ : std_logic;
signal \N__73940\ : std_logic;
signal \N__73939\ : std_logic;
signal \N__73936\ : std_logic;
signal \N__73933\ : std_logic;
signal \N__73930\ : std_logic;
signal \N__73927\ : std_logic;
signal \N__73924\ : std_logic;
signal \N__73921\ : std_logic;
signal \N__73918\ : std_logic;
signal \N__73915\ : std_logic;
signal \N__73908\ : std_logic;
signal \N__73905\ : std_logic;
signal \N__73902\ : std_logic;
signal \N__73901\ : std_logic;
signal \N__73900\ : std_logic;
signal \N__73899\ : std_logic;
signal \N__73896\ : std_logic;
signal \N__73893\ : std_logic;
signal \N__73890\ : std_logic;
signal \N__73887\ : std_logic;
signal \N__73884\ : std_logic;
signal \N__73881\ : std_logic;
signal \N__73876\ : std_logic;
signal \N__73873\ : std_logic;
signal \N__73868\ : std_logic;
signal \N__73863\ : std_logic;
signal \N__73862\ : std_logic;
signal \N__73861\ : std_logic;
signal \N__73858\ : std_logic;
signal \N__73855\ : std_logic;
signal \N__73854\ : std_logic;
signal \N__73851\ : std_logic;
signal \N__73848\ : std_logic;
signal \N__73843\ : std_logic;
signal \N__73840\ : std_logic;
signal \N__73837\ : std_logic;
signal \N__73834\ : std_logic;
signal \N__73831\ : std_logic;
signal \N__73828\ : std_logic;
signal \N__73825\ : std_logic;
signal \N__73822\ : std_logic;
signal \N__73817\ : std_logic;
signal \N__73814\ : std_logic;
signal \N__73809\ : std_logic;
signal \N__73806\ : std_logic;
signal \N__73803\ : std_logic;
signal \N__73800\ : std_logic;
signal \N__73797\ : std_logic;
signal \N__73796\ : std_logic;
signal \N__73793\ : std_logic;
signal \N__73790\ : std_logic;
signal \N__73787\ : std_logic;
signal \N__73784\ : std_logic;
signal \N__73779\ : std_logic;
signal \N__73776\ : std_logic;
signal \N__73773\ : std_logic;
signal \N__73772\ : std_logic;
signal \N__73769\ : std_logic;
signal \N__73766\ : std_logic;
signal \N__73763\ : std_logic;
signal \N__73760\ : std_logic;
signal \N__73755\ : std_logic;
signal \N__73752\ : std_logic;
signal \N__73751\ : std_logic;
signal \N__73750\ : std_logic;
signal \N__73747\ : std_logic;
signal \N__73744\ : std_logic;
signal \N__73741\ : std_logic;
signal \N__73738\ : std_logic;
signal \N__73735\ : std_logic;
signal \N__73734\ : std_logic;
signal \N__73727\ : std_logic;
signal \N__73724\ : std_logic;
signal \N__73719\ : std_logic;
signal \N__73718\ : std_logic;
signal \N__73717\ : std_logic;
signal \N__73716\ : std_logic;
signal \N__73715\ : std_logic;
signal \N__73714\ : std_logic;
signal \N__73711\ : std_logic;
signal \N__73710\ : std_logic;
signal \N__73709\ : std_logic;
signal \N__73708\ : std_logic;
signal \N__73707\ : std_logic;
signal \N__73706\ : std_logic;
signal \N__73705\ : std_logic;
signal \N__73704\ : std_logic;
signal \N__73703\ : std_logic;
signal \N__73702\ : std_logic;
signal \N__73697\ : std_logic;
signal \N__73696\ : std_logic;
signal \N__73695\ : std_logic;
signal \N__73694\ : std_logic;
signal \N__73693\ : std_logic;
signal \N__73692\ : std_logic;
signal \N__73691\ : std_logic;
signal \N__73690\ : std_logic;
signal \N__73689\ : std_logic;
signal \N__73688\ : std_logic;
signal \N__73687\ : std_logic;
signal \N__73686\ : std_logic;
signal \N__73685\ : std_logic;
signal \N__73684\ : std_logic;
signal \N__73681\ : std_logic;
signal \N__73670\ : std_logic;
signal \N__73669\ : std_logic;
signal \N__73668\ : std_logic;
signal \N__73667\ : std_logic;
signal \N__73666\ : std_logic;
signal \N__73665\ : std_logic;
signal \N__73662\ : std_logic;
signal \N__73659\ : std_logic;
signal \N__73658\ : std_logic;
signal \N__73655\ : std_logic;
signal \N__73652\ : std_logic;
signal \N__73651\ : std_logic;
signal \N__73644\ : std_logic;
signal \N__73641\ : std_logic;
signal \N__73630\ : std_logic;
signal \N__73623\ : std_logic;
signal \N__73620\ : std_logic;
signal \N__73615\ : std_logic;
signal \N__73612\ : std_logic;
signal \N__73611\ : std_logic;
signal \N__73610\ : std_logic;
signal \N__73609\ : std_logic;
signal \N__73608\ : std_logic;
signal \N__73605\ : std_logic;
signal \N__73602\ : std_logic;
signal \N__73599\ : std_logic;
signal \N__73598\ : std_logic;
signal \N__73597\ : std_logic;
signal \N__73596\ : std_logic;
signal \N__73595\ : std_logic;
signal \N__73590\ : std_logic;
signal \N__73587\ : std_logic;
signal \N__73582\ : std_logic;
signal \N__73579\ : std_logic;
signal \N__73576\ : std_logic;
signal \N__73573\ : std_logic;
signal \N__73570\ : std_logic;
signal \N__73567\ : std_logic;
signal \N__73564\ : std_logic;
signal \N__73561\ : std_logic;
signal \N__73558\ : std_logic;
signal \N__73551\ : std_logic;
signal \N__73548\ : std_logic;
signal \N__73543\ : std_logic;
signal \N__73534\ : std_logic;
signal \N__73529\ : std_logic;
signal \N__73526\ : std_logic;
signal \N__73523\ : std_logic;
signal \N__73522\ : std_logic;
signal \N__73521\ : std_logic;
signal \N__73520\ : std_logic;
signal \N__73519\ : std_logic;
signal \N__73518\ : std_logic;
signal \N__73513\ : std_logic;
signal \N__73506\ : std_logic;
signal \N__73503\ : std_logic;
signal \N__73500\ : std_logic;
signal \N__73497\ : std_logic;
signal \N__73492\ : std_logic;
signal \N__73489\ : std_logic;
signal \N__73484\ : std_logic;
signal \N__73479\ : std_logic;
signal \N__73472\ : std_logic;
signal \N__73467\ : std_logic;
signal \N__73464\ : std_logic;
signal \N__73461\ : std_logic;
signal \N__73458\ : std_logic;
signal \N__73453\ : std_logic;
signal \N__73450\ : std_logic;
signal \N__73447\ : std_logic;
signal \N__73444\ : std_logic;
signal \N__73441\ : std_logic;
signal \N__73436\ : std_logic;
signal \N__73431\ : std_logic;
signal \N__73424\ : std_logic;
signal \N__73401\ : std_logic;
signal \N__73400\ : std_logic;
signal \N__73397\ : std_logic;
signal \N__73396\ : std_logic;
signal \N__73393\ : std_logic;
signal \N__73392\ : std_logic;
signal \N__73389\ : std_logic;
signal \N__73386\ : std_logic;
signal \N__73383\ : std_logic;
signal \N__73380\ : std_logic;
signal \N__73377\ : std_logic;
signal \N__73374\ : std_logic;
signal \N__73369\ : std_logic;
signal \N__73366\ : std_logic;
signal \N__73361\ : std_logic;
signal \N__73356\ : std_logic;
signal \N__73353\ : std_logic;
signal \N__73350\ : std_logic;
signal \N__73349\ : std_logic;
signal \N__73348\ : std_logic;
signal \N__73347\ : std_logic;
signal \N__73346\ : std_logic;
signal \N__73343\ : std_logic;
signal \N__73338\ : std_logic;
signal \N__73337\ : std_logic;
signal \N__73336\ : std_logic;
signal \N__73335\ : std_logic;
signal \N__73332\ : std_logic;
signal \N__73331\ : std_logic;
signal \N__73330\ : std_logic;
signal \N__73327\ : std_logic;
signal \N__73326\ : std_logic;
signal \N__73321\ : std_logic;
signal \N__73316\ : std_logic;
signal \N__73313\ : std_logic;
signal \N__73308\ : std_logic;
signal \N__73307\ : std_logic;
signal \N__73304\ : std_logic;
signal \N__73301\ : std_logic;
signal \N__73300\ : std_logic;
signal \N__73299\ : std_logic;
signal \N__73298\ : std_logic;
signal \N__73295\ : std_logic;
signal \N__73294\ : std_logic;
signal \N__73293\ : std_logic;
signal \N__73292\ : std_logic;
signal \N__73291\ : std_logic;
signal \N__73290\ : std_logic;
signal \N__73289\ : std_logic;
signal \N__73286\ : std_logic;
signal \N__73283\ : std_logic;
signal \N__73280\ : std_logic;
signal \N__73277\ : std_logic;
signal \N__73276\ : std_logic;
signal \N__73273\ : std_logic;
signal \N__73270\ : std_logic;
signal \N__73267\ : std_logic;
signal \N__73264\ : std_logic;
signal \N__73261\ : std_logic;
signal \N__73258\ : std_logic;
signal \N__73255\ : std_logic;
signal \N__73250\ : std_logic;
signal \N__73245\ : std_logic;
signal \N__73242\ : std_logic;
signal \N__73239\ : std_logic;
signal \N__73234\ : std_logic;
signal \N__73229\ : std_logic;
signal \N__73226\ : std_logic;
signal \N__73223\ : std_logic;
signal \N__73220\ : std_logic;
signal \N__73215\ : std_logic;
signal \N__73214\ : std_logic;
signal \N__73211\ : std_logic;
signal \N__73210\ : std_logic;
signal \N__73209\ : std_logic;
signal \N__73208\ : std_logic;
signal \N__73207\ : std_logic;
signal \N__73202\ : std_logic;
signal \N__73201\ : std_logic;
signal \N__73196\ : std_logic;
signal \N__73187\ : std_logic;
signal \N__73182\ : std_logic;
signal \N__73179\ : std_logic;
signal \N__73176\ : std_logic;
signal \N__73173\ : std_logic;
signal \N__73170\ : std_logic;
signal \N__73167\ : std_logic;
signal \N__73160\ : std_logic;
signal \N__73157\ : std_logic;
signal \N__73156\ : std_logic;
signal \N__73155\ : std_logic;
signal \N__73154\ : std_logic;
signal \N__73153\ : std_logic;
signal \N__73150\ : std_logic;
signal \N__73147\ : std_logic;
signal \N__73144\ : std_logic;
signal \N__73137\ : std_logic;
signal \N__73134\ : std_logic;
signal \N__73131\ : std_logic;
signal \N__73124\ : std_logic;
signal \N__73121\ : std_logic;
signal \N__73118\ : std_logic;
signal \N__73113\ : std_logic;
signal \N__73110\ : std_logic;
signal \N__73103\ : std_logic;
signal \N__73096\ : std_logic;
signal \N__73083\ : std_logic;
signal \N__73082\ : std_logic;
signal \N__73081\ : std_logic;
signal \N__73078\ : std_logic;
signal \N__73075\ : std_logic;
signal \N__73072\ : std_logic;
signal \N__73067\ : std_logic;
signal \N__73064\ : std_logic;
signal \N__73059\ : std_logic;
signal \N__73056\ : std_logic;
signal \N__73055\ : std_logic;
signal \N__73052\ : std_logic;
signal \N__73049\ : std_logic;
signal \N__73046\ : std_logic;
signal \N__73043\ : std_logic;
signal \N__73038\ : std_logic;
signal \N__73035\ : std_logic;
signal \N__73034\ : std_logic;
signal \N__73033\ : std_logic;
signal \N__73030\ : std_logic;
signal \N__73027\ : std_logic;
signal \N__73024\ : std_logic;
signal \N__73021\ : std_logic;
signal \N__73020\ : std_logic;
signal \N__73015\ : std_logic;
signal \N__73012\ : std_logic;
signal \N__73009\ : std_logic;
signal \N__73006\ : std_logic;
signal \N__73003\ : std_logic;
signal \N__72996\ : std_logic;
signal \N__72993\ : std_logic;
signal \N__72992\ : std_logic;
signal \N__72991\ : std_logic;
signal \N__72990\ : std_logic;
signal \N__72989\ : std_logic;
signal \N__72986\ : std_logic;
signal \N__72983\ : std_logic;
signal \N__72982\ : std_logic;
signal \N__72981\ : std_logic;
signal \N__72980\ : std_logic;
signal \N__72979\ : std_logic;
signal \N__72978\ : std_logic;
signal \N__72977\ : std_logic;
signal \N__72974\ : std_logic;
signal \N__72971\ : std_logic;
signal \N__72968\ : std_logic;
signal \N__72967\ : std_logic;
signal \N__72966\ : std_logic;
signal \N__72965\ : std_logic;
signal \N__72964\ : std_logic;
signal \N__72961\ : std_logic;
signal \N__72956\ : std_logic;
signal \N__72949\ : std_logic;
signal \N__72946\ : std_logic;
signal \N__72943\ : std_logic;
signal \N__72942\ : std_logic;
signal \N__72941\ : std_logic;
signal \N__72940\ : std_logic;
signal \N__72939\ : std_logic;
signal \N__72938\ : std_logic;
signal \N__72937\ : std_logic;
signal \N__72936\ : std_logic;
signal \N__72935\ : std_logic;
signal \N__72932\ : std_logic;
signal \N__72929\ : std_logic;
signal \N__72926\ : std_logic;
signal \N__72925\ : std_logic;
signal \N__72924\ : std_logic;
signal \N__72923\ : std_logic;
signal \N__72920\ : std_logic;
signal \N__72917\ : std_logic;
signal \N__72912\ : std_logic;
signal \N__72909\ : std_logic;
signal \N__72906\ : std_logic;
signal \N__72903\ : std_logic;
signal \N__72900\ : std_logic;
signal \N__72899\ : std_logic;
signal \N__72898\ : std_logic;
signal \N__72893\ : std_logic;
signal \N__72890\ : std_logic;
signal \N__72887\ : std_logic;
signal \N__72884\ : std_logic;
signal \N__72881\ : std_logic;
signal \N__72880\ : std_logic;
signal \N__72875\ : std_logic;
signal \N__72872\ : std_logic;
signal \N__72869\ : std_logic;
signal \N__72866\ : std_logic;
signal \N__72863\ : std_logic;
signal \N__72862\ : std_logic;
signal \N__72861\ : std_logic;
signal \N__72860\ : std_logic;
signal \N__72857\ : std_logic;
signal \N__72848\ : std_logic;
signal \N__72845\ : std_logic;
signal \N__72838\ : std_logic;
signal \N__72835\ : std_logic;
signal \N__72832\ : std_logic;
signal \N__72829\ : std_logic;
signal \N__72826\ : std_logic;
signal \N__72821\ : std_logic;
signal \N__72816\ : std_logic;
signal \N__72813\ : std_logic;
signal \N__72810\ : std_logic;
signal \N__72805\ : std_logic;
signal \N__72800\ : std_logic;
signal \N__72797\ : std_logic;
signal \N__72792\ : std_logic;
signal \N__72789\ : std_logic;
signal \N__72786\ : std_logic;
signal \N__72781\ : std_logic;
signal \N__72774\ : std_logic;
signal \N__72771\ : std_logic;
signal \N__72768\ : std_logic;
signal \N__72765\ : std_logic;
signal \N__72762\ : std_logic;
signal \N__72759\ : std_logic;
signal \N__72754\ : std_logic;
signal \N__72751\ : std_logic;
signal \N__72748\ : std_logic;
signal \N__72745\ : std_logic;
signal \N__72740\ : std_logic;
signal \N__72737\ : std_logic;
signal \N__72734\ : std_logic;
signal \N__72729\ : std_logic;
signal \N__72722\ : std_logic;
signal \N__72717\ : std_logic;
signal \N__72712\ : std_logic;
signal \N__72705\ : std_logic;
signal \N__72702\ : std_logic;
signal \N__72693\ : std_logic;
signal \N__72690\ : std_logic;
signal \N__72689\ : std_logic;
signal \N__72686\ : std_logic;
signal \N__72683\ : std_logic;
signal \N__72682\ : std_logic;
signal \N__72681\ : std_logic;
signal \N__72678\ : std_logic;
signal \N__72675\ : std_logic;
signal \N__72672\ : std_logic;
signal \N__72669\ : std_logic;
signal \N__72666\ : std_logic;
signal \N__72663\ : std_logic;
signal \N__72660\ : std_logic;
signal \N__72657\ : std_logic;
signal \N__72654\ : std_logic;
signal \N__72651\ : std_logic;
signal \N__72642\ : std_logic;
signal \N__72639\ : std_logic;
signal \N__72638\ : std_logic;
signal \N__72635\ : std_logic;
signal \N__72632\ : std_logic;
signal \N__72631\ : std_logic;
signal \N__72626\ : std_logic;
signal \N__72623\ : std_logic;
signal \N__72620\ : std_logic;
signal \N__72617\ : std_logic;
signal \N__72612\ : std_logic;
signal \N__72609\ : std_logic;
signal \N__72606\ : std_logic;
signal \N__72603\ : std_logic;
signal \N__72600\ : std_logic;
signal \N__72597\ : std_logic;
signal \N__72594\ : std_logic;
signal \N__72591\ : std_logic;
signal \N__72588\ : std_logic;
signal \N__72587\ : std_logic;
signal \N__72586\ : std_logic;
signal \N__72585\ : std_logic;
signal \N__72582\ : std_logic;
signal \N__72581\ : std_logic;
signal \N__72578\ : std_logic;
signal \N__72577\ : std_logic;
signal \N__72574\ : std_logic;
signal \N__72571\ : std_logic;
signal \N__72570\ : std_logic;
signal \N__72567\ : std_logic;
signal \N__72564\ : std_logic;
signal \N__72563\ : std_logic;
signal \N__72560\ : std_logic;
signal \N__72559\ : std_logic;
signal \N__72556\ : std_logic;
signal \N__72553\ : std_logic;
signal \N__72550\ : std_logic;
signal \N__72547\ : std_logic;
signal \N__72542\ : std_logic;
signal \N__72539\ : std_logic;
signal \N__72536\ : std_logic;
signal \N__72533\ : std_logic;
signal \N__72530\ : std_logic;
signal \N__72529\ : std_logic;
signal \N__72528\ : std_logic;
signal \N__72521\ : std_logic;
signal \N__72518\ : std_logic;
signal \N__72515\ : std_logic;
signal \N__72508\ : std_logic;
signal \N__72503\ : std_logic;
signal \N__72500\ : std_logic;
signal \N__72489\ : std_logic;
signal \N__72486\ : std_logic;
signal \N__72483\ : std_logic;
signal \N__72482\ : std_logic;
signal \N__72479\ : std_logic;
signal \N__72476\ : std_logic;
signal \N__72473\ : std_logic;
signal \N__72472\ : std_logic;
signal \N__72469\ : std_logic;
signal \N__72468\ : std_logic;
signal \N__72465\ : std_logic;
signal \N__72464\ : std_logic;
signal \N__72463\ : std_logic;
signal \N__72460\ : std_logic;
signal \N__72457\ : std_logic;
signal \N__72454\ : std_logic;
signal \N__72451\ : std_logic;
signal \N__72448\ : std_logic;
signal \N__72445\ : std_logic;
signal \N__72442\ : std_logic;
signal \N__72439\ : std_logic;
signal \N__72436\ : std_logic;
signal \N__72433\ : std_logic;
signal \N__72430\ : std_logic;
signal \N__72417\ : std_logic;
signal \N__72414\ : std_logic;
signal \N__72413\ : std_logic;
signal \N__72410\ : std_logic;
signal \N__72407\ : std_logic;
signal \N__72404\ : std_logic;
signal \N__72401\ : std_logic;
signal \N__72398\ : std_logic;
signal \N__72397\ : std_logic;
signal \N__72396\ : std_logic;
signal \N__72393\ : std_logic;
signal \N__72390\ : std_logic;
signal \N__72387\ : std_logic;
signal \N__72384\ : std_logic;
signal \N__72377\ : std_logic;
signal \N__72372\ : std_logic;
signal \N__72371\ : std_logic;
signal \N__72370\ : std_logic;
signal \N__72367\ : std_logic;
signal \N__72366\ : std_logic;
signal \N__72361\ : std_logic;
signal \N__72360\ : std_logic;
signal \N__72357\ : std_logic;
signal \N__72354\ : std_logic;
signal \N__72351\ : std_logic;
signal \N__72348\ : std_logic;
signal \N__72347\ : std_logic;
signal \N__72342\ : std_logic;
signal \N__72337\ : std_logic;
signal \N__72334\ : std_logic;
signal \N__72329\ : std_logic;
signal \N__72326\ : std_logic;
signal \N__72321\ : std_logic;
signal \N__72320\ : std_logic;
signal \N__72319\ : std_logic;
signal \N__72318\ : std_logic;
signal \N__72315\ : std_logic;
signal \N__72310\ : std_logic;
signal \N__72309\ : std_logic;
signal \N__72306\ : std_logic;
signal \N__72303\ : std_logic;
signal \N__72300\ : std_logic;
signal \N__72299\ : std_logic;
signal \N__72296\ : std_logic;
signal \N__72293\ : std_logic;
signal \N__72288\ : std_logic;
signal \N__72285\ : std_logic;
signal \N__72284\ : std_logic;
signal \N__72283\ : std_logic;
signal \N__72280\ : std_logic;
signal \N__72277\ : std_logic;
signal \N__72274\ : std_logic;
signal \N__72271\ : std_logic;
signal \N__72268\ : std_logic;
signal \N__72265\ : std_logic;
signal \N__72252\ : std_logic;
signal \N__72251\ : std_logic;
signal \N__72246\ : std_logic;
signal \N__72243\ : std_logic;
signal \N__72242\ : std_logic;
signal \N__72239\ : std_logic;
signal \N__72238\ : std_logic;
signal \N__72237\ : std_logic;
signal \N__72234\ : std_logic;
signal \N__72231\ : std_logic;
signal \N__72226\ : std_logic;
signal \N__72219\ : std_logic;
signal \N__72216\ : std_logic;
signal \N__72215\ : std_logic;
signal \N__72214\ : std_logic;
signal \N__72211\ : std_logic;
signal \N__72210\ : std_logic;
signal \N__72207\ : std_logic;
signal \N__72206\ : std_logic;
signal \N__72203\ : std_logic;
signal \N__72200\ : std_logic;
signal \N__72197\ : std_logic;
signal \N__72196\ : std_logic;
signal \N__72195\ : std_logic;
signal \N__72192\ : std_logic;
signal \N__72187\ : std_logic;
signal \N__72182\ : std_logic;
signal \N__72179\ : std_logic;
signal \N__72176\ : std_logic;
signal \N__72165\ : std_logic;
signal \N__72162\ : std_logic;
signal \N__72161\ : std_logic;
signal \N__72158\ : std_logic;
signal \N__72155\ : std_logic;
signal \N__72154\ : std_logic;
signal \N__72153\ : std_logic;
signal \N__72152\ : std_logic;
signal \N__72149\ : std_logic;
signal \N__72146\ : std_logic;
signal \N__72143\ : std_logic;
signal \N__72138\ : std_logic;
signal \N__72135\ : std_logic;
signal \N__72130\ : std_logic;
signal \N__72123\ : std_logic;
signal \N__72120\ : std_logic;
signal \N__72117\ : std_logic;
signal \N__72114\ : std_logic;
signal \N__72111\ : std_logic;
signal \N__72110\ : std_logic;
signal \N__72107\ : std_logic;
signal \N__72104\ : std_logic;
signal \N__72103\ : std_logic;
signal \N__72100\ : std_logic;
signal \N__72095\ : std_logic;
signal \N__72090\ : std_logic;
signal \N__72089\ : std_logic;
signal \N__72088\ : std_logic;
signal \N__72085\ : std_logic;
signal \N__72082\ : std_logic;
signal \N__72079\ : std_logic;
signal \N__72078\ : std_logic;
signal \N__72075\ : std_logic;
signal \N__72072\ : std_logic;
signal \N__72067\ : std_logic;
signal \N__72060\ : std_logic;
signal \N__72057\ : std_logic;
signal \N__72054\ : std_logic;
signal \N__72051\ : std_logic;
signal \N__72050\ : std_logic;
signal \N__72049\ : std_logic;
signal \N__72046\ : std_logic;
signal \N__72041\ : std_logic;
signal \N__72036\ : std_logic;
signal \N__72033\ : std_logic;
signal \N__72032\ : std_logic;
signal \N__72029\ : std_logic;
signal \N__72026\ : std_logic;
signal \N__72021\ : std_logic;
signal \N__72018\ : std_logic;
signal \N__72017\ : std_logic;
signal \N__72014\ : std_logic;
signal \N__72011\ : std_logic;
signal \N__72006\ : std_logic;
signal \N__72003\ : std_logic;
signal \N__72002\ : std_logic;
signal \N__72001\ : std_logic;
signal \N__71998\ : std_logic;
signal \N__71995\ : std_logic;
signal \N__71992\ : std_logic;
signal \N__71989\ : std_logic;
signal \N__71988\ : std_logic;
signal \N__71981\ : std_logic;
signal \N__71978\ : std_logic;
signal \N__71975\ : std_logic;
signal \N__71970\ : std_logic;
signal \N__71969\ : std_logic;
signal \N__71968\ : std_logic;
signal \N__71967\ : std_logic;
signal \N__71966\ : std_logic;
signal \N__71963\ : std_logic;
signal \N__71960\ : std_logic;
signal \N__71959\ : std_logic;
signal \N__71958\ : std_logic;
signal \N__71957\ : std_logic;
signal \N__71954\ : std_logic;
signal \N__71953\ : std_logic;
signal \N__71950\ : std_logic;
signal \N__71947\ : std_logic;
signal \N__71946\ : std_logic;
signal \N__71945\ : std_logic;
signal \N__71944\ : std_logic;
signal \N__71943\ : std_logic;
signal \N__71940\ : std_logic;
signal \N__71939\ : std_logic;
signal \N__71938\ : std_logic;
signal \N__71937\ : std_logic;
signal \N__71936\ : std_logic;
signal \N__71931\ : std_logic;
signal \N__71928\ : std_logic;
signal \N__71925\ : std_logic;
signal \N__71922\ : std_logic;
signal \N__71921\ : std_logic;
signal \N__71918\ : std_logic;
signal \N__71917\ : std_logic;
signal \N__71916\ : std_logic;
signal \N__71915\ : std_logic;
signal \N__71914\ : std_logic;
signal \N__71913\ : std_logic;
signal \N__71910\ : std_logic;
signal \N__71907\ : std_logic;
signal \N__71906\ : std_logic;
signal \N__71903\ : std_logic;
signal \N__71902\ : std_logic;
signal \N__71897\ : std_logic;
signal \N__71894\ : std_logic;
signal \N__71891\ : std_logic;
signal \N__71888\ : std_logic;
signal \N__71887\ : std_logic;
signal \N__71884\ : std_logic;
signal \N__71879\ : std_logic;
signal \N__71876\ : std_logic;
signal \N__71875\ : std_logic;
signal \N__71872\ : std_logic;
signal \N__71867\ : std_logic;
signal \N__71866\ : std_logic;
signal \N__71863\ : std_logic;
signal \N__71860\ : std_logic;
signal \N__71855\ : std_logic;
signal \N__71850\ : std_logic;
signal \N__71847\ : std_logic;
signal \N__71842\ : std_logic;
signal \N__71837\ : std_logic;
signal \N__71834\ : std_logic;
signal \N__71831\ : std_logic;
signal \N__71828\ : std_logic;
signal \N__71825\ : std_logic;
signal \N__71822\ : std_logic;
signal \N__71817\ : std_logic;
signal \N__71816\ : std_logic;
signal \N__71811\ : std_logic;
signal \N__71808\ : std_logic;
signal \N__71805\ : std_logic;
signal \N__71802\ : std_logic;
signal \N__71799\ : std_logic;
signal \N__71796\ : std_logic;
signal \N__71793\ : std_logic;
signal \N__71790\ : std_logic;
signal \N__71787\ : std_logic;
signal \N__71782\ : std_logic;
signal \N__71781\ : std_logic;
signal \N__71778\ : std_logic;
signal \N__71773\ : std_logic;
signal \N__71768\ : std_logic;
signal \N__71763\ : std_logic;
signal \N__71762\ : std_logic;
signal \N__71761\ : std_logic;
signal \N__71758\ : std_logic;
signal \N__71753\ : std_logic;
signal \N__71744\ : std_logic;
signal \N__71741\ : std_logic;
signal \N__71734\ : std_logic;
signal \N__71731\ : std_logic;
signal \N__71726\ : std_logic;
signal \N__71723\ : std_logic;
signal \N__71720\ : std_logic;
signal \N__71715\ : std_logic;
signal \N__71712\ : std_logic;
signal \N__71709\ : std_logic;
signal \N__71706\ : std_logic;
signal \N__71701\ : std_logic;
signal \N__71692\ : std_logic;
signal \N__71679\ : std_logic;
signal \N__71676\ : std_logic;
signal \N__71675\ : std_logic;
signal \N__71674\ : std_logic;
signal \N__71673\ : std_logic;
signal \N__71670\ : std_logic;
signal \N__71667\ : std_logic;
signal \N__71662\ : std_logic;
signal \N__71659\ : std_logic;
signal \N__71656\ : std_logic;
signal \N__71653\ : std_logic;
signal \N__71646\ : std_logic;
signal \N__71645\ : std_logic;
signal \N__71642\ : std_logic;
signal \N__71639\ : std_logic;
signal \N__71636\ : std_logic;
signal \N__71635\ : std_logic;
signal \N__71632\ : std_logic;
signal \N__71631\ : std_logic;
signal \N__71628\ : std_logic;
signal \N__71627\ : std_logic;
signal \N__71624\ : std_logic;
signal \N__71621\ : std_logic;
signal \N__71618\ : std_logic;
signal \N__71615\ : std_logic;
signal \N__71612\ : std_logic;
signal \N__71609\ : std_logic;
signal \N__71606\ : std_logic;
signal \N__71603\ : std_logic;
signal \N__71598\ : std_logic;
signal \N__71589\ : std_logic;
signal \N__71588\ : std_logic;
signal \N__71585\ : std_logic;
signal \N__71582\ : std_logic;
signal \N__71579\ : std_logic;
signal \N__71576\ : std_logic;
signal \N__71573\ : std_logic;
signal \N__71572\ : std_logic;
signal \N__71569\ : std_logic;
signal \N__71566\ : std_logic;
signal \N__71563\ : std_logic;
signal \N__71560\ : std_logic;
signal \N__71553\ : std_logic;
signal \N__71552\ : std_logic;
signal \N__71549\ : std_logic;
signal \N__71546\ : std_logic;
signal \N__71545\ : std_logic;
signal \N__71544\ : std_logic;
signal \N__71543\ : std_logic;
signal \N__71542\ : std_logic;
signal \N__71539\ : std_logic;
signal \N__71538\ : std_logic;
signal \N__71537\ : std_logic;
signal \N__71536\ : std_logic;
signal \N__71533\ : std_logic;
signal \N__71530\ : std_logic;
signal \N__71529\ : std_logic;
signal \N__71526\ : std_logic;
signal \N__71523\ : std_logic;
signal \N__71520\ : std_logic;
signal \N__71519\ : std_logic;
signal \N__71516\ : std_logic;
signal \N__71513\ : std_logic;
signal \N__71510\ : std_logic;
signal \N__71507\ : std_logic;
signal \N__71506\ : std_logic;
signal \N__71505\ : std_logic;
signal \N__71504\ : std_logic;
signal \N__71499\ : std_logic;
signal \N__71496\ : std_logic;
signal \N__71493\ : std_logic;
signal \N__71490\ : std_logic;
signal \N__71487\ : std_logic;
signal \N__71484\ : std_logic;
signal \N__71483\ : std_logic;
signal \N__71482\ : std_logic;
signal \N__71477\ : std_logic;
signal \N__71474\ : std_logic;
signal \N__71473\ : std_logic;
signal \N__71472\ : std_logic;
signal \N__71471\ : std_logic;
signal \N__71468\ : std_logic;
signal \N__71465\ : std_logic;
signal \N__71462\ : std_logic;
signal \N__71459\ : std_logic;
signal \N__71458\ : std_logic;
signal \N__71457\ : std_logic;
signal \N__71456\ : std_logic;
signal \N__71455\ : std_logic;
signal \N__71454\ : std_logic;
signal \N__71451\ : std_logic;
signal \N__71448\ : std_logic;
signal \N__71445\ : std_logic;
signal \N__71442\ : std_logic;
signal \N__71437\ : std_logic;
signal \N__71432\ : std_logic;
signal \N__71429\ : std_logic;
signal \N__71428\ : std_logic;
signal \N__71425\ : std_logic;
signal \N__71418\ : std_logic;
signal \N__71409\ : std_logic;
signal \N__71406\ : std_logic;
signal \N__71403\ : std_logic;
signal \N__71398\ : std_logic;
signal \N__71395\ : std_logic;
signal \N__71394\ : std_logic;
signal \N__71391\ : std_logic;
signal \N__71388\ : std_logic;
signal \N__71379\ : std_logic;
signal \N__71376\ : std_logic;
signal \N__71373\ : std_logic;
signal \N__71372\ : std_logic;
signal \N__71369\ : std_logic;
signal \N__71366\ : std_logic;
signal \N__71355\ : std_logic;
signal \N__71352\ : std_logic;
signal \N__71351\ : std_logic;
signal \N__71350\ : std_logic;
signal \N__71349\ : std_logic;
signal \N__71348\ : std_logic;
signal \N__71347\ : std_logic;
signal \N__71344\ : std_logic;
signal \N__71341\ : std_logic;
signal \N__71338\ : std_logic;
signal \N__71333\ : std_logic;
signal \N__71330\ : std_logic;
signal \N__71321\ : std_logic;
signal \N__71310\ : std_logic;
signal \N__71295\ : std_logic;
signal \N__71292\ : std_logic;
signal \N__71289\ : std_logic;
signal \N__71286\ : std_logic;
signal \N__71283\ : std_logic;
signal \N__71280\ : std_logic;
signal \N__71277\ : std_logic;
signal \N__71274\ : std_logic;
signal \N__71271\ : std_logic;
signal \N__71270\ : std_logic;
signal \N__71269\ : std_logic;
signal \N__71268\ : std_logic;
signal \N__71265\ : std_logic;
signal \N__71260\ : std_logic;
signal \N__71257\ : std_logic;
signal \N__71254\ : std_logic;
signal \N__71247\ : std_logic;
signal \N__71246\ : std_logic;
signal \N__71243\ : std_logic;
signal \N__71242\ : std_logic;
signal \N__71239\ : std_logic;
signal \N__71236\ : std_logic;
signal \N__71233\ : std_logic;
signal \N__71230\ : std_logic;
signal \N__71225\ : std_logic;
signal \N__71220\ : std_logic;
signal \N__71219\ : std_logic;
signal \N__71216\ : std_logic;
signal \N__71213\ : std_logic;
signal \N__71210\ : std_logic;
signal \N__71209\ : std_logic;
signal \N__71206\ : std_logic;
signal \N__71203\ : std_logic;
signal \N__71200\ : std_logic;
signal \N__71197\ : std_logic;
signal \N__71192\ : std_logic;
signal \N__71187\ : std_logic;
signal \N__71184\ : std_logic;
signal \N__71181\ : std_logic;
signal \N__71178\ : std_logic;
signal \N__71177\ : std_logic;
signal \N__71176\ : std_logic;
signal \N__71175\ : std_logic;
signal \N__71172\ : std_logic;
signal \N__71169\ : std_logic;
signal \N__71166\ : std_logic;
signal \N__71163\ : std_logic;
signal \N__71158\ : std_logic;
signal \N__71155\ : std_logic;
signal \N__71148\ : std_logic;
signal \N__71145\ : std_logic;
signal \N__71142\ : std_logic;
signal \N__71139\ : std_logic;
signal \N__71136\ : std_logic;
signal \N__71133\ : std_logic;
signal \N__71130\ : std_logic;
signal \N__71127\ : std_logic;
signal \N__71126\ : std_logic;
signal \N__71123\ : std_logic;
signal \N__71120\ : std_logic;
signal \N__71119\ : std_logic;
signal \N__71118\ : std_logic;
signal \N__71117\ : std_logic;
signal \N__71116\ : std_logic;
signal \N__71115\ : std_logic;
signal \N__71114\ : std_logic;
signal \N__71113\ : std_logic;
signal \N__71110\ : std_logic;
signal \N__71107\ : std_logic;
signal \N__71104\ : std_logic;
signal \N__71101\ : std_logic;
signal \N__71100\ : std_logic;
signal \N__71099\ : std_logic;
signal \N__71096\ : std_logic;
signal \N__71095\ : std_logic;
signal \N__71094\ : std_logic;
signal \N__71093\ : std_logic;
signal \N__71092\ : std_logic;
signal \N__71091\ : std_logic;
signal \N__71088\ : std_logic;
signal \N__71081\ : std_logic;
signal \N__71080\ : std_logic;
signal \N__71079\ : std_logic;
signal \N__71078\ : std_logic;
signal \N__71077\ : std_logic;
signal \N__71068\ : std_logic;
signal \N__71065\ : std_logic;
signal \N__71062\ : std_logic;
signal \N__71059\ : std_logic;
signal \N__71054\ : std_logic;
signal \N__71051\ : std_logic;
signal \N__71046\ : std_logic;
signal \N__71041\ : std_logic;
signal \N__71036\ : std_logic;
signal \N__71033\ : std_logic;
signal \N__71032\ : std_logic;
signal \N__71031\ : std_logic;
signal \N__71030\ : std_logic;
signal \N__71027\ : std_logic;
signal \N__71024\ : std_logic;
signal \N__71019\ : std_logic;
signal \N__71016\ : std_logic;
signal \N__71005\ : std_logic;
signal \N__71002\ : std_logic;
signal \N__70999\ : std_logic;
signal \N__70994\ : std_logic;
signal \N__70989\ : std_logic;
signal \N__70982\ : std_logic;
signal \N__70971\ : std_logic;
signal \N__70968\ : std_logic;
signal \N__70965\ : std_logic;
signal \N__70962\ : std_logic;
signal \N__70959\ : std_logic;
signal \N__70958\ : std_logic;
signal \N__70955\ : std_logic;
signal \N__70952\ : std_logic;
signal \N__70949\ : std_logic;
signal \N__70946\ : std_logic;
signal \N__70943\ : std_logic;
signal \N__70940\ : std_logic;
signal \N__70937\ : std_logic;
signal \N__70932\ : std_logic;
signal \N__70929\ : std_logic;
signal \N__70926\ : std_logic;
signal \N__70923\ : std_logic;
signal \N__70922\ : std_logic;
signal \N__70919\ : std_logic;
signal \N__70916\ : std_logic;
signal \N__70915\ : std_logic;
signal \N__70910\ : std_logic;
signal \N__70907\ : std_logic;
signal \N__70902\ : std_logic;
signal \N__70899\ : std_logic;
signal \N__70896\ : std_logic;
signal \N__70893\ : std_logic;
signal \N__70890\ : std_logic;
signal \N__70887\ : std_logic;
signal \N__70886\ : std_logic;
signal \N__70885\ : std_logic;
signal \N__70880\ : std_logic;
signal \N__70877\ : std_logic;
signal \N__70876\ : std_logic;
signal \N__70873\ : std_logic;
signal \N__70870\ : std_logic;
signal \N__70867\ : std_logic;
signal \N__70864\ : std_logic;
signal \N__70861\ : std_logic;
signal \N__70854\ : std_logic;
signal \N__70851\ : std_logic;
signal \N__70850\ : std_logic;
signal \N__70849\ : std_logic;
signal \N__70848\ : std_logic;
signal \N__70847\ : std_logic;
signal \N__70844\ : std_logic;
signal \N__70841\ : std_logic;
signal \N__70838\ : std_logic;
signal \N__70835\ : std_logic;
signal \N__70832\ : std_logic;
signal \N__70827\ : std_logic;
signal \N__70818\ : std_logic;
signal \N__70815\ : std_logic;
signal \N__70812\ : std_logic;
signal \N__70809\ : std_logic;
signal \N__70808\ : std_logic;
signal \N__70805\ : std_logic;
signal \N__70802\ : std_logic;
signal \N__70799\ : std_logic;
signal \N__70796\ : std_logic;
signal \N__70793\ : std_logic;
signal \N__70788\ : std_logic;
signal \N__70787\ : std_logic;
signal \N__70784\ : std_logic;
signal \N__70781\ : std_logic;
signal \N__70778\ : std_logic;
signal \N__70775\ : std_logic;
signal \N__70774\ : std_logic;
signal \N__70771\ : std_logic;
signal \N__70768\ : std_logic;
signal \N__70765\ : std_logic;
signal \N__70760\ : std_logic;
signal \N__70757\ : std_logic;
signal \N__70754\ : std_logic;
signal \N__70749\ : std_logic;
signal \N__70746\ : std_logic;
signal \N__70743\ : std_logic;
signal \N__70742\ : std_logic;
signal \N__70741\ : std_logic;
signal \N__70738\ : std_logic;
signal \N__70735\ : std_logic;
signal \N__70732\ : std_logic;
signal \N__70727\ : std_logic;
signal \N__70724\ : std_logic;
signal \N__70721\ : std_logic;
signal \N__70716\ : std_logic;
signal \N__70715\ : std_logic;
signal \N__70712\ : std_logic;
signal \N__70709\ : std_logic;
signal \N__70706\ : std_logic;
signal \N__70701\ : std_logic;
signal \N__70698\ : std_logic;
signal \N__70695\ : std_logic;
signal \N__70694\ : std_logic;
signal \N__70691\ : std_logic;
signal \N__70688\ : std_logic;
signal \N__70683\ : std_logic;
signal \N__70680\ : std_logic;
signal \N__70677\ : std_logic;
signal \N__70674\ : std_logic;
signal \N__70673\ : std_logic;
signal \N__70672\ : std_logic;
signal \N__70669\ : std_logic;
signal \N__70666\ : std_logic;
signal \N__70663\ : std_logic;
signal \N__70660\ : std_logic;
signal \N__70659\ : std_logic;
signal \N__70658\ : std_logic;
signal \N__70655\ : std_logic;
signal \N__70652\ : std_logic;
signal \N__70649\ : std_logic;
signal \N__70646\ : std_logic;
signal \N__70645\ : std_logic;
signal \N__70642\ : std_logic;
signal \N__70637\ : std_logic;
signal \N__70632\ : std_logic;
signal \N__70627\ : std_logic;
signal \N__70620\ : std_logic;
signal \N__70619\ : std_logic;
signal \N__70618\ : std_logic;
signal \N__70615\ : std_logic;
signal \N__70612\ : std_logic;
signal \N__70609\ : std_logic;
signal \N__70602\ : std_logic;
signal \N__70599\ : std_logic;
signal \N__70598\ : std_logic;
signal \N__70595\ : std_logic;
signal \N__70592\ : std_logic;
signal \N__70591\ : std_logic;
signal \N__70588\ : std_logic;
signal \N__70585\ : std_logic;
signal \N__70582\ : std_logic;
signal \N__70575\ : std_logic;
signal \N__70572\ : std_logic;
signal \N__70571\ : std_logic;
signal \N__70568\ : std_logic;
signal \N__70565\ : std_logic;
signal \N__70562\ : std_logic;
signal \N__70559\ : std_logic;
signal \N__70556\ : std_logic;
signal \N__70551\ : std_logic;
signal \N__70550\ : std_logic;
signal \N__70549\ : std_logic;
signal \N__70548\ : std_logic;
signal \N__70545\ : std_logic;
signal \N__70542\ : std_logic;
signal \N__70537\ : std_logic;
signal \N__70534\ : std_logic;
signal \N__70531\ : std_logic;
signal \N__70528\ : std_logic;
signal \N__70527\ : std_logic;
signal \N__70524\ : std_logic;
signal \N__70519\ : std_logic;
signal \N__70516\ : std_logic;
signal \N__70513\ : std_logic;
signal \N__70506\ : std_logic;
signal \N__70505\ : std_logic;
signal \N__70502\ : std_logic;
signal \N__70499\ : std_logic;
signal \N__70498\ : std_logic;
signal \N__70495\ : std_logic;
signal \N__70492\ : std_logic;
signal \N__70489\ : std_logic;
signal \N__70482\ : std_logic;
signal \N__70479\ : std_logic;
signal \N__70476\ : std_logic;
signal \N__70473\ : std_logic;
signal \N__70470\ : std_logic;
signal \N__70469\ : std_logic;
signal \N__70466\ : std_logic;
signal \N__70463\ : std_logic;
signal \N__70458\ : std_logic;
signal \N__70455\ : std_logic;
signal \N__70452\ : std_logic;
signal \N__70449\ : std_logic;
signal \N__70446\ : std_logic;
signal \N__70445\ : std_logic;
signal \N__70444\ : std_logic;
signal \N__70443\ : std_logic;
signal \N__70440\ : std_logic;
signal \N__70439\ : std_logic;
signal \N__70432\ : std_logic;
signal \N__70429\ : std_logic;
signal \N__70426\ : std_logic;
signal \N__70425\ : std_logic;
signal \N__70422\ : std_logic;
signal \N__70417\ : std_logic;
signal \N__70414\ : std_logic;
signal \N__70411\ : std_logic;
signal \N__70408\ : std_logic;
signal \N__70401\ : std_logic;
signal \N__70400\ : std_logic;
signal \N__70397\ : std_logic;
signal \N__70394\ : std_logic;
signal \N__70391\ : std_logic;
signal \N__70388\ : std_logic;
signal \N__70387\ : std_logic;
signal \N__70384\ : std_logic;
signal \N__70381\ : std_logic;
signal \N__70378\ : std_logic;
signal \N__70373\ : std_logic;
signal \N__70368\ : std_logic;
signal \N__70365\ : std_logic;
signal \N__70362\ : std_logic;
signal \N__70359\ : std_logic;
signal \N__70356\ : std_logic;
signal \N__70353\ : std_logic;
signal \N__70352\ : std_logic;
signal \N__70349\ : std_logic;
signal \N__70348\ : std_logic;
signal \N__70347\ : std_logic;
signal \N__70344\ : std_logic;
signal \N__70341\ : std_logic;
signal \N__70338\ : std_logic;
signal \N__70335\ : std_logic;
signal \N__70332\ : std_logic;
signal \N__70329\ : std_logic;
signal \N__70328\ : std_logic;
signal \N__70325\ : std_logic;
signal \N__70322\ : std_logic;
signal \N__70319\ : std_logic;
signal \N__70316\ : std_logic;
signal \N__70313\ : std_logic;
signal \N__70310\ : std_logic;
signal \N__70299\ : std_logic;
signal \N__70298\ : std_logic;
signal \N__70297\ : std_logic;
signal \N__70294\ : std_logic;
signal \N__70291\ : std_logic;
signal \N__70288\ : std_logic;
signal \N__70285\ : std_logic;
signal \N__70284\ : std_logic;
signal \N__70281\ : std_logic;
signal \N__70278\ : std_logic;
signal \N__70277\ : std_logic;
signal \N__70274\ : std_logic;
signal \N__70271\ : std_logic;
signal \N__70268\ : std_logic;
signal \N__70265\ : std_logic;
signal \N__70264\ : std_logic;
signal \N__70261\ : std_logic;
signal \N__70258\ : std_logic;
signal \N__70253\ : std_logic;
signal \N__70250\ : std_logic;
signal \N__70247\ : std_logic;
signal \N__70244\ : std_logic;
signal \N__70233\ : std_logic;
signal \N__70230\ : std_logic;
signal \N__70229\ : std_logic;
signal \N__70226\ : std_logic;
signal \N__70225\ : std_logic;
signal \N__70222\ : std_logic;
signal \N__70219\ : std_logic;
signal \N__70216\ : std_logic;
signal \N__70215\ : std_logic;
signal \N__70212\ : std_logic;
signal \N__70209\ : std_logic;
signal \N__70206\ : std_logic;
signal \N__70203\ : std_logic;
signal \N__70194\ : std_logic;
signal \N__70193\ : std_logic;
signal \N__70188\ : std_logic;
signal \N__70187\ : std_logic;
signal \N__70186\ : std_logic;
signal \N__70183\ : std_logic;
signal \N__70180\ : std_logic;
signal \N__70179\ : std_logic;
signal \N__70178\ : std_logic;
signal \N__70175\ : std_logic;
signal \N__70174\ : std_logic;
signal \N__70173\ : std_logic;
signal \N__70172\ : std_logic;
signal \N__70171\ : std_logic;
signal \N__70170\ : std_logic;
signal \N__70169\ : std_logic;
signal \N__70168\ : std_logic;
signal \N__70167\ : std_logic;
signal \N__70166\ : std_logic;
signal \N__70165\ : std_logic;
signal \N__70164\ : std_logic;
signal \N__70159\ : std_logic;
signal \N__70156\ : std_logic;
signal \N__70155\ : std_logic;
signal \N__70154\ : std_logic;
signal \N__70153\ : std_logic;
signal \N__70152\ : std_logic;
signal \N__70151\ : std_logic;
signal \N__70150\ : std_logic;
signal \N__70149\ : std_logic;
signal \N__70148\ : std_logic;
signal \N__70147\ : std_logic;
signal \N__70146\ : std_logic;
signal \N__70145\ : std_logic;
signal \N__70144\ : std_logic;
signal \N__70143\ : std_logic;
signal \N__70142\ : std_logic;
signal \N__70141\ : std_logic;
signal \N__70140\ : std_logic;
signal \N__70139\ : std_logic;
signal \N__70138\ : std_logic;
signal \N__70131\ : std_logic;
signal \N__70128\ : std_logic;
signal \N__70121\ : std_logic;
signal \N__70116\ : std_logic;
signal \N__70107\ : std_logic;
signal \N__70102\ : std_logic;
signal \N__70097\ : std_logic;
signal \N__70094\ : std_logic;
signal \N__70091\ : std_logic;
signal \N__70088\ : std_logic;
signal \N__70087\ : std_logic;
signal \N__70084\ : std_logic;
signal \N__70083\ : std_logic;
signal \N__70082\ : std_logic;
signal \N__70081\ : std_logic;
signal \N__70080\ : std_logic;
signal \N__70079\ : std_logic;
signal \N__70078\ : std_logic;
signal \N__70075\ : std_logic;
signal \N__70070\ : std_logic;
signal \N__70063\ : std_logic;
signal \N__70058\ : std_logic;
signal \N__70055\ : std_logic;
signal \N__70048\ : std_logic;
signal \N__70045\ : std_logic;
signal \N__70038\ : std_logic;
signal \N__70031\ : std_logic;
signal \N__70024\ : std_logic;
signal \N__70023\ : std_logic;
signal \N__70022\ : std_logic;
signal \N__70019\ : std_logic;
signal \N__70018\ : std_logic;
signal \N__70017\ : std_logic;
signal \N__70016\ : std_logic;
signal \N__70015\ : std_logic;
signal \N__70014\ : std_logic;
signal \N__70005\ : std_logic;
signal \N__69998\ : std_logic;
signal \N__69993\ : std_logic;
signal \N__69988\ : std_logic;
signal \N__69979\ : std_logic;
signal \N__69974\ : std_logic;
signal \N__69969\ : std_logic;
signal \N__69966\ : std_logic;
signal \N__69963\ : std_logic;
signal \N__69954\ : std_logic;
signal \N__69951\ : std_logic;
signal \N__69946\ : std_logic;
signal \N__69941\ : std_logic;
signal \N__69938\ : std_logic;
signal \N__69935\ : std_logic;
signal \N__69928\ : std_logic;
signal \N__69925\ : std_logic;
signal \N__69920\ : std_logic;
signal \N__69917\ : std_logic;
signal \N__69912\ : std_logic;
signal \N__69903\ : std_logic;
signal \N__69902\ : std_logic;
signal \N__69899\ : std_logic;
signal \N__69898\ : std_logic;
signal \N__69895\ : std_logic;
signal \N__69894\ : std_logic;
signal \N__69891\ : std_logic;
signal \N__69888\ : std_logic;
signal \N__69885\ : std_logic;
signal \N__69884\ : std_logic;
signal \N__69881\ : std_logic;
signal \N__69878\ : std_logic;
signal \N__69873\ : std_logic;
signal \N__69870\ : std_logic;
signal \N__69867\ : std_logic;
signal \N__69862\ : std_logic;
signal \N__69861\ : std_logic;
signal \N__69860\ : std_logic;
signal \N__69857\ : std_logic;
signal \N__69852\ : std_logic;
signal \N__69847\ : std_logic;
signal \N__69844\ : std_logic;
signal \N__69837\ : std_logic;
signal \N__69834\ : std_logic;
signal \N__69833\ : std_logic;
signal \N__69832\ : std_logic;
signal \N__69829\ : std_logic;
signal \N__69826\ : std_logic;
signal \N__69825\ : std_logic;
signal \N__69822\ : std_logic;
signal \N__69819\ : std_logic;
signal \N__69814\ : std_logic;
signal \N__69811\ : std_logic;
signal \N__69804\ : std_logic;
signal \N__69801\ : std_logic;
signal \N__69800\ : std_logic;
signal \N__69797\ : std_logic;
signal \N__69794\ : std_logic;
signal \N__69793\ : std_logic;
signal \N__69792\ : std_logic;
signal \N__69789\ : std_logic;
signal \N__69788\ : std_logic;
signal \N__69785\ : std_logic;
signal \N__69780\ : std_logic;
signal \N__69777\ : std_logic;
signal \N__69774\ : std_logic;
signal \N__69765\ : std_logic;
signal \N__69762\ : std_logic;
signal \N__69761\ : std_logic;
signal \N__69760\ : std_logic;
signal \N__69759\ : std_logic;
signal \N__69758\ : std_logic;
signal \N__69755\ : std_logic;
signal \N__69752\ : std_logic;
signal \N__69747\ : std_logic;
signal \N__69744\ : std_logic;
signal \N__69741\ : std_logic;
signal \N__69738\ : std_logic;
signal \N__69735\ : std_logic;
signal \N__69732\ : std_logic;
signal \N__69729\ : std_logic;
signal \N__69728\ : std_logic;
signal \N__69725\ : std_logic;
signal \N__69720\ : std_logic;
signal \N__69717\ : std_logic;
signal \N__69714\ : std_logic;
signal \N__69709\ : std_logic;
signal \N__69702\ : std_logic;
signal \N__69701\ : std_logic;
signal \N__69700\ : std_logic;
signal \N__69697\ : std_logic;
signal \N__69694\ : std_logic;
signal \N__69693\ : std_logic;
signal \N__69690\ : std_logic;
signal \N__69687\ : std_logic;
signal \N__69684\ : std_logic;
signal \N__69681\ : std_logic;
signal \N__69672\ : std_logic;
signal \N__69669\ : std_logic;
signal \N__69666\ : std_logic;
signal \N__69663\ : std_logic;
signal \N__69660\ : std_logic;
signal \N__69657\ : std_logic;
signal \N__69654\ : std_logic;
signal \N__69651\ : std_logic;
signal \N__69648\ : std_logic;
signal \N__69645\ : std_logic;
signal \N__69644\ : std_logic;
signal \N__69641\ : std_logic;
signal \N__69640\ : std_logic;
signal \N__69637\ : std_logic;
signal \N__69634\ : std_logic;
signal \N__69631\ : std_logic;
signal \N__69630\ : std_logic;
signal \N__69627\ : std_logic;
signal \N__69624\ : std_logic;
signal \N__69619\ : std_logic;
signal \N__69616\ : std_logic;
signal \N__69609\ : std_logic;
signal \N__69608\ : std_logic;
signal \N__69605\ : std_logic;
signal \N__69602\ : std_logic;
signal \N__69599\ : std_logic;
signal \N__69596\ : std_logic;
signal \N__69593\ : std_logic;
signal \N__69590\ : std_logic;
signal \N__69585\ : std_logic;
signal \N__69584\ : std_logic;
signal \N__69583\ : std_logic;
signal \N__69582\ : std_logic;
signal \N__69581\ : std_logic;
signal \N__69580\ : std_logic;
signal \N__69577\ : std_logic;
signal \N__69574\ : std_logic;
signal \N__69567\ : std_logic;
signal \N__69564\ : std_logic;
signal \N__69561\ : std_logic;
signal \N__69558\ : std_logic;
signal \N__69557\ : std_logic;
signal \N__69554\ : std_logic;
signal \N__69551\ : std_logic;
signal \N__69550\ : std_logic;
signal \N__69549\ : std_logic;
signal \N__69548\ : std_logic;
signal \N__69547\ : std_logic;
signal \N__69546\ : std_logic;
signal \N__69543\ : std_logic;
signal \N__69540\ : std_logic;
signal \N__69537\ : std_logic;
signal \N__69532\ : std_logic;
signal \N__69525\ : std_logic;
signal \N__69522\ : std_logic;
signal \N__69519\ : std_logic;
signal \N__69504\ : std_logic;
signal \N__69501\ : std_logic;
signal \N__69500\ : std_logic;
signal \N__69495\ : std_logic;
signal \N__69492\ : std_logic;
signal \N__69491\ : std_logic;
signal \N__69488\ : std_logic;
signal \N__69485\ : std_logic;
signal \N__69482\ : std_logic;
signal \N__69481\ : std_logic;
signal \N__69480\ : std_logic;
signal \N__69475\ : std_logic;
signal \N__69472\ : std_logic;
signal \N__69469\ : std_logic;
signal \N__69462\ : std_logic;
signal \N__69461\ : std_logic;
signal \N__69460\ : std_logic;
signal \N__69459\ : std_logic;
signal \N__69454\ : std_logic;
signal \N__69451\ : std_logic;
signal \N__69450\ : std_logic;
signal \N__69447\ : std_logic;
signal \N__69444\ : std_logic;
signal \N__69441\ : std_logic;
signal \N__69438\ : std_logic;
signal \N__69437\ : std_logic;
signal \N__69434\ : std_logic;
signal \N__69431\ : std_logic;
signal \N__69426\ : std_logic;
signal \N__69423\ : std_logic;
signal \N__69420\ : std_logic;
signal \N__69415\ : std_logic;
signal \N__69412\ : std_logic;
signal \N__69411\ : std_logic;
signal \N__69410\ : std_logic;
signal \N__69407\ : std_logic;
signal \N__69402\ : std_logic;
signal \N__69399\ : std_logic;
signal \N__69396\ : std_logic;
signal \N__69387\ : std_logic;
signal \N__69384\ : std_logic;
signal \N__69381\ : std_logic;
signal \N__69380\ : std_logic;
signal \N__69377\ : std_logic;
signal \N__69376\ : std_logic;
signal \N__69373\ : std_logic;
signal \N__69370\ : std_logic;
signal \N__69367\ : std_logic;
signal \N__69364\ : std_logic;
signal \N__69363\ : std_logic;
signal \N__69362\ : std_logic;
signal \N__69355\ : std_logic;
signal \N__69354\ : std_logic;
signal \N__69351\ : std_logic;
signal \N__69348\ : std_logic;
signal \N__69345\ : std_logic;
signal \N__69342\ : std_logic;
signal \N__69337\ : std_logic;
signal \N__69330\ : std_logic;
signal \N__69329\ : std_logic;
signal \N__69326\ : std_logic;
signal \N__69325\ : std_logic;
signal \N__69322\ : std_logic;
signal \N__69321\ : std_logic;
signal \N__69320\ : std_logic;
signal \N__69317\ : std_logic;
signal \N__69314\ : std_logic;
signal \N__69313\ : std_logic;
signal \N__69310\ : std_logic;
signal \N__69305\ : std_logic;
signal \N__69302\ : std_logic;
signal \N__69301\ : std_logic;
signal \N__69298\ : std_logic;
signal \N__69295\ : std_logic;
signal \N__69288\ : std_logic;
signal \N__69285\ : std_logic;
signal \N__69276\ : std_logic;
signal \N__69275\ : std_logic;
signal \N__69272\ : std_logic;
signal \N__69267\ : std_logic;
signal \N__69264\ : std_logic;
signal \N__69263\ : std_logic;
signal \N__69262\ : std_logic;
signal \N__69255\ : std_logic;
signal \N__69252\ : std_logic;
signal \N__69249\ : std_logic;
signal \N__69246\ : std_logic;
signal \N__69243\ : std_logic;
signal \N__69240\ : std_logic;
signal \N__69237\ : std_logic;
signal \N__69236\ : std_logic;
signal \N__69235\ : std_logic;
signal \N__69228\ : std_logic;
signal \N__69227\ : std_logic;
signal \N__69226\ : std_logic;
signal \N__69225\ : std_logic;
signal \N__69224\ : std_logic;
signal \N__69223\ : std_logic;
signal \N__69220\ : std_logic;
signal \N__69215\ : std_logic;
signal \N__69212\ : std_logic;
signal \N__69211\ : std_logic;
signal \N__69210\ : std_logic;
signal \N__69205\ : std_logic;
signal \N__69204\ : std_logic;
signal \N__69201\ : std_logic;
signal \N__69200\ : std_logic;
signal \N__69199\ : std_logic;
signal \N__69196\ : std_logic;
signal \N__69195\ : std_logic;
signal \N__69194\ : std_logic;
signal \N__69191\ : std_logic;
signal \N__69186\ : std_logic;
signal \N__69185\ : std_logic;
signal \N__69184\ : std_logic;
signal \N__69183\ : std_logic;
signal \N__69182\ : std_logic;
signal \N__69181\ : std_logic;
signal \N__69180\ : std_logic;
signal \N__69177\ : std_logic;
signal \N__69174\ : std_logic;
signal \N__69171\ : std_logic;
signal \N__69170\ : std_logic;
signal \N__69167\ : std_logic;
signal \N__69166\ : std_logic;
signal \N__69163\ : std_logic;
signal \N__69162\ : std_logic;
signal \N__69161\ : std_logic;
signal \N__69158\ : std_logic;
signal \N__69157\ : std_logic;
signal \N__69156\ : std_logic;
signal \N__69151\ : std_logic;
signal \N__69150\ : std_logic;
signal \N__69147\ : std_logic;
signal \N__69144\ : std_logic;
signal \N__69141\ : std_logic;
signal \N__69136\ : std_logic;
signal \N__69129\ : std_logic;
signal \N__69124\ : std_logic;
signal \N__69121\ : std_logic;
signal \N__69118\ : std_logic;
signal \N__69117\ : std_logic;
signal \N__69112\ : std_logic;
signal \N__69109\ : std_logic;
signal \N__69104\ : std_logic;
signal \N__69101\ : std_logic;
signal \N__69098\ : std_logic;
signal \N__69095\ : std_logic;
signal \N__69092\ : std_logic;
signal \N__69091\ : std_logic;
signal \N__69088\ : std_logic;
signal \N__69085\ : std_logic;
signal \N__69078\ : std_logic;
signal \N__69075\ : std_logic;
signal \N__69072\ : std_logic;
signal \N__69069\ : std_logic;
signal \N__69068\ : std_logic;
signal \N__69065\ : std_logic;
signal \N__69062\ : std_logic;
signal \N__69059\ : std_logic;
signal \N__69050\ : std_logic;
signal \N__69047\ : std_logic;
signal \N__69044\ : std_logic;
signal \N__69041\ : std_logic;
signal \N__69038\ : std_logic;
signal \N__69035\ : std_logic;
signal \N__69032\ : std_logic;
signal \N__69025\ : std_logic;
signal \N__69022\ : std_logic;
signal \N__69019\ : std_logic;
signal \N__69012\ : std_logic;
signal \N__69007\ : std_logic;
signal \N__69000\ : std_logic;
signal \N__68995\ : std_logic;
signal \N__68982\ : std_logic;
signal \N__68979\ : std_logic;
signal \N__68976\ : std_logic;
signal \N__68973\ : std_logic;
signal \N__68970\ : std_logic;
signal \N__68969\ : std_logic;
signal \N__68966\ : std_logic;
signal \N__68963\ : std_logic;
signal \N__68960\ : std_logic;
signal \N__68959\ : std_logic;
signal \N__68958\ : std_logic;
signal \N__68957\ : std_logic;
signal \N__68954\ : std_logic;
signal \N__68951\ : std_logic;
signal \N__68948\ : std_logic;
signal \N__68945\ : std_logic;
signal \N__68942\ : std_logic;
signal \N__68931\ : std_logic;
signal \N__68928\ : std_logic;
signal \N__68927\ : std_logic;
signal \N__68924\ : std_logic;
signal \N__68923\ : std_logic;
signal \N__68920\ : std_logic;
signal \N__68917\ : std_logic;
signal \N__68914\ : std_logic;
signal \N__68911\ : std_logic;
signal \N__68908\ : std_logic;
signal \N__68901\ : std_logic;
signal \N__68900\ : std_logic;
signal \N__68895\ : std_logic;
signal \N__68892\ : std_logic;
signal \N__68889\ : std_logic;
signal \N__68886\ : std_logic;
signal \N__68883\ : std_logic;
signal \N__68880\ : std_logic;
signal \N__68879\ : std_logic;
signal \N__68876\ : std_logic;
signal \N__68873\ : std_logic;
signal \N__68870\ : std_logic;
signal \N__68867\ : std_logic;
signal \N__68864\ : std_logic;
signal \N__68861\ : std_logic;
signal \N__68858\ : std_logic;
signal \N__68855\ : std_logic;
signal \N__68850\ : std_logic;
signal \N__68849\ : std_logic;
signal \N__68848\ : std_logic;
signal \N__68847\ : std_logic;
signal \N__68846\ : std_logic;
signal \N__68845\ : std_logic;
signal \N__68844\ : std_logic;
signal \N__68843\ : std_logic;
signal \N__68842\ : std_logic;
signal \N__68841\ : std_logic;
signal \N__68840\ : std_logic;
signal \N__68837\ : std_logic;
signal \N__68832\ : std_logic;
signal \N__68829\ : std_logic;
signal \N__68826\ : std_logic;
signal \N__68821\ : std_logic;
signal \N__68814\ : std_logic;
signal \N__68811\ : std_logic;
signal \N__68796\ : std_logic;
signal \N__68795\ : std_logic;
signal \N__68794\ : std_logic;
signal \N__68793\ : std_logic;
signal \N__68790\ : std_logic;
signal \N__68787\ : std_logic;
signal \N__68782\ : std_logic;
signal \N__68781\ : std_logic;
signal \N__68780\ : std_logic;
signal \N__68777\ : std_logic;
signal \N__68774\ : std_logic;
signal \N__68771\ : std_logic;
signal \N__68766\ : std_logic;
signal \N__68757\ : std_logic;
signal \N__68756\ : std_logic;
signal \N__68753\ : std_logic;
signal \N__68752\ : std_logic;
signal \N__68751\ : std_logic;
signal \N__68750\ : std_logic;
signal \N__68749\ : std_logic;
signal \N__68746\ : std_logic;
signal \N__68743\ : std_logic;
signal \N__68740\ : std_logic;
signal \N__68737\ : std_logic;
signal \N__68734\ : std_logic;
signal \N__68733\ : std_logic;
signal \N__68732\ : std_logic;
signal \N__68729\ : std_logic;
signal \N__68728\ : std_logic;
signal \N__68727\ : std_logic;
signal \N__68726\ : std_logic;
signal \N__68723\ : std_logic;
signal \N__68716\ : std_logic;
signal \N__68713\ : std_logic;
signal \N__68710\ : std_logic;
signal \N__68707\ : std_logic;
signal \N__68702\ : std_logic;
signal \N__68699\ : std_logic;
signal \N__68696\ : std_logic;
signal \N__68679\ : std_logic;
signal \N__68678\ : std_logic;
signal \N__68677\ : std_logic;
signal \N__68672\ : std_logic;
signal \N__68671\ : std_logic;
signal \N__68670\ : std_logic;
signal \N__68669\ : std_logic;
signal \N__68666\ : std_logic;
signal \N__68663\ : std_logic;
signal \N__68660\ : std_logic;
signal \N__68655\ : std_logic;
signal \N__68646\ : std_logic;
signal \N__68645\ : std_logic;
signal \N__68642\ : std_logic;
signal \N__68639\ : std_logic;
signal \N__68634\ : std_logic;
signal \N__68633\ : std_logic;
signal \N__68628\ : std_logic;
signal \N__68625\ : std_logic;
signal \N__68624\ : std_logic;
signal \N__68623\ : std_logic;
signal \N__68622\ : std_logic;
signal \N__68619\ : std_logic;
signal \N__68612\ : std_logic;
signal \N__68607\ : std_logic;
signal \N__68604\ : std_logic;
signal \N__68601\ : std_logic;
signal \N__68600\ : std_logic;
signal \N__68597\ : std_logic;
signal \N__68594\ : std_logic;
signal \N__68593\ : std_logic;
signal \N__68588\ : std_logic;
signal \N__68585\ : std_logic;
signal \N__68582\ : std_logic;
signal \N__68579\ : std_logic;
signal \N__68576\ : std_logic;
signal \N__68571\ : std_logic;
signal \N__68570\ : std_logic;
signal \N__68567\ : std_logic;
signal \N__68564\ : std_logic;
signal \N__68559\ : std_logic;
signal \N__68556\ : std_logic;
signal \N__68555\ : std_logic;
signal \N__68552\ : std_logic;
signal \N__68549\ : std_logic;
signal \N__68546\ : std_logic;
signal \N__68545\ : std_logic;
signal \N__68544\ : std_logic;
signal \N__68543\ : std_logic;
signal \N__68542\ : std_logic;
signal \N__68539\ : std_logic;
signal \N__68536\ : std_logic;
signal \N__68533\ : std_logic;
signal \N__68532\ : std_logic;
signal \N__68531\ : std_logic;
signal \N__68528\ : std_logic;
signal \N__68527\ : std_logic;
signal \N__68524\ : std_logic;
signal \N__68521\ : std_logic;
signal \N__68518\ : std_logic;
signal \N__68513\ : std_logic;
signal \N__68512\ : std_logic;
signal \N__68511\ : std_logic;
signal \N__68510\ : std_logic;
signal \N__68507\ : std_logic;
signal \N__68504\ : std_logic;
signal \N__68501\ : std_logic;
signal \N__68498\ : std_logic;
signal \N__68497\ : std_logic;
signal \N__68496\ : std_logic;
signal \N__68495\ : std_logic;
signal \N__68490\ : std_logic;
signal \N__68485\ : std_logic;
signal \N__68482\ : std_logic;
signal \N__68477\ : std_logic;
signal \N__68472\ : std_logic;
signal \N__68467\ : std_logic;
signal \N__68464\ : std_logic;
signal \N__68459\ : std_logic;
signal \N__68442\ : std_logic;
signal \N__68441\ : std_logic;
signal \N__68438\ : std_logic;
signal \N__68437\ : std_logic;
signal \N__68434\ : std_logic;
signal \N__68433\ : std_logic;
signal \N__68432\ : std_logic;
signal \N__68429\ : std_logic;
signal \N__68426\ : std_logic;
signal \N__68423\ : std_logic;
signal \N__68422\ : std_logic;
signal \N__68419\ : std_logic;
signal \N__68416\ : std_logic;
signal \N__68411\ : std_logic;
signal \N__68408\ : std_logic;
signal \N__68405\ : std_logic;
signal \N__68402\ : std_logic;
signal \N__68399\ : std_logic;
signal \N__68396\ : std_logic;
signal \N__68395\ : std_logic;
signal \N__68390\ : std_logic;
signal \N__68387\ : std_logic;
signal \N__68382\ : std_logic;
signal \N__68379\ : std_logic;
signal \N__68370\ : std_logic;
signal \N__68367\ : std_logic;
signal \N__68366\ : std_logic;
signal \N__68365\ : std_logic;
signal \N__68362\ : std_logic;
signal \N__68359\ : std_logic;
signal \N__68356\ : std_logic;
signal \N__68353\ : std_logic;
signal \N__68350\ : std_logic;
signal \N__68349\ : std_logic;
signal \N__68346\ : std_logic;
signal \N__68343\ : std_logic;
signal \N__68340\ : std_logic;
signal \N__68337\ : std_logic;
signal \N__68334\ : std_logic;
signal \N__68331\ : std_logic;
signal \N__68328\ : std_logic;
signal \N__68319\ : std_logic;
signal \N__68316\ : std_logic;
signal \N__68313\ : std_logic;
signal \N__68312\ : std_logic;
signal \N__68311\ : std_logic;
signal \N__68308\ : std_logic;
signal \N__68305\ : std_logic;
signal \N__68302\ : std_logic;
signal \N__68295\ : std_logic;
signal \N__68292\ : std_logic;
signal \N__68289\ : std_logic;
signal \N__68286\ : std_logic;
signal \N__68283\ : std_logic;
signal \N__68280\ : std_logic;
signal \N__68279\ : std_logic;
signal \N__68278\ : std_logic;
signal \N__68275\ : std_logic;
signal \N__68270\ : std_logic;
signal \N__68267\ : std_logic;
signal \N__68262\ : std_logic;
signal \N__68261\ : std_logic;
signal \N__68258\ : std_logic;
signal \N__68255\ : std_logic;
signal \N__68252\ : std_logic;
signal \N__68247\ : std_logic;
signal \N__68244\ : std_logic;
signal \N__68241\ : std_logic;
signal \N__68240\ : std_logic;
signal \N__68237\ : std_logic;
signal \N__68232\ : std_logic;
signal \N__68229\ : std_logic;
signal \N__68228\ : std_logic;
signal \N__68223\ : std_logic;
signal \N__68220\ : std_logic;
signal \N__68217\ : std_logic;
signal \N__68216\ : std_logic;
signal \N__68215\ : std_logic;
signal \N__68212\ : std_logic;
signal \N__68209\ : std_logic;
signal \N__68206\ : std_logic;
signal \N__68203\ : std_logic;
signal \N__68200\ : std_logic;
signal \N__68197\ : std_logic;
signal \N__68190\ : std_logic;
signal \N__68189\ : std_logic;
signal \N__68186\ : std_logic;
signal \N__68183\ : std_logic;
signal \N__68180\ : std_logic;
signal \N__68177\ : std_logic;
signal \N__68174\ : std_logic;
signal \N__68171\ : std_logic;
signal \N__68168\ : std_logic;
signal \N__68163\ : std_logic;
signal \N__68162\ : std_logic;
signal \N__68161\ : std_logic;
signal \N__68160\ : std_logic;
signal \N__68157\ : std_logic;
signal \N__68150\ : std_logic;
signal \N__68145\ : std_logic;
signal \N__68142\ : std_logic;
signal \N__68141\ : std_logic;
signal \N__68140\ : std_logic;
signal \N__68137\ : std_logic;
signal \N__68132\ : std_logic;
signal \N__68127\ : std_logic;
signal \N__68126\ : std_logic;
signal \N__68123\ : std_logic;
signal \N__68122\ : std_logic;
signal \N__68121\ : std_logic;
signal \N__68120\ : std_logic;
signal \N__68117\ : std_logic;
signal \N__68114\ : std_logic;
signal \N__68111\ : std_logic;
signal \N__68110\ : std_logic;
signal \N__68109\ : std_logic;
signal \N__68108\ : std_logic;
signal \N__68105\ : std_logic;
signal \N__68102\ : std_logic;
signal \N__68097\ : std_logic;
signal \N__68096\ : std_logic;
signal \N__68095\ : std_logic;
signal \N__68094\ : std_logic;
signal \N__68093\ : std_logic;
signal \N__68090\ : std_logic;
signal \N__68083\ : std_logic;
signal \N__68082\ : std_logic;
signal \N__68081\ : std_logic;
signal \N__68078\ : std_logic;
signal \N__68073\ : std_logic;
signal \N__68068\ : std_logic;
signal \N__68063\ : std_logic;
signal \N__68058\ : std_logic;
signal \N__68053\ : std_logic;
signal \N__68040\ : std_logic;
signal \N__68039\ : std_logic;
signal \N__68038\ : std_logic;
signal \N__68035\ : std_logic;
signal \N__68034\ : std_logic;
signal \N__68031\ : std_logic;
signal \N__68030\ : std_logic;
signal \N__68029\ : std_logic;
signal \N__68028\ : std_logic;
signal \N__68025\ : std_logic;
signal \N__68022\ : std_logic;
signal \N__68019\ : std_logic;
signal \N__68014\ : std_logic;
signal \N__68009\ : std_logic;
signal \N__67998\ : std_logic;
signal \N__67995\ : std_logic;
signal \N__67992\ : std_logic;
signal \N__67989\ : std_logic;
signal \N__67986\ : std_logic;
signal \N__67985\ : std_logic;
signal \N__67984\ : std_logic;
signal \N__67981\ : std_logic;
signal \N__67978\ : std_logic;
signal \N__67975\ : std_logic;
signal \N__67972\ : std_logic;
signal \N__67969\ : std_logic;
signal \N__67968\ : std_logic;
signal \N__67967\ : std_logic;
signal \N__67964\ : std_logic;
signal \N__67959\ : std_logic;
signal \N__67956\ : std_logic;
signal \N__67953\ : std_logic;
signal \N__67944\ : std_logic;
signal \N__67943\ : std_logic;
signal \N__67942\ : std_logic;
signal \N__67941\ : std_logic;
signal \N__67938\ : std_logic;
signal \N__67935\ : std_logic;
signal \N__67934\ : std_logic;
signal \N__67931\ : std_logic;
signal \N__67928\ : std_logic;
signal \N__67925\ : std_logic;
signal \N__67922\ : std_logic;
signal \N__67919\ : std_logic;
signal \N__67916\ : std_logic;
signal \N__67915\ : std_logic;
signal \N__67914\ : std_logic;
signal \N__67911\ : std_logic;
signal \N__67908\ : std_logic;
signal \N__67903\ : std_logic;
signal \N__67900\ : std_logic;
signal \N__67895\ : std_logic;
signal \N__67884\ : std_logic;
signal \N__67883\ : std_logic;
signal \N__67880\ : std_logic;
signal \N__67877\ : std_logic;
signal \N__67874\ : std_logic;
signal \N__67873\ : std_logic;
signal \N__67870\ : std_logic;
signal \N__67867\ : std_logic;
signal \N__67864\ : std_logic;
signal \N__67863\ : std_logic;
signal \N__67862\ : std_logic;
signal \N__67859\ : std_logic;
signal \N__67856\ : std_logic;
signal \N__67853\ : std_logic;
signal \N__67850\ : std_logic;
signal \N__67847\ : std_logic;
signal \N__67844\ : std_logic;
signal \N__67841\ : std_logic;
signal \N__67838\ : std_logic;
signal \N__67835\ : std_logic;
signal \N__67824\ : std_logic;
signal \N__67821\ : std_logic;
signal \N__67820\ : std_logic;
signal \N__67819\ : std_logic;
signal \N__67816\ : std_logic;
signal \N__67813\ : std_logic;
signal \N__67810\ : std_logic;
signal \N__67805\ : std_logic;
signal \N__67802\ : std_logic;
signal \N__67797\ : std_logic;
signal \N__67794\ : std_logic;
signal \N__67793\ : std_logic;
signal \N__67792\ : std_logic;
signal \N__67789\ : std_logic;
signal \N__67786\ : std_logic;
signal \N__67783\ : std_logic;
signal \N__67780\ : std_logic;
signal \N__67773\ : std_logic;
signal \N__67770\ : std_logic;
signal \N__67767\ : std_logic;
signal \N__67764\ : std_logic;
signal \N__67761\ : std_logic;
signal \N__67758\ : std_logic;
signal \N__67755\ : std_logic;
signal \N__67752\ : std_logic;
signal \N__67749\ : std_logic;
signal \N__67748\ : std_logic;
signal \N__67745\ : std_logic;
signal \N__67742\ : std_logic;
signal \N__67739\ : std_logic;
signal \N__67736\ : std_logic;
signal \N__67733\ : std_logic;
signal \N__67730\ : std_logic;
signal \N__67725\ : std_logic;
signal \N__67722\ : std_logic;
signal \N__67719\ : std_logic;
signal \N__67716\ : std_logic;
signal \N__67713\ : std_logic;
signal \N__67710\ : std_logic;
signal \N__67707\ : std_logic;
signal \N__67706\ : std_logic;
signal \N__67703\ : std_logic;
signal \N__67700\ : std_logic;
signal \N__67695\ : std_logic;
signal \N__67692\ : std_logic;
signal \N__67689\ : std_logic;
signal \N__67686\ : std_logic;
signal \N__67683\ : std_logic;
signal \N__67680\ : std_logic;
signal \N__67677\ : std_logic;
signal \N__67674\ : std_logic;
signal \N__67671\ : std_logic;
signal \N__67668\ : std_logic;
signal \N__67665\ : std_logic;
signal \N__67664\ : std_logic;
signal \N__67661\ : std_logic;
signal \N__67658\ : std_logic;
signal \N__67657\ : std_logic;
signal \N__67652\ : std_logic;
signal \N__67649\ : std_logic;
signal \N__67648\ : std_logic;
signal \N__67645\ : std_logic;
signal \N__67644\ : std_logic;
signal \N__67641\ : std_logic;
signal \N__67640\ : std_logic;
signal \N__67637\ : std_logic;
signal \N__67634\ : std_logic;
signal \N__67631\ : std_logic;
signal \N__67628\ : std_logic;
signal \N__67625\ : std_logic;
signal \N__67622\ : std_logic;
signal \N__67621\ : std_logic;
signal \N__67620\ : std_logic;
signal \N__67617\ : std_logic;
signal \N__67614\ : std_logic;
signal \N__67607\ : std_logic;
signal \N__67602\ : std_logic;
signal \N__67593\ : std_logic;
signal \N__67592\ : std_logic;
signal \N__67591\ : std_logic;
signal \N__67588\ : std_logic;
signal \N__67585\ : std_logic;
signal \N__67582\ : std_logic;
signal \N__67577\ : std_logic;
signal \N__67574\ : std_logic;
signal \N__67571\ : std_logic;
signal \N__67566\ : std_logic;
signal \N__67563\ : std_logic;
signal \N__67560\ : std_logic;
signal \N__67559\ : std_logic;
signal \N__67556\ : std_logic;
signal \N__67553\ : std_logic;
signal \N__67552\ : std_logic;
signal \N__67551\ : std_logic;
signal \N__67550\ : std_logic;
signal \N__67549\ : std_logic;
signal \N__67544\ : std_logic;
signal \N__67539\ : std_logic;
signal \N__67536\ : std_logic;
signal \N__67533\ : std_logic;
signal \N__67532\ : std_logic;
signal \N__67529\ : std_logic;
signal \N__67522\ : std_logic;
signal \N__67519\ : std_logic;
signal \N__67516\ : std_logic;
signal \N__67513\ : std_logic;
signal \N__67506\ : std_logic;
signal \N__67505\ : std_logic;
signal \N__67502\ : std_logic;
signal \N__67501\ : std_logic;
signal \N__67500\ : std_logic;
signal \N__67499\ : std_logic;
signal \N__67496\ : std_logic;
signal \N__67493\ : std_logic;
signal \N__67492\ : std_logic;
signal \N__67491\ : std_logic;
signal \N__67488\ : std_logic;
signal \N__67483\ : std_logic;
signal \N__67480\ : std_logic;
signal \N__67477\ : std_logic;
signal \N__67472\ : std_logic;
signal \N__67461\ : std_logic;
signal \N__67458\ : std_logic;
signal \N__67455\ : std_logic;
signal \N__67452\ : std_logic;
signal \N__67449\ : std_logic;
signal \N__67446\ : std_logic;
signal \N__67443\ : std_logic;
signal \N__67440\ : std_logic;
signal \N__67437\ : std_logic;
signal \N__67434\ : std_logic;
signal \N__67431\ : std_logic;
signal \N__67428\ : std_logic;
signal \N__67425\ : std_logic;
signal \N__67422\ : std_logic;
signal \N__67419\ : std_logic;
signal \N__67416\ : std_logic;
signal \N__67415\ : std_logic;
signal \N__67412\ : std_logic;
signal \N__67409\ : std_logic;
signal \N__67406\ : std_logic;
signal \N__67403\ : std_logic;
signal \N__67398\ : std_logic;
signal \N__67395\ : std_logic;
signal \N__67392\ : std_logic;
signal \N__67389\ : std_logic;
signal \N__67386\ : std_logic;
signal \N__67383\ : std_logic;
signal \N__67380\ : std_logic;
signal \N__67377\ : std_logic;
signal \N__67376\ : std_logic;
signal \N__67373\ : std_logic;
signal \N__67370\ : std_logic;
signal \N__67365\ : std_logic;
signal \N__67362\ : std_logic;
signal \N__67361\ : std_logic;
signal \N__67358\ : std_logic;
signal \N__67355\ : std_logic;
signal \N__67352\ : std_logic;
signal \N__67351\ : std_logic;
signal \N__67348\ : std_logic;
signal \N__67345\ : std_logic;
signal \N__67342\ : std_logic;
signal \N__67335\ : std_logic;
signal \N__67332\ : std_logic;
signal \N__67329\ : std_logic;
signal \N__67328\ : std_logic;
signal \N__67327\ : std_logic;
signal \N__67324\ : std_logic;
signal \N__67321\ : std_logic;
signal \N__67318\ : std_logic;
signal \N__67315\ : std_logic;
signal \N__67314\ : std_logic;
signal \N__67313\ : std_logic;
signal \N__67310\ : std_logic;
signal \N__67307\ : std_logic;
signal \N__67304\ : std_logic;
signal \N__67301\ : std_logic;
signal \N__67298\ : std_logic;
signal \N__67297\ : std_logic;
signal \N__67296\ : std_logic;
signal \N__67287\ : std_logic;
signal \N__67284\ : std_logic;
signal \N__67281\ : std_logic;
signal \N__67278\ : std_logic;
signal \N__67275\ : std_logic;
signal \N__67272\ : std_logic;
signal \N__67269\ : std_logic;
signal \N__67260\ : std_logic;
signal \N__67257\ : std_logic;
signal \N__67256\ : std_logic;
signal \N__67255\ : std_logic;
signal \N__67252\ : std_logic;
signal \N__67251\ : std_logic;
signal \N__67250\ : std_logic;
signal \N__67249\ : std_logic;
signal \N__67248\ : std_logic;
signal \N__67243\ : std_logic;
signal \N__67240\ : std_logic;
signal \N__67235\ : std_logic;
signal \N__67230\ : std_logic;
signal \N__67223\ : std_logic;
signal \N__67218\ : std_logic;
signal \N__67215\ : std_logic;
signal \N__67214\ : std_logic;
signal \N__67213\ : std_logic;
signal \N__67212\ : std_logic;
signal \N__67209\ : std_logic;
signal \N__67204\ : std_logic;
signal \N__67201\ : std_logic;
signal \N__67194\ : std_logic;
signal \N__67193\ : std_logic;
signal \N__67190\ : std_logic;
signal \N__67187\ : std_logic;
signal \N__67184\ : std_logic;
signal \N__67181\ : std_logic;
signal \N__67180\ : std_logic;
signal \N__67177\ : std_logic;
signal \N__67174\ : std_logic;
signal \N__67171\ : std_logic;
signal \N__67164\ : std_logic;
signal \N__67163\ : std_logic;
signal \N__67160\ : std_logic;
signal \N__67157\ : std_logic;
signal \N__67152\ : std_logic;
signal \N__67151\ : std_logic;
signal \N__67150\ : std_logic;
signal \N__67149\ : std_logic;
signal \N__67148\ : std_logic;
signal \N__67147\ : std_logic;
signal \N__67144\ : std_logic;
signal \N__67141\ : std_logic;
signal \N__67140\ : std_logic;
signal \N__67137\ : std_logic;
signal \N__67128\ : std_logic;
signal \N__67125\ : std_logic;
signal \N__67122\ : std_logic;
signal \N__67121\ : std_logic;
signal \N__67118\ : std_logic;
signal \N__67115\ : std_logic;
signal \N__67112\ : std_logic;
signal \N__67109\ : std_logic;
signal \N__67106\ : std_logic;
signal \N__67099\ : std_logic;
signal \N__67096\ : std_logic;
signal \N__67089\ : std_logic;
signal \N__67086\ : std_logic;
signal \N__67083\ : std_logic;
signal \N__67082\ : std_logic;
signal \N__67079\ : std_logic;
signal \N__67076\ : std_logic;
signal \N__67071\ : std_logic;
signal \N__67070\ : std_logic;
signal \N__67067\ : std_logic;
signal \N__67064\ : std_logic;
signal \N__67061\ : std_logic;
signal \N__67056\ : std_logic;
signal \N__67055\ : std_logic;
signal \N__67052\ : std_logic;
signal \N__67049\ : std_logic;
signal \N__67046\ : std_logic;
signal \N__67043\ : std_logic;
signal \N__67038\ : std_logic;
signal \N__67037\ : std_logic;
signal \N__67034\ : std_logic;
signal \N__67033\ : std_logic;
signal \N__67030\ : std_logic;
signal \N__67027\ : std_logic;
signal \N__67024\ : std_logic;
signal \N__67021\ : std_logic;
signal \N__67018\ : std_logic;
signal \N__67015\ : std_logic;
signal \N__67012\ : std_logic;
signal \N__67005\ : std_logic;
signal \N__67002\ : std_logic;
signal \N__66999\ : std_logic;
signal \N__66998\ : std_logic;
signal \N__66995\ : std_logic;
signal \N__66992\ : std_logic;
signal \N__66987\ : std_logic;
signal \N__66986\ : std_logic;
signal \N__66985\ : std_logic;
signal \N__66984\ : std_logic;
signal \N__66979\ : std_logic;
signal \N__66976\ : std_logic;
signal \N__66973\ : std_logic;
signal \N__66970\ : std_logic;
signal \N__66965\ : std_logic;
signal \N__66962\ : std_logic;
signal \N__66957\ : std_logic;
signal \N__66954\ : std_logic;
signal \N__66951\ : std_logic;
signal \N__66950\ : std_logic;
signal \N__66947\ : std_logic;
signal \N__66944\ : std_logic;
signal \N__66939\ : std_logic;
signal \N__66936\ : std_logic;
signal \N__66933\ : std_logic;
signal \N__66930\ : std_logic;
signal \N__66929\ : std_logic;
signal \N__66926\ : std_logic;
signal \N__66923\ : std_logic;
signal \N__66920\ : std_logic;
signal \N__66919\ : std_logic;
signal \N__66916\ : std_logic;
signal \N__66913\ : std_logic;
signal \N__66910\ : std_logic;
signal \N__66903\ : std_logic;
signal \N__66900\ : std_logic;
signal \N__66899\ : std_logic;
signal \N__66898\ : std_logic;
signal \N__66897\ : std_logic;
signal \N__66894\ : std_logic;
signal \N__66893\ : std_logic;
signal \N__66890\ : std_logic;
signal \N__66887\ : std_logic;
signal \N__66884\ : std_logic;
signal \N__66881\ : std_logic;
signal \N__66878\ : std_logic;
signal \N__66875\ : std_logic;
signal \N__66872\ : std_logic;
signal \N__66871\ : std_logic;
signal \N__66864\ : std_logic;
signal \N__66863\ : std_logic;
signal \N__66858\ : std_logic;
signal \N__66855\ : std_logic;
signal \N__66852\ : std_logic;
signal \N__66849\ : std_logic;
signal \N__66846\ : std_logic;
signal \N__66841\ : std_logic;
signal \N__66838\ : std_logic;
signal \N__66831\ : std_logic;
signal \N__66828\ : std_logic;
signal \N__66827\ : std_logic;
signal \N__66824\ : std_logic;
signal \N__66821\ : std_logic;
signal \N__66818\ : std_logic;
signal \N__66813\ : std_logic;
signal \N__66812\ : std_logic;
signal \N__66811\ : std_logic;
signal \N__66808\ : std_logic;
signal \N__66807\ : std_logic;
signal \N__66802\ : std_logic;
signal \N__66799\ : std_logic;
signal \N__66796\ : std_logic;
signal \N__66793\ : std_logic;
signal \N__66790\ : std_logic;
signal \N__66787\ : std_logic;
signal \N__66784\ : std_logic;
signal \N__66781\ : std_logic;
signal \N__66776\ : std_logic;
signal \N__66771\ : std_logic;
signal \N__66768\ : std_logic;
signal \N__66765\ : std_logic;
signal \N__66762\ : std_logic;
signal \N__66759\ : std_logic;
signal \N__66756\ : std_logic;
signal \N__66753\ : std_logic;
signal \N__66752\ : std_logic;
signal \N__66751\ : std_logic;
signal \N__66750\ : std_logic;
signal \N__66747\ : std_logic;
signal \N__66746\ : std_logic;
signal \N__66743\ : std_logic;
signal \N__66740\ : std_logic;
signal \N__66737\ : std_logic;
signal \N__66734\ : std_logic;
signal \N__66731\ : std_logic;
signal \N__66724\ : std_logic;
signal \N__66721\ : std_logic;
signal \N__66714\ : std_logic;
signal \N__66711\ : std_logic;
signal \N__66710\ : std_logic;
signal \N__66709\ : std_logic;
signal \N__66706\ : std_logic;
signal \N__66703\ : std_logic;
signal \N__66700\ : std_logic;
signal \N__66697\ : std_logic;
signal \N__66694\ : std_logic;
signal \N__66687\ : std_logic;
signal \N__66684\ : std_logic;
signal \N__66681\ : std_logic;
signal \N__66678\ : std_logic;
signal \N__66675\ : std_logic;
signal \N__66672\ : std_logic;
signal \N__66669\ : std_logic;
signal \N__66666\ : std_logic;
signal \N__66663\ : std_logic;
signal \N__66662\ : std_logic;
signal \N__66661\ : std_logic;
signal \N__66658\ : std_logic;
signal \N__66655\ : std_logic;
signal \N__66654\ : std_logic;
signal \N__66651\ : std_logic;
signal \N__66650\ : std_logic;
signal \N__66647\ : std_logic;
signal \N__66644\ : std_logic;
signal \N__66641\ : std_logic;
signal \N__66638\ : std_logic;
signal \N__66637\ : std_logic;
signal \N__66634\ : std_logic;
signal \N__66629\ : std_logic;
signal \N__66624\ : std_logic;
signal \N__66621\ : std_logic;
signal \N__66612\ : std_logic;
signal \N__66609\ : std_logic;
signal \N__66608\ : std_logic;
signal \N__66605\ : std_logic;
signal \N__66602\ : std_logic;
signal \N__66597\ : std_logic;
signal \N__66594\ : std_logic;
signal \N__66593\ : std_logic;
signal \N__66590\ : std_logic;
signal \N__66587\ : std_logic;
signal \N__66584\ : std_logic;
signal \N__66579\ : std_logic;
signal \N__66576\ : std_logic;
signal \N__66573\ : std_logic;
signal \N__66570\ : std_logic;
signal \N__66569\ : std_logic;
signal \N__66566\ : std_logic;
signal \N__66565\ : std_logic;
signal \N__66562\ : std_logic;
signal \N__66559\ : std_logic;
signal \N__66556\ : std_logic;
signal \N__66553\ : std_logic;
signal \N__66552\ : std_logic;
signal \N__66549\ : std_logic;
signal \N__66546\ : std_logic;
signal \N__66543\ : std_logic;
signal \N__66540\ : std_logic;
signal \N__66537\ : std_logic;
signal \N__66532\ : std_logic;
signal \N__66525\ : std_logic;
signal \N__66522\ : std_logic;
signal \N__66521\ : std_logic;
signal \N__66518\ : std_logic;
signal \N__66517\ : std_logic;
signal \N__66514\ : std_logic;
signal \N__66511\ : std_logic;
signal \N__66506\ : std_logic;
signal \N__66501\ : std_logic;
signal \N__66500\ : std_logic;
signal \N__66497\ : std_logic;
signal \N__66496\ : std_logic;
signal \N__66495\ : std_logic;
signal \N__66492\ : std_logic;
signal \N__66487\ : std_logic;
signal \N__66484\ : std_logic;
signal \N__66481\ : std_logic;
signal \N__66478\ : std_logic;
signal \N__66475\ : std_logic;
signal \N__66470\ : std_logic;
signal \N__66465\ : std_logic;
signal \N__66464\ : std_logic;
signal \N__66461\ : std_logic;
signal \N__66458\ : std_logic;
signal \N__66455\ : std_logic;
signal \N__66452\ : std_logic;
signal \N__66447\ : std_logic;
signal \N__66444\ : std_logic;
signal \N__66441\ : std_logic;
signal \N__66438\ : std_logic;
signal \N__66435\ : std_logic;
signal \N__66432\ : std_logic;
signal \N__66431\ : std_logic;
signal \N__66430\ : std_logic;
signal \N__66427\ : std_logic;
signal \N__66426\ : std_logic;
signal \N__66425\ : std_logic;
signal \N__66422\ : std_logic;
signal \N__66419\ : std_logic;
signal \N__66416\ : std_logic;
signal \N__66411\ : std_logic;
signal \N__66408\ : std_logic;
signal \N__66403\ : std_logic;
signal \N__66396\ : std_logic;
signal \N__66393\ : std_logic;
signal \N__66392\ : std_logic;
signal \N__66389\ : std_logic;
signal \N__66386\ : std_logic;
signal \N__66381\ : std_logic;
signal \N__66378\ : std_logic;
signal \N__66375\ : std_logic;
signal \N__66372\ : std_logic;
signal \N__66369\ : std_logic;
signal \N__66366\ : std_logic;
signal \N__66365\ : std_logic;
signal \N__66364\ : std_logic;
signal \N__66361\ : std_logic;
signal \N__66356\ : std_logic;
signal \N__66355\ : std_logic;
signal \N__66352\ : std_logic;
signal \N__66349\ : std_logic;
signal \N__66346\ : std_logic;
signal \N__66339\ : std_logic;
signal \N__66336\ : std_logic;
signal \N__66335\ : std_logic;
signal \N__66334\ : std_logic;
signal \N__66333\ : std_logic;
signal \N__66330\ : std_logic;
signal \N__66327\ : std_logic;
signal \N__66322\ : std_logic;
signal \N__66315\ : std_logic;
signal \N__66312\ : std_logic;
signal \N__66309\ : std_logic;
signal \N__66306\ : std_logic;
signal \N__66303\ : std_logic;
signal \N__66302\ : std_logic;
signal \N__66299\ : std_logic;
signal \N__66296\ : std_logic;
signal \N__66293\ : std_logic;
signal \N__66288\ : std_logic;
signal \N__66285\ : std_logic;
signal \N__66282\ : std_logic;
signal \N__66279\ : std_logic;
signal \N__66276\ : std_logic;
signal \N__66273\ : std_logic;
signal \N__66272\ : std_logic;
signal \N__66271\ : std_logic;
signal \N__66268\ : std_logic;
signal \N__66265\ : std_logic;
signal \N__66262\ : std_logic;
signal \N__66259\ : std_logic;
signal \N__66256\ : std_logic;
signal \N__66253\ : std_logic;
signal \N__66246\ : std_logic;
signal \N__66243\ : std_logic;
signal \N__66242\ : std_logic;
signal \N__66239\ : std_logic;
signal \N__66236\ : std_logic;
signal \N__66233\ : std_logic;
signal \N__66228\ : std_logic;
signal \N__66227\ : std_logic;
signal \N__66224\ : std_logic;
signal \N__66221\ : std_logic;
signal \N__66220\ : std_logic;
signal \N__66217\ : std_logic;
signal \N__66214\ : std_logic;
signal \N__66211\ : std_logic;
signal \N__66208\ : std_logic;
signal \N__66205\ : std_logic;
signal \N__66202\ : std_logic;
signal \N__66199\ : std_logic;
signal \N__66196\ : std_logic;
signal \N__66189\ : std_logic;
signal \N__66186\ : std_logic;
signal \N__66183\ : std_logic;
signal \N__66180\ : std_logic;
signal \N__66177\ : std_logic;
signal \N__66174\ : std_logic;
signal \N__66173\ : std_logic;
signal \N__66170\ : std_logic;
signal \N__66167\ : std_logic;
signal \N__66162\ : std_logic;
signal \N__66161\ : std_logic;
signal \N__66160\ : std_logic;
signal \N__66157\ : std_logic;
signal \N__66154\ : std_logic;
signal \N__66151\ : std_logic;
signal \N__66146\ : std_logic;
signal \N__66143\ : std_logic;
signal \N__66138\ : std_logic;
signal \N__66135\ : std_logic;
signal \N__66134\ : std_logic;
signal \N__66133\ : std_logic;
signal \N__66130\ : std_logic;
signal \N__66125\ : std_logic;
signal \N__66122\ : std_logic;
signal \N__66117\ : std_logic;
signal \N__66116\ : std_logic;
signal \N__66113\ : std_logic;
signal \N__66110\ : std_logic;
signal \N__66107\ : std_logic;
signal \N__66102\ : std_logic;
signal \N__66099\ : std_logic;
signal \N__66098\ : std_logic;
signal \N__66097\ : std_logic;
signal \N__66096\ : std_logic;
signal \N__66093\ : std_logic;
signal \N__66090\ : std_logic;
signal \N__66087\ : std_logic;
signal \N__66084\ : std_logic;
signal \N__66081\ : std_logic;
signal \N__66078\ : std_logic;
signal \N__66073\ : std_logic;
signal \N__66070\ : std_logic;
signal \N__66063\ : std_logic;
signal \N__66060\ : std_logic;
signal \N__66057\ : std_logic;
signal \N__66054\ : std_logic;
signal \N__66053\ : std_logic;
signal \N__66052\ : std_logic;
signal \N__66049\ : std_logic;
signal \N__66044\ : std_logic;
signal \N__66041\ : std_logic;
signal \N__66038\ : std_logic;
signal \N__66033\ : std_logic;
signal \N__66032\ : std_logic;
signal \N__66027\ : std_logic;
signal \N__66024\ : std_logic;
signal \N__66021\ : std_logic;
signal \N__66018\ : std_logic;
signal \N__66017\ : std_logic;
signal \N__66016\ : std_logic;
signal \N__66011\ : std_logic;
signal \N__66010\ : std_logic;
signal \N__66007\ : std_logic;
signal \N__66006\ : std_logic;
signal \N__66003\ : std_logic;
signal \N__66000\ : std_logic;
signal \N__65995\ : std_logic;
signal \N__65988\ : std_logic;
signal \N__65987\ : std_logic;
signal \N__65984\ : std_logic;
signal \N__65981\ : std_logic;
signal \N__65980\ : std_logic;
signal \N__65977\ : std_logic;
signal \N__65972\ : std_logic;
signal \N__65969\ : std_logic;
signal \N__65964\ : std_logic;
signal \N__65961\ : std_logic;
signal \N__65960\ : std_logic;
signal \N__65959\ : std_logic;
signal \N__65956\ : std_logic;
signal \N__65953\ : std_logic;
signal \N__65950\ : std_logic;
signal \N__65947\ : std_logic;
signal \N__65944\ : std_logic;
signal \N__65941\ : std_logic;
signal \N__65938\ : std_logic;
signal \N__65931\ : std_logic;
signal \N__65928\ : std_logic;
signal \N__65927\ : std_logic;
signal \N__65924\ : std_logic;
signal \N__65921\ : std_logic;
signal \N__65918\ : std_logic;
signal \N__65915\ : std_logic;
signal \N__65910\ : std_logic;
signal \N__65907\ : std_logic;
signal \N__65904\ : std_logic;
signal \N__65903\ : std_logic;
signal \N__65902\ : std_logic;
signal \N__65899\ : std_logic;
signal \N__65896\ : std_logic;
signal \N__65893\ : std_logic;
signal \N__65888\ : std_logic;
signal \N__65885\ : std_logic;
signal \N__65884\ : std_logic;
signal \N__65881\ : std_logic;
signal \N__65878\ : std_logic;
signal \N__65875\ : std_logic;
signal \N__65872\ : std_logic;
signal \N__65869\ : std_logic;
signal \N__65862\ : std_logic;
signal \N__65861\ : std_logic;
signal \N__65858\ : std_logic;
signal \N__65855\ : std_logic;
signal \N__65854\ : std_logic;
signal \N__65853\ : std_logic;
signal \N__65850\ : std_logic;
signal \N__65847\ : std_logic;
signal \N__65846\ : std_logic;
signal \N__65841\ : std_logic;
signal \N__65836\ : std_logic;
signal \N__65835\ : std_logic;
signal \N__65832\ : std_logic;
signal \N__65829\ : std_logic;
signal \N__65826\ : std_logic;
signal \N__65823\ : std_logic;
signal \N__65814\ : std_logic;
signal \N__65811\ : std_logic;
signal \N__65808\ : std_logic;
signal \N__65805\ : std_logic;
signal \N__65802\ : std_logic;
signal \N__65799\ : std_logic;
signal \N__65798\ : std_logic;
signal \N__65795\ : std_logic;
signal \N__65792\ : std_logic;
signal \N__65787\ : std_logic;
signal \N__65786\ : std_logic;
signal \N__65783\ : std_logic;
signal \N__65780\ : std_logic;
signal \N__65779\ : std_logic;
signal \N__65776\ : std_logic;
signal \N__65773\ : std_logic;
signal \N__65772\ : std_logic;
signal \N__65769\ : std_logic;
signal \N__65766\ : std_logic;
signal \N__65763\ : std_logic;
signal \N__65760\ : std_logic;
signal \N__65757\ : std_logic;
signal \N__65748\ : std_logic;
signal \N__65747\ : std_logic;
signal \N__65744\ : std_logic;
signal \N__65741\ : std_logic;
signal \N__65738\ : std_logic;
signal \N__65735\ : std_logic;
signal \N__65732\ : std_logic;
signal \N__65729\ : std_logic;
signal \N__65726\ : std_logic;
signal \N__65721\ : std_logic;
signal \N__65718\ : std_logic;
signal \N__65717\ : std_logic;
signal \N__65714\ : std_logic;
signal \N__65711\ : std_logic;
signal \N__65706\ : std_logic;
signal \N__65705\ : std_logic;
signal \N__65704\ : std_logic;
signal \N__65703\ : std_logic;
signal \N__65698\ : std_logic;
signal \N__65697\ : std_logic;
signal \N__65696\ : std_logic;
signal \N__65691\ : std_logic;
signal \N__65688\ : std_logic;
signal \N__65685\ : std_logic;
signal \N__65682\ : std_logic;
signal \N__65679\ : std_logic;
signal \N__65678\ : std_logic;
signal \N__65675\ : std_logic;
signal \N__65670\ : std_logic;
signal \N__65667\ : std_logic;
signal \N__65664\ : std_logic;
signal \N__65655\ : std_logic;
signal \N__65654\ : std_logic;
signal \N__65651\ : std_logic;
signal \N__65646\ : std_logic;
signal \N__65643\ : std_logic;
signal \N__65640\ : std_logic;
signal \N__65639\ : std_logic;
signal \N__65638\ : std_logic;
signal \N__65637\ : std_logic;
signal \N__65634\ : std_logic;
signal \N__65633\ : std_logic;
signal \N__65632\ : std_logic;
signal \N__65631\ : std_logic;
signal \N__65630\ : std_logic;
signal \N__65627\ : std_logic;
signal \N__65624\ : std_logic;
signal \N__65621\ : std_logic;
signal \N__65618\ : std_logic;
signal \N__65613\ : std_logic;
signal \N__65608\ : std_logic;
signal \N__65595\ : std_logic;
signal \N__65592\ : std_logic;
signal \N__65591\ : std_logic;
signal \N__65588\ : std_logic;
signal \N__65585\ : std_logic;
signal \N__65580\ : std_logic;
signal \N__65577\ : std_logic;
signal \N__65576\ : std_logic;
signal \N__65573\ : std_logic;
signal \N__65570\ : std_logic;
signal \N__65567\ : std_logic;
signal \N__65564\ : std_logic;
signal \N__65561\ : std_logic;
signal \N__65558\ : std_logic;
signal \N__65553\ : std_logic;
signal \N__65550\ : std_logic;
signal \N__65549\ : std_logic;
signal \N__65546\ : std_logic;
signal \N__65543\ : std_logic;
signal \N__65538\ : std_logic;
signal \N__65535\ : std_logic;
signal \N__65532\ : std_logic;
signal \N__65529\ : std_logic;
signal \N__65526\ : std_logic;
signal \N__65525\ : std_logic;
signal \N__65522\ : std_logic;
signal \N__65519\ : std_logic;
signal \N__65516\ : std_logic;
signal \N__65511\ : std_logic;
signal \N__65510\ : std_logic;
signal \N__65507\ : std_logic;
signal \N__65504\ : std_logic;
signal \N__65501\ : std_logic;
signal \N__65498\ : std_logic;
signal \N__65493\ : std_logic;
signal \N__65492\ : std_logic;
signal \N__65489\ : std_logic;
signal \N__65486\ : std_logic;
signal \N__65481\ : std_logic;
signal \N__65478\ : std_logic;
signal \N__65475\ : std_logic;
signal \N__65472\ : std_logic;
signal \N__65469\ : std_logic;
signal \N__65466\ : std_logic;
signal \N__65463\ : std_logic;
signal \N__65460\ : std_logic;
signal \N__65457\ : std_logic;
signal \N__65454\ : std_logic;
signal \N__65453\ : std_logic;
signal \N__65450\ : std_logic;
signal \N__65447\ : std_logic;
signal \N__65444\ : std_logic;
signal \N__65441\ : std_logic;
signal \N__65436\ : std_logic;
signal \N__65435\ : std_logic;
signal \N__65430\ : std_logic;
signal \N__65427\ : std_logic;
signal \N__65426\ : std_logic;
signal \N__65423\ : std_logic;
signal \N__65420\ : std_logic;
signal \N__65419\ : std_logic;
signal \N__65416\ : std_logic;
signal \N__65413\ : std_logic;
signal \N__65410\ : std_logic;
signal \N__65407\ : std_logic;
signal \N__65406\ : std_logic;
signal \N__65405\ : std_logic;
signal \N__65398\ : std_logic;
signal \N__65395\ : std_logic;
signal \N__65392\ : std_logic;
signal \N__65385\ : std_logic;
signal \N__65382\ : std_logic;
signal \N__65379\ : std_logic;
signal \N__65376\ : std_logic;
signal \N__65373\ : std_logic;
signal \N__65370\ : std_logic;
signal \N__65369\ : std_logic;
signal \N__65368\ : std_logic;
signal \N__65365\ : std_logic;
signal \N__65362\ : std_logic;
signal \N__65359\ : std_logic;
signal \N__65356\ : std_logic;
signal \N__65353\ : std_logic;
signal \N__65350\ : std_logic;
signal \N__65347\ : std_logic;
signal \N__65344\ : std_logic;
signal \N__65337\ : std_logic;
signal \N__65336\ : std_logic;
signal \N__65335\ : std_logic;
signal \N__65332\ : std_logic;
signal \N__65331\ : std_logic;
signal \N__65328\ : std_logic;
signal \N__65327\ : std_logic;
signal \N__65324\ : std_logic;
signal \N__65319\ : std_logic;
signal \N__65316\ : std_logic;
signal \N__65313\ : std_logic;
signal \N__65304\ : std_logic;
signal \N__65301\ : std_logic;
signal \N__65298\ : std_logic;
signal \N__65297\ : std_logic;
signal \N__65296\ : std_logic;
signal \N__65295\ : std_logic;
signal \N__65292\ : std_logic;
signal \N__65287\ : std_logic;
signal \N__65286\ : std_logic;
signal \N__65283\ : std_logic;
signal \N__65278\ : std_logic;
signal \N__65275\ : std_logic;
signal \N__65272\ : std_logic;
signal \N__65269\ : std_logic;
signal \N__65266\ : std_logic;
signal \N__65263\ : std_logic;
signal \N__65260\ : std_logic;
signal \N__65253\ : std_logic;
signal \N__65250\ : std_logic;
signal \N__65247\ : std_logic;
signal \N__65244\ : std_logic;
signal \N__65241\ : std_logic;
signal \N__65238\ : std_logic;
signal \N__65235\ : std_logic;
signal \N__65232\ : std_logic;
signal \N__65229\ : std_logic;
signal \N__65226\ : std_logic;
signal \N__65223\ : std_logic;
signal \N__65222\ : std_logic;
signal \N__65221\ : std_logic;
signal \N__65220\ : std_logic;
signal \N__65217\ : std_logic;
signal \N__65214\ : std_logic;
signal \N__65209\ : std_logic;
signal \N__65202\ : std_logic;
signal \N__65201\ : std_logic;
signal \N__65200\ : std_logic;
signal \N__65197\ : std_logic;
signal \N__65194\ : std_logic;
signal \N__65193\ : std_logic;
signal \N__65190\ : std_logic;
signal \N__65185\ : std_logic;
signal \N__65184\ : std_logic;
signal \N__65181\ : std_logic;
signal \N__65178\ : std_logic;
signal \N__65175\ : std_logic;
signal \N__65172\ : std_logic;
signal \N__65163\ : std_logic;
signal \N__65160\ : std_logic;
signal \N__65157\ : std_logic;
signal \N__65154\ : std_logic;
signal \N__65151\ : std_logic;
signal \N__65150\ : std_logic;
signal \N__65147\ : std_logic;
signal \N__65144\ : std_logic;
signal \N__65143\ : std_logic;
signal \N__65140\ : std_logic;
signal \N__65137\ : std_logic;
signal \N__65134\ : std_logic;
signal \N__65127\ : std_logic;
signal \N__65126\ : std_logic;
signal \N__65121\ : std_logic;
signal \N__65118\ : std_logic;
signal \N__65115\ : std_logic;
signal \N__65112\ : std_logic;
signal \N__65111\ : std_logic;
signal \N__65110\ : std_logic;
signal \N__65109\ : std_logic;
signal \N__65108\ : std_logic;
signal \N__65105\ : std_logic;
signal \N__65102\ : std_logic;
signal \N__65097\ : std_logic;
signal \N__65096\ : std_logic;
signal \N__65093\ : std_logic;
signal \N__65088\ : std_logic;
signal \N__65085\ : std_logic;
signal \N__65082\ : std_logic;
signal \N__65079\ : std_logic;
signal \N__65074\ : std_logic;
signal \N__65073\ : std_logic;
signal \N__65070\ : std_logic;
signal \N__65069\ : std_logic;
signal \N__65068\ : std_logic;
signal \N__65065\ : std_logic;
signal \N__65062\ : std_logic;
signal \N__65059\ : std_logic;
signal \N__65056\ : std_logic;
signal \N__65051\ : std_logic;
signal \N__65040\ : std_logic;
signal \N__65039\ : std_logic;
signal \N__65036\ : std_logic;
signal \N__65035\ : std_logic;
signal \N__65032\ : std_logic;
signal \N__65029\ : std_logic;
signal \N__65026\ : std_logic;
signal \N__65023\ : std_logic;
signal \N__65020\ : std_logic;
signal \N__65017\ : std_logic;
signal \N__65010\ : std_logic;
signal \N__65009\ : std_logic;
signal \N__65006\ : std_logic;
signal \N__65003\ : std_logic;
signal \N__65000\ : std_logic;
signal \N__64997\ : std_logic;
signal \N__64994\ : std_logic;
signal \N__64989\ : std_logic;
signal \N__64988\ : std_logic;
signal \N__64987\ : std_logic;
signal \N__64986\ : std_logic;
signal \N__64983\ : std_logic;
signal \N__64980\ : std_logic;
signal \N__64977\ : std_logic;
signal \N__64974\ : std_logic;
signal \N__64971\ : std_logic;
signal \N__64968\ : std_logic;
signal \N__64967\ : std_logic;
signal \N__64966\ : std_logic;
signal \N__64965\ : std_logic;
signal \N__64962\ : std_logic;
signal \N__64959\ : std_logic;
signal \N__64956\ : std_logic;
signal \N__64953\ : std_logic;
signal \N__64950\ : std_logic;
signal \N__64947\ : std_logic;
signal \N__64944\ : std_logic;
signal \N__64939\ : std_logic;
signal \N__64936\ : std_logic;
signal \N__64931\ : std_logic;
signal \N__64928\ : std_logic;
signal \N__64923\ : std_logic;
signal \N__64914\ : std_logic;
signal \N__64911\ : std_logic;
signal \N__64908\ : std_logic;
signal \N__64905\ : std_logic;
signal \N__64902\ : std_logic;
signal \N__64901\ : std_logic;
signal \N__64898\ : std_logic;
signal \N__64897\ : std_logic;
signal \N__64894\ : std_logic;
signal \N__64891\ : std_logic;
signal \N__64888\ : std_logic;
signal \N__64885\ : std_logic;
signal \N__64884\ : std_logic;
signal \N__64883\ : std_logic;
signal \N__64880\ : std_logic;
signal \N__64877\ : std_logic;
signal \N__64874\ : std_logic;
signal \N__64873\ : std_logic;
signal \N__64868\ : std_logic;
signal \N__64863\ : std_logic;
signal \N__64860\ : std_logic;
signal \N__64857\ : std_logic;
signal \N__64854\ : std_logic;
signal \N__64851\ : std_logic;
signal \N__64848\ : std_logic;
signal \N__64839\ : std_logic;
signal \N__64838\ : std_logic;
signal \N__64835\ : std_logic;
signal \N__64834\ : std_logic;
signal \N__64831\ : std_logic;
signal \N__64828\ : std_logic;
signal \N__64827\ : std_logic;
signal \N__64824\ : std_logic;
signal \N__64821\ : std_logic;
signal \N__64820\ : std_logic;
signal \N__64819\ : std_logic;
signal \N__64818\ : std_logic;
signal \N__64817\ : std_logic;
signal \N__64814\ : std_logic;
signal \N__64811\ : std_logic;
signal \N__64808\ : std_logic;
signal \N__64805\ : std_logic;
signal \N__64796\ : std_logic;
signal \N__64793\ : std_logic;
signal \N__64788\ : std_logic;
signal \N__64779\ : std_logic;
signal \N__64778\ : std_logic;
signal \N__64777\ : std_logic;
signal \N__64774\ : std_logic;
signal \N__64773\ : std_logic;
signal \N__64772\ : std_logic;
signal \N__64769\ : std_logic;
signal \N__64768\ : std_logic;
signal \N__64765\ : std_logic;
signal \N__64764\ : std_logic;
signal \N__64761\ : std_logic;
signal \N__64756\ : std_logic;
signal \N__64755\ : std_logic;
signal \N__64752\ : std_logic;
signal \N__64749\ : std_logic;
signal \N__64746\ : std_logic;
signal \N__64743\ : std_logic;
signal \N__64738\ : std_logic;
signal \N__64737\ : std_logic;
signal \N__64734\ : std_logic;
signal \N__64733\ : std_logic;
signal \N__64728\ : std_logic;
signal \N__64725\ : std_logic;
signal \N__64724\ : std_logic;
signal \N__64719\ : std_logic;
signal \N__64716\ : std_logic;
signal \N__64713\ : std_logic;
signal \N__64710\ : std_logic;
signal \N__64705\ : std_logic;
signal \N__64702\ : std_logic;
signal \N__64697\ : std_logic;
signal \N__64686\ : std_logic;
signal \N__64683\ : std_logic;
signal \N__64680\ : std_logic;
signal \N__64677\ : std_logic;
signal \N__64674\ : std_logic;
signal \N__64673\ : std_logic;
signal \N__64670\ : std_logic;
signal \N__64667\ : std_logic;
signal \N__64662\ : std_logic;
signal \N__64659\ : std_logic;
signal \N__64656\ : std_logic;
signal \N__64655\ : std_logic;
signal \N__64652\ : std_logic;
signal \N__64649\ : std_logic;
signal \N__64644\ : std_logic;
signal \N__64641\ : std_logic;
signal \N__64638\ : std_logic;
signal \N__64635\ : std_logic;
signal \N__64634\ : std_logic;
signal \N__64633\ : std_logic;
signal \N__64630\ : std_logic;
signal \N__64625\ : std_logic;
signal \N__64622\ : std_logic;
signal \N__64619\ : std_logic;
signal \N__64614\ : std_logic;
signal \N__64613\ : std_logic;
signal \N__64610\ : std_logic;
signal \N__64607\ : std_logic;
signal \N__64606\ : std_logic;
signal \N__64605\ : std_logic;
signal \N__64602\ : std_logic;
signal \N__64599\ : std_logic;
signal \N__64596\ : std_logic;
signal \N__64593\ : std_logic;
signal \N__64590\ : std_logic;
signal \N__64585\ : std_logic;
signal \N__64582\ : std_logic;
signal \N__64581\ : std_logic;
signal \N__64578\ : std_logic;
signal \N__64573\ : std_logic;
signal \N__64570\ : std_logic;
signal \N__64563\ : std_logic;
signal \N__64562\ : std_logic;
signal \N__64557\ : std_logic;
signal \N__64554\ : std_logic;
signal \N__64551\ : std_logic;
signal \N__64548\ : std_logic;
signal \N__64545\ : std_logic;
signal \N__64544\ : std_logic;
signal \N__64541\ : std_logic;
signal \N__64538\ : std_logic;
signal \N__64535\ : std_logic;
signal \N__64532\ : std_logic;
signal \N__64531\ : std_logic;
signal \N__64530\ : std_logic;
signal \N__64529\ : std_logic;
signal \N__64524\ : std_logic;
signal \N__64521\ : std_logic;
signal \N__64516\ : std_logic;
signal \N__64513\ : std_logic;
signal \N__64506\ : std_logic;
signal \N__64503\ : std_logic;
signal \N__64502\ : std_logic;
signal \N__64501\ : std_logic;
signal \N__64498\ : std_logic;
signal \N__64495\ : std_logic;
signal \N__64492\ : std_logic;
signal \N__64491\ : std_logic;
signal \N__64490\ : std_logic;
signal \N__64487\ : std_logic;
signal \N__64484\ : std_logic;
signal \N__64481\ : std_logic;
signal \N__64478\ : std_logic;
signal \N__64475\ : std_logic;
signal \N__64472\ : std_logic;
signal \N__64465\ : std_logic;
signal \N__64458\ : std_logic;
signal \N__64457\ : std_logic;
signal \N__64454\ : std_logic;
signal \N__64451\ : std_logic;
signal \N__64450\ : std_logic;
signal \N__64447\ : std_logic;
signal \N__64444\ : std_logic;
signal \N__64441\ : std_logic;
signal \N__64440\ : std_logic;
signal \N__64437\ : std_logic;
signal \N__64434\ : std_logic;
signal \N__64431\ : std_logic;
signal \N__64428\ : std_logic;
signal \N__64423\ : std_logic;
signal \N__64416\ : std_logic;
signal \N__64413\ : std_logic;
signal \N__64410\ : std_logic;
signal \N__64409\ : std_logic;
signal \N__64406\ : std_logic;
signal \N__64403\ : std_logic;
signal \N__64400\ : std_logic;
signal \N__64397\ : std_logic;
signal \N__64394\ : std_logic;
signal \N__64389\ : std_logic;
signal \N__64386\ : std_logic;
signal \N__64383\ : std_logic;
signal \N__64380\ : std_logic;
signal \N__64377\ : std_logic;
signal \N__64374\ : std_logic;
signal \N__64373\ : std_logic;
signal \N__64370\ : std_logic;
signal \N__64367\ : std_logic;
signal \N__64364\ : std_logic;
signal \N__64361\ : std_logic;
signal \N__64360\ : std_logic;
signal \N__64355\ : std_logic;
signal \N__64352\ : std_logic;
signal \N__64347\ : std_logic;
signal \N__64346\ : std_logic;
signal \N__64345\ : std_logic;
signal \N__64342\ : std_logic;
signal \N__64341\ : std_logic;
signal \N__64340\ : std_logic;
signal \N__64337\ : std_logic;
signal \N__64334\ : std_logic;
signal \N__64331\ : std_logic;
signal \N__64328\ : std_logic;
signal \N__64325\ : std_logic;
signal \N__64322\ : std_logic;
signal \N__64317\ : std_logic;
signal \N__64314\ : std_logic;
signal \N__64311\ : std_logic;
signal \N__64306\ : std_logic;
signal \N__64303\ : std_logic;
signal \N__64300\ : std_logic;
signal \N__64293\ : std_logic;
signal \N__64290\ : std_logic;
signal \N__64287\ : std_logic;
signal \N__64284\ : std_logic;
signal \N__64283\ : std_logic;
signal \N__64280\ : std_logic;
signal \N__64275\ : std_logic;
signal \N__64272\ : std_logic;
signal \N__64269\ : std_logic;
signal \N__64266\ : std_logic;
signal \N__64263\ : std_logic;
signal \N__64262\ : std_logic;
signal \N__64261\ : std_logic;
signal \N__64260\ : std_logic;
signal \N__64259\ : std_logic;
signal \N__64256\ : std_logic;
signal \N__64251\ : std_logic;
signal \N__64246\ : std_logic;
signal \N__64239\ : std_logic;
signal \N__64236\ : std_logic;
signal \N__64233\ : std_logic;
signal \N__64230\ : std_logic;
signal \N__64229\ : std_logic;
signal \N__64226\ : std_logic;
signal \N__64223\ : std_logic;
signal \N__64220\ : std_logic;
signal \N__64217\ : std_logic;
signal \N__64212\ : std_logic;
signal \N__64211\ : std_logic;
signal \N__64206\ : std_logic;
signal \N__64203\ : std_logic;
signal \N__64200\ : std_logic;
signal \N__64197\ : std_logic;
signal \N__64194\ : std_logic;
signal \N__64191\ : std_logic;
signal \N__64188\ : std_logic;
signal \N__64185\ : std_logic;
signal \N__64182\ : std_logic;
signal \N__64179\ : std_logic;
signal \N__64178\ : std_logic;
signal \N__64177\ : std_logic;
signal \N__64174\ : std_logic;
signal \N__64169\ : std_logic;
signal \N__64168\ : std_logic;
signal \N__64165\ : std_logic;
signal \N__64162\ : std_logic;
signal \N__64159\ : std_logic;
signal \N__64158\ : std_logic;
signal \N__64153\ : std_logic;
signal \N__64148\ : std_logic;
signal \N__64143\ : std_logic;
signal \N__64140\ : std_logic;
signal \N__64139\ : std_logic;
signal \N__64138\ : std_logic;
signal \N__64135\ : std_logic;
signal \N__64134\ : std_logic;
signal \N__64133\ : std_logic;
signal \N__64130\ : std_logic;
signal \N__64127\ : std_logic;
signal \N__64124\ : std_logic;
signal \N__64121\ : std_logic;
signal \N__64118\ : std_logic;
signal \N__64115\ : std_logic;
signal \N__64112\ : std_logic;
signal \N__64107\ : std_logic;
signal \N__64104\ : std_logic;
signal \N__64099\ : std_logic;
signal \N__64096\ : std_logic;
signal \N__64089\ : std_logic;
signal \N__64086\ : std_logic;
signal \N__64085\ : std_logic;
signal \N__64082\ : std_logic;
signal \N__64079\ : std_logic;
signal \N__64076\ : std_logic;
signal \N__64073\ : std_logic;
signal \N__64068\ : std_logic;
signal \N__64065\ : std_logic;
signal \N__64062\ : std_logic;
signal \N__64059\ : std_logic;
signal \N__64056\ : std_logic;
signal \N__64053\ : std_logic;
signal \N__64050\ : std_logic;
signal \N__64049\ : std_logic;
signal \N__64048\ : std_logic;
signal \N__64045\ : std_logic;
signal \N__64042\ : std_logic;
signal \N__64039\ : std_logic;
signal \N__64034\ : std_logic;
signal \N__64033\ : std_logic;
signal \N__64030\ : std_logic;
signal \N__64027\ : std_logic;
signal \N__64024\ : std_logic;
signal \N__64017\ : std_logic;
signal \N__64014\ : std_logic;
signal \N__64013\ : std_logic;
signal \N__64012\ : std_logic;
signal \N__64009\ : std_logic;
signal \N__64008\ : std_logic;
signal \N__64007\ : std_logic;
signal \N__64006\ : std_logic;
signal \N__64003\ : std_logic;
signal \N__64000\ : std_logic;
signal \N__63997\ : std_logic;
signal \N__63994\ : std_logic;
signal \N__63989\ : std_logic;
signal \N__63986\ : std_logic;
signal \N__63983\ : std_logic;
signal \N__63972\ : std_logic;
signal \N__63969\ : std_logic;
signal \N__63966\ : std_logic;
signal \N__63965\ : std_logic;
signal \N__63962\ : std_logic;
signal \N__63961\ : std_logic;
signal \N__63958\ : std_logic;
signal \N__63955\ : std_logic;
signal \N__63952\ : std_logic;
signal \N__63945\ : std_logic;
signal \N__63942\ : std_logic;
signal \N__63939\ : std_logic;
signal \N__63936\ : std_logic;
signal \N__63933\ : std_logic;
signal \N__63932\ : std_logic;
signal \N__63929\ : std_logic;
signal \N__63926\ : std_logic;
signal \N__63921\ : std_logic;
signal \N__63918\ : std_logic;
signal \N__63917\ : std_logic;
signal \N__63914\ : std_logic;
signal \N__63911\ : std_logic;
signal \N__63908\ : std_logic;
signal \N__63907\ : std_logic;
signal \N__63906\ : std_logic;
signal \N__63903\ : std_logic;
signal \N__63900\ : std_logic;
signal \N__63895\ : std_logic;
signal \N__63888\ : std_logic;
signal \N__63885\ : std_logic;
signal \N__63882\ : std_logic;
signal \N__63879\ : std_logic;
signal \N__63878\ : std_logic;
signal \N__63877\ : std_logic;
signal \N__63874\ : std_logic;
signal \N__63871\ : std_logic;
signal \N__63868\ : std_logic;
signal \N__63865\ : std_logic;
signal \N__63860\ : std_logic;
signal \N__63855\ : std_logic;
signal \N__63852\ : std_logic;
signal \N__63849\ : std_logic;
signal \N__63848\ : std_logic;
signal \N__63847\ : std_logic;
signal \N__63846\ : std_logic;
signal \N__63843\ : std_logic;
signal \N__63838\ : std_logic;
signal \N__63835\ : std_logic;
signal \N__63828\ : std_logic;
signal \N__63825\ : std_logic;
signal \N__63824\ : std_logic;
signal \N__63821\ : std_logic;
signal \N__63818\ : std_logic;
signal \N__63813\ : std_logic;
signal \N__63810\ : std_logic;
signal \N__63807\ : std_logic;
signal \N__63804\ : std_logic;
signal \N__63803\ : std_logic;
signal \N__63798\ : std_logic;
signal \N__63795\ : std_logic;
signal \N__63792\ : std_logic;
signal \N__63791\ : std_logic;
signal \N__63790\ : std_logic;
signal \N__63789\ : std_logic;
signal \N__63788\ : std_logic;
signal \N__63787\ : std_logic;
signal \N__63786\ : std_logic;
signal \N__63783\ : std_logic;
signal \N__63782\ : std_logic;
signal \N__63779\ : std_logic;
signal \N__63776\ : std_logic;
signal \N__63771\ : std_logic;
signal \N__63768\ : std_logic;
signal \N__63765\ : std_logic;
signal \N__63762\ : std_logic;
signal \N__63759\ : std_logic;
signal \N__63750\ : std_logic;
signal \N__63741\ : std_logic;
signal \N__63740\ : std_logic;
signal \N__63739\ : std_logic;
signal \N__63736\ : std_logic;
signal \N__63735\ : std_logic;
signal \N__63732\ : std_logic;
signal \N__63731\ : std_logic;
signal \N__63728\ : std_logic;
signal \N__63727\ : std_logic;
signal \N__63724\ : std_logic;
signal \N__63719\ : std_logic;
signal \N__63716\ : std_logic;
signal \N__63713\ : std_logic;
signal \N__63710\ : std_logic;
signal \N__63705\ : std_logic;
signal \N__63702\ : std_logic;
signal \N__63697\ : std_logic;
signal \N__63694\ : std_logic;
signal \N__63687\ : std_logic;
signal \N__63686\ : std_logic;
signal \N__63685\ : std_logic;
signal \N__63684\ : std_logic;
signal \N__63681\ : std_logic;
signal \N__63680\ : std_logic;
signal \N__63677\ : std_logic;
signal \N__63672\ : std_logic;
signal \N__63669\ : std_logic;
signal \N__63666\ : std_logic;
signal \N__63657\ : std_logic;
signal \N__63654\ : std_logic;
signal \N__63653\ : std_logic;
signal \N__63650\ : std_logic;
signal \N__63647\ : std_logic;
signal \N__63642\ : std_logic;
signal \N__63639\ : std_logic;
signal \N__63636\ : std_logic;
signal \N__63635\ : std_logic;
signal \N__63634\ : std_logic;
signal \N__63631\ : std_logic;
signal \N__63626\ : std_logic;
signal \N__63621\ : std_logic;
signal \N__63618\ : std_logic;
signal \N__63615\ : std_logic;
signal \N__63612\ : std_logic;
signal \N__63609\ : std_logic;
signal \N__63606\ : std_logic;
signal \N__63603\ : std_logic;
signal \N__63600\ : std_logic;
signal \N__63599\ : std_logic;
signal \N__63598\ : std_logic;
signal \N__63595\ : std_logic;
signal \N__63592\ : std_logic;
signal \N__63589\ : std_logic;
signal \N__63582\ : std_logic;
signal \N__63579\ : std_logic;
signal \N__63576\ : std_logic;
signal \N__63573\ : std_logic;
signal \N__63570\ : std_logic;
signal \N__63567\ : std_logic;
signal \N__63564\ : std_logic;
signal \N__63561\ : std_logic;
signal \N__63560\ : std_logic;
signal \N__63557\ : std_logic;
signal \N__63554\ : std_logic;
signal \N__63551\ : std_logic;
signal \N__63548\ : std_logic;
signal \N__63543\ : std_logic;
signal \N__63542\ : std_logic;
signal \N__63539\ : std_logic;
signal \N__63536\ : std_logic;
signal \N__63533\ : std_logic;
signal \N__63530\ : std_logic;
signal \N__63527\ : std_logic;
signal \N__63524\ : std_logic;
signal \N__63523\ : std_logic;
signal \N__63522\ : std_logic;
signal \N__63517\ : std_logic;
signal \N__63512\ : std_logic;
signal \N__63507\ : std_logic;
signal \N__63506\ : std_logic;
signal \N__63503\ : std_logic;
signal \N__63500\ : std_logic;
signal \N__63499\ : std_logic;
signal \N__63496\ : std_logic;
signal \N__63493\ : std_logic;
signal \N__63490\ : std_logic;
signal \N__63487\ : std_logic;
signal \N__63484\ : std_logic;
signal \N__63479\ : std_logic;
signal \N__63474\ : std_logic;
signal \N__63471\ : std_logic;
signal \N__63468\ : std_logic;
signal \N__63465\ : std_logic;
signal \N__63464\ : std_logic;
signal \N__63461\ : std_logic;
signal \N__63458\ : std_logic;
signal \N__63453\ : std_logic;
signal \N__63450\ : std_logic;
signal \N__63447\ : std_logic;
signal \N__63444\ : std_logic;
signal \N__63441\ : std_logic;
signal \N__63440\ : std_logic;
signal \N__63437\ : std_logic;
signal \N__63434\ : std_logic;
signal \N__63431\ : std_logic;
signal \N__63430\ : std_logic;
signal \N__63427\ : std_logic;
signal \N__63424\ : std_logic;
signal \N__63421\ : std_logic;
signal \N__63418\ : std_logic;
signal \N__63413\ : std_logic;
signal \N__63412\ : std_logic;
signal \N__63409\ : std_logic;
signal \N__63406\ : std_logic;
signal \N__63403\ : std_logic;
signal \N__63400\ : std_logic;
signal \N__63397\ : std_logic;
signal \N__63394\ : std_logic;
signal \N__63391\ : std_logic;
signal \N__63388\ : std_logic;
signal \N__63381\ : std_logic;
signal \N__63380\ : std_logic;
signal \N__63379\ : std_logic;
signal \N__63378\ : std_logic;
signal \N__63375\ : std_logic;
signal \N__63372\ : std_logic;
signal \N__63367\ : std_logic;
signal \N__63364\ : std_logic;
signal \N__63359\ : std_logic;
signal \N__63356\ : std_logic;
signal \N__63353\ : std_logic;
signal \N__63348\ : std_logic;
signal \N__63347\ : std_logic;
signal \N__63346\ : std_logic;
signal \N__63345\ : std_logic;
signal \N__63342\ : std_logic;
signal \N__63339\ : std_logic;
signal \N__63332\ : std_logic;
signal \N__63329\ : std_logic;
signal \N__63328\ : std_logic;
signal \N__63325\ : std_logic;
signal \N__63322\ : std_logic;
signal \N__63319\ : std_logic;
signal \N__63316\ : std_logic;
signal \N__63313\ : std_logic;
signal \N__63306\ : std_logic;
signal \N__63303\ : std_logic;
signal \N__63300\ : std_logic;
signal \N__63299\ : std_logic;
signal \N__63296\ : std_logic;
signal \N__63295\ : std_logic;
signal \N__63292\ : std_logic;
signal \N__63289\ : std_logic;
signal \N__63286\ : std_logic;
signal \N__63279\ : std_logic;
signal \N__63276\ : std_logic;
signal \N__63273\ : std_logic;
signal \N__63270\ : std_logic;
signal \N__63267\ : std_logic;
signal \N__63264\ : std_logic;
signal \N__63263\ : std_logic;
signal \N__63260\ : std_logic;
signal \N__63257\ : std_logic;
signal \N__63254\ : std_logic;
signal \N__63251\ : std_logic;
signal \N__63246\ : std_logic;
signal \N__63243\ : std_logic;
signal \N__63242\ : std_logic;
signal \N__63241\ : std_logic;
signal \N__63240\ : std_logic;
signal \N__63237\ : std_logic;
signal \N__63234\ : std_logic;
signal \N__63231\ : std_logic;
signal \N__63230\ : std_logic;
signal \N__63227\ : std_logic;
signal \N__63226\ : std_logic;
signal \N__63223\ : std_logic;
signal \N__63218\ : std_logic;
signal \N__63215\ : std_logic;
signal \N__63212\ : std_logic;
signal \N__63211\ : std_logic;
signal \N__63208\ : std_logic;
signal \N__63203\ : std_logic;
signal \N__63198\ : std_logic;
signal \N__63195\ : std_logic;
signal \N__63192\ : std_logic;
signal \N__63185\ : std_logic;
signal \N__63182\ : std_logic;
signal \N__63179\ : std_logic;
signal \N__63174\ : std_logic;
signal \N__63171\ : std_logic;
signal \N__63170\ : std_logic;
signal \N__63167\ : std_logic;
signal \N__63164\ : std_logic;
signal \N__63159\ : std_logic;
signal \N__63156\ : std_logic;
signal \N__63153\ : std_logic;
signal \N__63152\ : std_logic;
signal \N__63149\ : std_logic;
signal \N__63148\ : std_logic;
signal \N__63145\ : std_logic;
signal \N__63142\ : std_logic;
signal \N__63141\ : std_logic;
signal \N__63138\ : std_logic;
signal \N__63135\ : std_logic;
signal \N__63132\ : std_logic;
signal \N__63129\ : std_logic;
signal \N__63120\ : std_logic;
signal \N__63117\ : std_logic;
signal \N__63114\ : std_logic;
signal \N__63111\ : std_logic;
signal \N__63108\ : std_logic;
signal \N__63107\ : std_logic;
signal \N__63102\ : std_logic;
signal \N__63099\ : std_logic;
signal \N__63096\ : std_logic;
signal \N__63093\ : std_logic;
signal \N__63090\ : std_logic;
signal \N__63089\ : std_logic;
signal \N__63086\ : std_logic;
signal \N__63083\ : std_logic;
signal \N__63080\ : std_logic;
signal \N__63077\ : std_logic;
signal \N__63074\ : std_logic;
signal \N__63069\ : std_logic;
signal \N__63066\ : std_logic;
signal \N__63063\ : std_logic;
signal \N__63060\ : std_logic;
signal \N__63057\ : std_logic;
signal \N__63054\ : std_logic;
signal \N__63051\ : std_logic;
signal \N__63048\ : std_logic;
signal \N__63045\ : std_logic;
signal \N__63042\ : std_logic;
signal \N__63039\ : std_logic;
signal \N__63036\ : std_logic;
signal \N__63033\ : std_logic;
signal \N__63032\ : std_logic;
signal \N__63029\ : std_logic;
signal \N__63026\ : std_logic;
signal \N__63021\ : std_logic;
signal \N__63018\ : std_logic;
signal \N__63015\ : std_logic;
signal \N__63012\ : std_logic;
signal \N__63011\ : std_logic;
signal \N__63008\ : std_logic;
signal \N__63005\ : std_logic;
signal \N__63002\ : std_logic;
signal \N__62999\ : std_logic;
signal \N__62994\ : std_logic;
signal \N__62991\ : std_logic;
signal \N__62988\ : std_logic;
signal \N__62985\ : std_logic;
signal \N__62982\ : std_logic;
signal \N__62981\ : std_logic;
signal \N__62980\ : std_logic;
signal \N__62977\ : std_logic;
signal \N__62974\ : std_logic;
signal \N__62971\ : std_logic;
signal \N__62968\ : std_logic;
signal \N__62965\ : std_logic;
signal \N__62962\ : std_logic;
signal \N__62959\ : std_logic;
signal \N__62956\ : std_logic;
signal \N__62953\ : std_logic;
signal \N__62948\ : std_logic;
signal \N__62943\ : std_logic;
signal \N__62940\ : std_logic;
signal \N__62939\ : std_logic;
signal \N__62934\ : std_logic;
signal \N__62931\ : std_logic;
signal \N__62928\ : std_logic;
signal \N__62927\ : std_logic;
signal \N__62924\ : std_logic;
signal \N__62921\ : std_logic;
signal \N__62920\ : std_logic;
signal \N__62919\ : std_logic;
signal \N__62916\ : std_logic;
signal \N__62911\ : std_logic;
signal \N__62908\ : std_logic;
signal \N__62905\ : std_logic;
signal \N__62900\ : std_logic;
signal \N__62895\ : std_logic;
signal \N__62894\ : std_logic;
signal \N__62891\ : std_logic;
signal \N__62888\ : std_logic;
signal \N__62887\ : std_logic;
signal \N__62886\ : std_logic;
signal \N__62881\ : std_logic;
signal \N__62876\ : std_logic;
signal \N__62875\ : std_logic;
signal \N__62872\ : std_logic;
signal \N__62869\ : std_logic;
signal \N__62866\ : std_logic;
signal \N__62859\ : std_logic;
signal \N__62858\ : std_logic;
signal \N__62855\ : std_logic;
signal \N__62854\ : std_logic;
signal \N__62849\ : std_logic;
signal \N__62848\ : std_logic;
signal \N__62847\ : std_logic;
signal \N__62844\ : std_logic;
signal \N__62841\ : std_logic;
signal \N__62838\ : std_logic;
signal \N__62835\ : std_logic;
signal \N__62832\ : std_logic;
signal \N__62829\ : std_logic;
signal \N__62826\ : std_logic;
signal \N__62823\ : std_logic;
signal \N__62820\ : std_logic;
signal \N__62815\ : std_logic;
signal \N__62808\ : std_logic;
signal \N__62807\ : std_logic;
signal \N__62806\ : std_logic;
signal \N__62803\ : std_logic;
signal \N__62800\ : std_logic;
signal \N__62799\ : std_logic;
signal \N__62796\ : std_logic;
signal \N__62795\ : std_logic;
signal \N__62792\ : std_logic;
signal \N__62787\ : std_logic;
signal \N__62784\ : std_logic;
signal \N__62781\ : std_logic;
signal \N__62774\ : std_logic;
signal \N__62769\ : std_logic;
signal \N__62768\ : std_logic;
signal \N__62767\ : std_logic;
signal \N__62766\ : std_logic;
signal \N__62759\ : std_logic;
signal \N__62758\ : std_logic;
signal \N__62757\ : std_logic;
signal \N__62756\ : std_logic;
signal \N__62753\ : std_logic;
signal \N__62750\ : std_logic;
signal \N__62743\ : std_logic;
signal \N__62742\ : std_logic;
signal \N__62735\ : std_logic;
signal \N__62732\ : std_logic;
signal \N__62727\ : std_logic;
signal \N__62724\ : std_logic;
signal \N__62721\ : std_logic;
signal \N__62720\ : std_logic;
signal \N__62715\ : std_logic;
signal \N__62712\ : std_logic;
signal \N__62711\ : std_logic;
signal \N__62710\ : std_logic;
signal \N__62705\ : std_logic;
signal \N__62702\ : std_logic;
signal \N__62699\ : std_logic;
signal \N__62696\ : std_logic;
signal \N__62693\ : std_logic;
signal \N__62688\ : std_logic;
signal \N__62687\ : std_logic;
signal \N__62686\ : std_logic;
signal \N__62683\ : std_logic;
signal \N__62682\ : std_logic;
signal \N__62677\ : std_logic;
signal \N__62674\ : std_logic;
signal \N__62671\ : std_logic;
signal \N__62668\ : std_logic;
signal \N__62667\ : std_logic;
signal \N__62666\ : std_logic;
signal \N__62663\ : std_logic;
signal \N__62658\ : std_logic;
signal \N__62655\ : std_logic;
signal \N__62652\ : std_logic;
signal \N__62643\ : std_logic;
signal \N__62640\ : std_logic;
signal \N__62639\ : std_logic;
signal \N__62638\ : std_logic;
signal \N__62635\ : std_logic;
signal \N__62632\ : std_logic;
signal \N__62629\ : std_logic;
signal \N__62624\ : std_logic;
signal \N__62621\ : std_logic;
signal \N__62616\ : std_logic;
signal \N__62615\ : std_logic;
signal \N__62614\ : std_logic;
signal \N__62613\ : std_logic;
signal \N__62610\ : std_logic;
signal \N__62607\ : std_logic;
signal \N__62604\ : std_logic;
signal \N__62603\ : std_logic;
signal \N__62598\ : std_logic;
signal \N__62595\ : std_logic;
signal \N__62592\ : std_logic;
signal \N__62591\ : std_logic;
signal \N__62588\ : std_logic;
signal \N__62585\ : std_logic;
signal \N__62582\ : std_logic;
signal \N__62579\ : std_logic;
signal \N__62574\ : std_logic;
signal \N__62571\ : std_logic;
signal \N__62566\ : std_logic;
signal \N__62559\ : std_logic;
signal \N__62556\ : std_logic;
signal \N__62553\ : std_logic;
signal \N__62550\ : std_logic;
signal \N__62549\ : std_logic;
signal \N__62546\ : std_logic;
signal \N__62543\ : std_logic;
signal \N__62538\ : std_logic;
signal \N__62535\ : std_logic;
signal \N__62532\ : std_logic;
signal \N__62529\ : std_logic;
signal \N__62528\ : std_logic;
signal \N__62527\ : std_logic;
signal \N__62526\ : std_logic;
signal \N__62523\ : std_logic;
signal \N__62518\ : std_logic;
signal \N__62515\ : std_logic;
signal \N__62512\ : std_logic;
signal \N__62509\ : std_logic;
signal \N__62506\ : std_logic;
signal \N__62503\ : std_logic;
signal \N__62500\ : std_logic;
signal \N__62493\ : std_logic;
signal \N__62490\ : std_logic;
signal \N__62487\ : std_logic;
signal \N__62484\ : std_logic;
signal \N__62483\ : std_logic;
signal \N__62480\ : std_logic;
signal \N__62477\ : std_logic;
signal \N__62476\ : std_logic;
signal \N__62471\ : std_logic;
signal \N__62468\ : std_logic;
signal \N__62463\ : std_logic;
signal \N__62460\ : std_logic;
signal \N__62459\ : std_logic;
signal \N__62458\ : std_logic;
signal \N__62455\ : std_logic;
signal \N__62452\ : std_logic;
signal \N__62449\ : std_logic;
signal \N__62446\ : std_logic;
signal \N__62445\ : std_logic;
signal \N__62442\ : std_logic;
signal \N__62439\ : std_logic;
signal \N__62436\ : std_logic;
signal \N__62433\ : std_logic;
signal \N__62424\ : std_logic;
signal \N__62423\ : std_logic;
signal \N__62420\ : std_logic;
signal \N__62417\ : std_logic;
signal \N__62412\ : std_logic;
signal \N__62411\ : std_logic;
signal \N__62408\ : std_logic;
signal \N__62407\ : std_logic;
signal \N__62404\ : std_logic;
signal \N__62401\ : std_logic;
signal \N__62398\ : std_logic;
signal \N__62397\ : std_logic;
signal \N__62396\ : std_logic;
signal \N__62389\ : std_logic;
signal \N__62386\ : std_logic;
signal \N__62383\ : std_logic;
signal \N__62380\ : std_logic;
signal \N__62379\ : std_logic;
signal \N__62376\ : std_logic;
signal \N__62371\ : std_logic;
signal \N__62368\ : std_logic;
signal \N__62361\ : std_logic;
signal \N__62360\ : std_logic;
signal \N__62357\ : std_logic;
signal \N__62356\ : std_logic;
signal \N__62355\ : std_logic;
signal \N__62354\ : std_logic;
signal \N__62353\ : std_logic;
signal \N__62350\ : std_logic;
signal \N__62345\ : std_logic;
signal \N__62338\ : std_logic;
signal \N__62331\ : std_logic;
signal \N__62328\ : std_logic;
signal \N__62325\ : std_logic;
signal \N__62322\ : std_logic;
signal \N__62319\ : std_logic;
signal \N__62318\ : std_logic;
signal \N__62317\ : std_logic;
signal \N__62316\ : std_logic;
signal \N__62313\ : std_logic;
signal \N__62310\ : std_logic;
signal \N__62309\ : std_logic;
signal \N__62306\ : std_logic;
signal \N__62303\ : std_logic;
signal \N__62300\ : std_logic;
signal \N__62297\ : std_logic;
signal \N__62296\ : std_logic;
signal \N__62295\ : std_logic;
signal \N__62294\ : std_logic;
signal \N__62291\ : std_logic;
signal \N__62286\ : std_logic;
signal \N__62281\ : std_logic;
signal \N__62278\ : std_logic;
signal \N__62275\ : std_logic;
signal \N__62272\ : std_logic;
signal \N__62271\ : std_logic;
signal \N__62268\ : std_logic;
signal \N__62265\ : std_logic;
signal \N__62262\ : std_logic;
signal \N__62259\ : std_logic;
signal \N__62254\ : std_logic;
signal \N__62253\ : std_logic;
signal \N__62250\ : std_logic;
signal \N__62245\ : std_logic;
signal \N__62244\ : std_logic;
signal \N__62241\ : std_logic;
signal \N__62236\ : std_logic;
signal \N__62233\ : std_logic;
signal \N__62228\ : std_logic;
signal \N__62225\ : std_logic;
signal \N__62222\ : std_logic;
signal \N__62219\ : std_logic;
signal \N__62216\ : std_logic;
signal \N__62213\ : std_logic;
signal \N__62210\ : std_logic;
signal \N__62207\ : std_logic;
signal \N__62204\ : std_logic;
signal \N__62201\ : std_logic;
signal \N__62198\ : std_logic;
signal \N__62197\ : std_logic;
signal \N__62194\ : std_logic;
signal \N__62191\ : std_logic;
signal \N__62188\ : std_logic;
signal \N__62185\ : std_logic;
signal \N__62182\ : std_logic;
signal \N__62179\ : std_logic;
signal \N__62166\ : std_logic;
signal \N__62163\ : std_logic;
signal \N__62160\ : std_logic;
signal \N__62157\ : std_logic;
signal \N__62154\ : std_logic;
signal \N__62151\ : std_logic;
signal \N__62148\ : std_logic;
signal \N__62145\ : std_logic;
signal \N__62142\ : std_logic;
signal \N__62141\ : std_logic;
signal \N__62136\ : std_logic;
signal \N__62133\ : std_logic;
signal \N__62132\ : std_logic;
signal \N__62127\ : std_logic;
signal \N__62124\ : std_logic;
signal \N__62123\ : std_logic;
signal \N__62120\ : std_logic;
signal \N__62119\ : std_logic;
signal \N__62116\ : std_logic;
signal \N__62113\ : std_logic;
signal \N__62110\ : std_logic;
signal \N__62107\ : std_logic;
signal \N__62102\ : std_logic;
signal \N__62099\ : std_logic;
signal \N__62096\ : std_logic;
signal \N__62091\ : std_logic;
signal \N__62088\ : std_logic;
signal \N__62085\ : std_logic;
signal \N__62084\ : std_logic;
signal \N__62081\ : std_logic;
signal \N__62078\ : std_logic;
signal \N__62075\ : std_logic;
signal \N__62072\ : std_logic;
signal \N__62071\ : std_logic;
signal \N__62070\ : std_logic;
signal \N__62069\ : std_logic;
signal \N__62064\ : std_logic;
signal \N__62057\ : std_logic;
signal \N__62052\ : std_logic;
signal \N__62049\ : std_logic;
signal \N__62046\ : std_logic;
signal \N__62043\ : std_logic;
signal \N__62040\ : std_logic;
signal \N__62037\ : std_logic;
signal \N__62034\ : std_logic;
signal \N__62033\ : std_logic;
signal \N__62030\ : std_logic;
signal \N__62027\ : std_logic;
signal \N__62022\ : std_logic;
signal \N__62019\ : std_logic;
signal \N__62016\ : std_logic;
signal \N__62013\ : std_logic;
signal \N__62010\ : std_logic;
signal \N__62009\ : std_logic;
signal \N__62006\ : std_logic;
signal \N__62003\ : std_logic;
signal \N__62000\ : std_logic;
signal \N__61995\ : std_logic;
signal \N__61992\ : std_logic;
signal \N__61991\ : std_logic;
signal \N__61988\ : std_logic;
signal \N__61987\ : std_logic;
signal \N__61984\ : std_logic;
signal \N__61981\ : std_logic;
signal \N__61978\ : std_logic;
signal \N__61975\ : std_logic;
signal \N__61972\ : std_logic;
signal \N__61969\ : std_logic;
signal \N__61962\ : std_logic;
signal \N__61959\ : std_logic;
signal \N__61956\ : std_logic;
signal \N__61953\ : std_logic;
signal \N__61950\ : std_logic;
signal \N__61949\ : std_logic;
signal \N__61946\ : std_logic;
signal \N__61943\ : std_logic;
signal \N__61938\ : std_logic;
signal \N__61935\ : std_logic;
signal \N__61934\ : std_logic;
signal \N__61931\ : std_logic;
signal \N__61928\ : std_logic;
signal \N__61927\ : std_logic;
signal \N__61926\ : std_logic;
signal \N__61921\ : std_logic;
signal \N__61916\ : std_logic;
signal \N__61913\ : std_logic;
signal \N__61910\ : std_logic;
signal \N__61905\ : std_logic;
signal \N__61902\ : std_logic;
signal \N__61901\ : std_logic;
signal \N__61898\ : std_logic;
signal \N__61897\ : std_logic;
signal \N__61894\ : std_logic;
signal \N__61891\ : std_logic;
signal \N__61890\ : std_logic;
signal \N__61887\ : std_logic;
signal \N__61884\ : std_logic;
signal \N__61881\ : std_logic;
signal \N__61878\ : std_logic;
signal \N__61875\ : std_logic;
signal \N__61872\ : std_logic;
signal \N__61867\ : std_logic;
signal \N__61860\ : std_logic;
signal \N__61859\ : std_logic;
signal \N__61856\ : std_logic;
signal \N__61853\ : std_logic;
signal \N__61852\ : std_logic;
signal \N__61851\ : std_logic;
signal \N__61846\ : std_logic;
signal \N__61841\ : std_logic;
signal \N__61838\ : std_logic;
signal \N__61833\ : std_logic;
signal \N__61830\ : std_logic;
signal \N__61827\ : std_logic;
signal \N__61824\ : std_logic;
signal \N__61821\ : std_logic;
signal \N__61818\ : std_logic;
signal \N__61815\ : std_logic;
signal \N__61812\ : std_logic;
signal \N__61811\ : std_logic;
signal \N__61808\ : std_logic;
signal \N__61805\ : std_logic;
signal \N__61800\ : std_logic;
signal \N__61797\ : std_logic;
signal \N__61796\ : std_logic;
signal \N__61793\ : std_logic;
signal \N__61792\ : std_logic;
signal \N__61789\ : std_logic;
signal \N__61786\ : std_logic;
signal \N__61783\ : std_logic;
signal \N__61782\ : std_logic;
signal \N__61781\ : std_logic;
signal \N__61774\ : std_logic;
signal \N__61771\ : std_logic;
signal \N__61768\ : std_logic;
signal \N__61767\ : std_logic;
signal \N__61762\ : std_logic;
signal \N__61759\ : std_logic;
signal \N__61756\ : std_logic;
signal \N__61753\ : std_logic;
signal \N__61746\ : std_logic;
signal \N__61745\ : std_logic;
signal \N__61742\ : std_logic;
signal \N__61741\ : std_logic;
signal \N__61740\ : std_logic;
signal \N__61739\ : std_logic;
signal \N__61738\ : std_logic;
signal \N__61735\ : std_logic;
signal \N__61732\ : std_logic;
signal \N__61725\ : std_logic;
signal \N__61720\ : std_logic;
signal \N__61719\ : std_logic;
signal \N__61716\ : std_logic;
signal \N__61711\ : std_logic;
signal \N__61708\ : std_logic;
signal \N__61703\ : std_logic;
signal \N__61698\ : std_logic;
signal \N__61695\ : std_logic;
signal \N__61692\ : std_logic;
signal \N__61691\ : std_logic;
signal \N__61688\ : std_logic;
signal \N__61685\ : std_logic;
signal \N__61680\ : std_logic;
signal \N__61677\ : std_logic;
signal \N__61674\ : std_logic;
signal \N__61671\ : std_logic;
signal \N__61668\ : std_logic;
signal \N__61665\ : std_logic;
signal \N__61662\ : std_logic;
signal \N__61659\ : std_logic;
signal \N__61658\ : std_logic;
signal \N__61655\ : std_logic;
signal \N__61652\ : std_logic;
signal \N__61649\ : std_logic;
signal \N__61648\ : std_logic;
signal \N__61645\ : std_logic;
signal \N__61642\ : std_logic;
signal \N__61639\ : std_logic;
signal \N__61634\ : std_logic;
signal \N__61629\ : std_logic;
signal \N__61626\ : std_logic;
signal \N__61623\ : std_logic;
signal \N__61620\ : std_logic;
signal \N__61617\ : std_logic;
signal \N__61616\ : std_logic;
signal \N__61613\ : std_logic;
signal \N__61610\ : std_logic;
signal \N__61607\ : std_logic;
signal \N__61604\ : std_logic;
signal \N__61601\ : std_logic;
signal \N__61596\ : std_logic;
signal \N__61593\ : std_logic;
signal \N__61590\ : std_logic;
signal \N__61589\ : std_logic;
signal \N__61586\ : std_logic;
signal \N__61583\ : std_logic;
signal \N__61582\ : std_logic;
signal \N__61579\ : std_logic;
signal \N__61576\ : std_logic;
signal \N__61573\ : std_logic;
signal \N__61570\ : std_logic;
signal \N__61567\ : std_logic;
signal \N__61560\ : std_logic;
signal \N__61557\ : std_logic;
signal \N__61554\ : std_logic;
signal \N__61553\ : std_logic;
signal \N__61552\ : std_logic;
signal \N__61549\ : std_logic;
signal \N__61548\ : std_logic;
signal \N__61545\ : std_logic;
signal \N__61542\ : std_logic;
signal \N__61541\ : std_logic;
signal \N__61538\ : std_logic;
signal \N__61535\ : std_logic;
signal \N__61530\ : std_logic;
signal \N__61527\ : std_logic;
signal \N__61524\ : std_logic;
signal \N__61521\ : std_logic;
signal \N__61518\ : std_logic;
signal \N__61515\ : std_logic;
signal \N__61512\ : std_logic;
signal \N__61503\ : std_logic;
signal \N__61500\ : std_logic;
signal \N__61497\ : std_logic;
signal \N__61494\ : std_logic;
signal \N__61491\ : std_logic;
signal \N__61488\ : std_logic;
signal \N__61487\ : std_logic;
signal \N__61482\ : std_logic;
signal \N__61479\ : std_logic;
signal \N__61476\ : std_logic;
signal \N__61475\ : std_logic;
signal \N__61470\ : std_logic;
signal \N__61467\ : std_logic;
signal \N__61466\ : std_logic;
signal \N__61463\ : std_logic;
signal \N__61460\ : std_logic;
signal \N__61457\ : std_logic;
signal \N__61454\ : std_logic;
signal \N__61451\ : std_logic;
signal \N__61448\ : std_logic;
signal \N__61443\ : std_logic;
signal \N__61440\ : std_logic;
signal \N__61437\ : std_logic;
signal \N__61434\ : std_logic;
signal \N__61433\ : std_logic;
signal \N__61430\ : std_logic;
signal \N__61429\ : std_logic;
signal \N__61426\ : std_logic;
signal \N__61425\ : std_logic;
signal \N__61424\ : std_logic;
signal \N__61421\ : std_logic;
signal \N__61418\ : std_logic;
signal \N__61415\ : std_logic;
signal \N__61412\ : std_logic;
signal \N__61409\ : std_logic;
signal \N__61404\ : std_logic;
signal \N__61399\ : std_logic;
signal \N__61392\ : std_logic;
signal \N__61391\ : std_logic;
signal \N__61388\ : std_logic;
signal \N__61385\ : std_logic;
signal \N__61384\ : std_logic;
signal \N__61381\ : std_logic;
signal \N__61380\ : std_logic;
signal \N__61377\ : std_logic;
signal \N__61374\ : std_logic;
signal \N__61371\ : std_logic;
signal \N__61368\ : std_logic;
signal \N__61363\ : std_logic;
signal \N__61360\ : std_logic;
signal \N__61357\ : std_logic;
signal \N__61352\ : std_logic;
signal \N__61347\ : std_logic;
signal \N__61344\ : std_logic;
signal \N__61341\ : std_logic;
signal \N__61338\ : std_logic;
signal \N__61335\ : std_logic;
signal \N__61334\ : std_logic;
signal \N__61333\ : std_logic;
signal \N__61330\ : std_logic;
signal \N__61327\ : std_logic;
signal \N__61324\ : std_logic;
signal \N__61321\ : std_logic;
signal \N__61316\ : std_logic;
signal \N__61313\ : std_logic;
signal \N__61310\ : std_logic;
signal \N__61305\ : std_logic;
signal \N__61302\ : std_logic;
signal \N__61299\ : std_logic;
signal \N__61298\ : std_logic;
signal \N__61295\ : std_logic;
signal \N__61294\ : std_logic;
signal \N__61293\ : std_logic;
signal \N__61292\ : std_logic;
signal \N__61289\ : std_logic;
signal \N__61288\ : std_logic;
signal \N__61285\ : std_logic;
signal \N__61282\ : std_logic;
signal \N__61277\ : std_logic;
signal \N__61272\ : std_logic;
signal \N__61263\ : std_logic;
signal \N__61262\ : std_logic;
signal \N__61259\ : std_logic;
signal \N__61256\ : std_logic;
signal \N__61255\ : std_logic;
signal \N__61252\ : std_logic;
signal \N__61249\ : std_logic;
signal \N__61246\ : std_logic;
signal \N__61245\ : std_logic;
signal \N__61242\ : std_logic;
signal \N__61239\ : std_logic;
signal \N__61236\ : std_logic;
signal \N__61235\ : std_logic;
signal \N__61232\ : std_logic;
signal \N__61227\ : std_logic;
signal \N__61224\ : std_logic;
signal \N__61221\ : std_logic;
signal \N__61212\ : std_logic;
signal \N__61209\ : std_logic;
signal \N__61206\ : std_logic;
signal \N__61203\ : std_logic;
signal \N__61200\ : std_logic;
signal \N__61197\ : std_logic;
signal \N__61194\ : std_logic;
signal \N__61191\ : std_logic;
signal \N__61188\ : std_logic;
signal \N__61185\ : std_logic;
signal \N__61182\ : std_logic;
signal \N__61179\ : std_logic;
signal \N__61176\ : std_logic;
signal \N__61175\ : std_logic;
signal \N__61172\ : std_logic;
signal \N__61169\ : std_logic;
signal \N__61166\ : std_logic;
signal \N__61163\ : std_logic;
signal \N__61160\ : std_logic;
signal \N__61157\ : std_logic;
signal \N__61152\ : std_logic;
signal \N__61149\ : std_logic;
signal \N__61146\ : std_logic;
signal \N__61143\ : std_logic;
signal \N__61142\ : std_logic;
signal \N__61139\ : std_logic;
signal \N__61136\ : std_logic;
signal \N__61133\ : std_logic;
signal \N__61128\ : std_logic;
signal \N__61125\ : std_logic;
signal \N__61122\ : std_logic;
signal \N__61119\ : std_logic;
signal \N__61116\ : std_logic;
signal \N__61113\ : std_logic;
signal \N__61112\ : std_logic;
signal \N__61111\ : std_logic;
signal \N__61104\ : std_logic;
signal \N__61101\ : std_logic;
signal \N__61098\ : std_logic;
signal \N__61095\ : std_logic;
signal \N__61094\ : std_logic;
signal \N__61091\ : std_logic;
signal \N__61088\ : std_logic;
signal \N__61083\ : std_logic;
signal \N__61080\ : std_logic;
signal \N__61077\ : std_logic;
signal \N__61074\ : std_logic;
signal \N__61071\ : std_logic;
signal \N__61068\ : std_logic;
signal \N__61065\ : std_logic;
signal \N__61064\ : std_logic;
signal \N__61061\ : std_logic;
signal \N__61058\ : std_logic;
signal \N__61057\ : std_logic;
signal \N__61054\ : std_logic;
signal \N__61051\ : std_logic;
signal \N__61048\ : std_logic;
signal \N__61045\ : std_logic;
signal \N__61044\ : std_logic;
signal \N__61043\ : std_logic;
signal \N__61040\ : std_logic;
signal \N__61037\ : std_logic;
signal \N__61036\ : std_logic;
signal \N__61035\ : std_logic;
signal \N__61032\ : std_logic;
signal \N__61031\ : std_logic;
signal \N__61030\ : std_logic;
signal \N__61025\ : std_logic;
signal \N__61020\ : std_logic;
signal \N__61017\ : std_logic;
signal \N__61014\ : std_logic;
signal \N__61011\ : std_logic;
signal \N__61008\ : std_logic;
signal \N__61005\ : std_logic;
signal \N__60998\ : std_logic;
signal \N__60987\ : std_logic;
signal \N__60984\ : std_logic;
signal \N__60981\ : std_logic;
signal \N__60978\ : std_logic;
signal \N__60975\ : std_logic;
signal \N__60972\ : std_logic;
signal \N__60969\ : std_logic;
signal \N__60966\ : std_logic;
signal \N__60963\ : std_logic;
signal \N__60960\ : std_logic;
signal \N__60957\ : std_logic;
signal \N__60954\ : std_logic;
signal \N__60953\ : std_logic;
signal \N__60952\ : std_logic;
signal \N__60949\ : std_logic;
signal \N__60946\ : std_logic;
signal \N__60943\ : std_logic;
signal \N__60942\ : std_logic;
signal \N__60939\ : std_logic;
signal \N__60934\ : std_logic;
signal \N__60931\ : std_logic;
signal \N__60924\ : std_logic;
signal \N__60921\ : std_logic;
signal \N__60918\ : std_logic;
signal \N__60915\ : std_logic;
signal \N__60912\ : std_logic;
signal \N__60909\ : std_logic;
signal \N__60906\ : std_logic;
signal \N__60905\ : std_logic;
signal \N__60900\ : std_logic;
signal \N__60899\ : std_logic;
signal \N__60896\ : std_logic;
signal \N__60895\ : std_logic;
signal \N__60892\ : std_logic;
signal \N__60891\ : std_logic;
signal \N__60888\ : std_logic;
signal \N__60885\ : std_logic;
signal \N__60884\ : std_logic;
signal \N__60883\ : std_logic;
signal \N__60882\ : std_logic;
signal \N__60877\ : std_logic;
signal \N__60874\ : std_logic;
signal \N__60867\ : std_logic;
signal \N__60864\ : std_logic;
signal \N__60855\ : std_logic;
signal \N__60854\ : std_logic;
signal \N__60851\ : std_logic;
signal \N__60850\ : std_logic;
signal \N__60847\ : std_logic;
signal \N__60844\ : std_logic;
signal \N__60841\ : std_logic;
signal \N__60836\ : std_logic;
signal \N__60835\ : std_logic;
signal \N__60834\ : std_logic;
signal \N__60829\ : std_logic;
signal \N__60824\ : std_logic;
signal \N__60819\ : std_logic;
signal \N__60818\ : std_logic;
signal \N__60817\ : std_logic;
signal \N__60814\ : std_logic;
signal \N__60809\ : std_logic;
signal \N__60806\ : std_logic;
signal \N__60803\ : std_logic;
signal \N__60798\ : std_logic;
signal \N__60797\ : std_logic;
signal \N__60796\ : std_logic;
signal \N__60793\ : std_logic;
signal \N__60792\ : std_logic;
signal \N__60789\ : std_logic;
signal \N__60786\ : std_logic;
signal \N__60783\ : std_logic;
signal \N__60780\ : std_logic;
signal \N__60775\ : std_logic;
signal \N__60774\ : std_logic;
signal \N__60773\ : std_logic;
signal \N__60770\ : std_logic;
signal \N__60765\ : std_logic;
signal \N__60760\ : std_logic;
signal \N__60753\ : std_logic;
signal \N__60750\ : std_logic;
signal \N__60747\ : std_logic;
signal \N__60746\ : std_logic;
signal \N__60743\ : std_logic;
signal \N__60742\ : std_logic;
signal \N__60741\ : std_logic;
signal \N__60738\ : std_logic;
signal \N__60737\ : std_logic;
signal \N__60734\ : std_logic;
signal \N__60731\ : std_logic;
signal \N__60728\ : std_logic;
signal \N__60723\ : std_logic;
signal \N__60714\ : std_logic;
signal \N__60711\ : std_logic;
signal \N__60708\ : std_logic;
signal \N__60705\ : std_logic;
signal \N__60702\ : std_logic;
signal \N__60699\ : std_logic;
signal \N__60696\ : std_logic;
signal \N__60693\ : std_logic;
signal \N__60690\ : std_logic;
signal \N__60687\ : std_logic;
signal \N__60686\ : std_logic;
signal \N__60683\ : std_logic;
signal \N__60680\ : std_logic;
signal \N__60677\ : std_logic;
signal \N__60674\ : std_logic;
signal \N__60671\ : std_logic;
signal \N__60666\ : std_logic;
signal \N__60663\ : std_logic;
signal \N__60660\ : std_logic;
signal \N__60657\ : std_logic;
signal \N__60654\ : std_logic;
signal \N__60651\ : std_logic;
signal \N__60648\ : std_logic;
signal \N__60645\ : std_logic;
signal \N__60644\ : std_logic;
signal \N__60641\ : std_logic;
signal \N__60638\ : std_logic;
signal \N__60637\ : std_logic;
signal \N__60636\ : std_logic;
signal \N__60635\ : std_logic;
signal \N__60634\ : std_logic;
signal \N__60633\ : std_logic;
signal \N__60632\ : std_logic;
signal \N__60631\ : std_logic;
signal \N__60628\ : std_logic;
signal \N__60625\ : std_logic;
signal \N__60620\ : std_logic;
signal \N__60617\ : std_logic;
signal \N__60610\ : std_logic;
signal \N__60607\ : std_logic;
signal \N__60594\ : std_logic;
signal \N__60591\ : std_logic;
signal \N__60588\ : std_logic;
signal \N__60585\ : std_logic;
signal \N__60582\ : std_logic;
signal \N__60579\ : std_logic;
signal \N__60576\ : std_logic;
signal \N__60573\ : std_logic;
signal \N__60570\ : std_logic;
signal \N__60567\ : std_logic;
signal \N__60566\ : std_logic;
signal \N__60563\ : std_logic;
signal \N__60562\ : std_logic;
signal \N__60559\ : std_logic;
signal \N__60558\ : std_logic;
signal \N__60557\ : std_logic;
signal \N__60554\ : std_logic;
signal \N__60553\ : std_logic;
signal \N__60552\ : std_logic;
signal \N__60549\ : std_logic;
signal \N__60548\ : std_logic;
signal \N__60547\ : std_logic;
signal \N__60546\ : std_logic;
signal \N__60545\ : std_logic;
signal \N__60542\ : std_logic;
signal \N__60537\ : std_logic;
signal \N__60536\ : std_logic;
signal \N__60535\ : std_logic;
signal \N__60534\ : std_logic;
signal \N__60533\ : std_logic;
signal \N__60530\ : std_logic;
signal \N__60527\ : std_logic;
signal \N__60524\ : std_logic;
signal \N__60521\ : std_logic;
signal \N__60518\ : std_logic;
signal \N__60515\ : std_logic;
signal \N__60512\ : std_logic;
signal \N__60511\ : std_logic;
signal \N__60508\ : std_logic;
signal \N__60507\ : std_logic;
signal \N__60504\ : std_logic;
signal \N__60501\ : std_logic;
signal \N__60494\ : std_logic;
signal \N__60491\ : std_logic;
signal \N__60490\ : std_logic;
signal \N__60481\ : std_logic;
signal \N__60478\ : std_logic;
signal \N__60475\ : std_logic;
signal \N__60470\ : std_logic;
signal \N__60465\ : std_logic;
signal \N__60458\ : std_logic;
signal \N__60453\ : std_logic;
signal \N__60438\ : std_logic;
signal \N__60435\ : std_logic;
signal \N__60432\ : std_logic;
signal \N__60431\ : std_logic;
signal \N__60428\ : std_logic;
signal \N__60427\ : std_logic;
signal \N__60424\ : std_logic;
signal \N__60421\ : std_logic;
signal \N__60418\ : std_logic;
signal \N__60417\ : std_logic;
signal \N__60416\ : std_logic;
signal \N__60415\ : std_logic;
signal \N__60414\ : std_logic;
signal \N__60413\ : std_logic;
signal \N__60410\ : std_logic;
signal \N__60409\ : std_logic;
signal \N__60408\ : std_logic;
signal \N__60405\ : std_logic;
signal \N__60394\ : std_logic;
signal \N__60391\ : std_logic;
signal \N__60388\ : std_logic;
signal \N__60387\ : std_logic;
signal \N__60386\ : std_logic;
signal \N__60385\ : std_logic;
signal \N__60382\ : std_logic;
signal \N__60379\ : std_logic;
signal \N__60378\ : std_logic;
signal \N__60377\ : std_logic;
signal \N__60372\ : std_logic;
signal \N__60369\ : std_logic;
signal \N__60366\ : std_logic;
signal \N__60363\ : std_logic;
signal \N__60360\ : std_logic;
signal \N__60357\ : std_logic;
signal \N__60354\ : std_logic;
signal \N__60347\ : std_logic;
signal \N__60342\ : std_logic;
signal \N__60327\ : std_logic;
signal \N__60324\ : std_logic;
signal \N__60321\ : std_logic;
signal \N__60318\ : std_logic;
signal \N__60315\ : std_logic;
signal \N__60312\ : std_logic;
signal \N__60309\ : std_logic;
signal \N__60306\ : std_logic;
signal \N__60305\ : std_logic;
signal \N__60304\ : std_logic;
signal \N__60303\ : std_logic;
signal \N__60302\ : std_logic;
signal \N__60301\ : std_logic;
signal \N__60298\ : std_logic;
signal \N__60297\ : std_logic;
signal \N__60296\ : std_logic;
signal \N__60295\ : std_logic;
signal \N__60292\ : std_logic;
signal \N__60289\ : std_logic;
signal \N__60284\ : std_logic;
signal \N__60283\ : std_logic;
signal \N__60280\ : std_logic;
signal \N__60277\ : std_logic;
signal \N__60274\ : std_logic;
signal \N__60269\ : std_logic;
signal \N__60266\ : std_logic;
signal \N__60261\ : std_logic;
signal \N__60258\ : std_logic;
signal \N__60243\ : std_logic;
signal \N__60240\ : std_logic;
signal \N__60239\ : std_logic;
signal \N__60236\ : std_logic;
signal \N__60235\ : std_logic;
signal \N__60234\ : std_logic;
signal \N__60231\ : std_logic;
signal \N__60230\ : std_logic;
signal \N__60229\ : std_logic;
signal \N__60228\ : std_logic;
signal \N__60227\ : std_logic;
signal \N__60224\ : std_logic;
signal \N__60219\ : std_logic;
signal \N__60212\ : std_logic;
signal \N__60209\ : std_logic;
signal \N__60208\ : std_logic;
signal \N__60205\ : std_logic;
signal \N__60204\ : std_logic;
signal \N__60203\ : std_logic;
signal \N__60198\ : std_logic;
signal \N__60195\ : std_logic;
signal \N__60188\ : std_logic;
signal \N__60187\ : std_logic;
signal \N__60186\ : std_logic;
signal \N__60183\ : std_logic;
signal \N__60180\ : std_logic;
signal \N__60173\ : std_logic;
signal \N__60168\ : std_logic;
signal \N__60159\ : std_logic;
signal \N__60156\ : std_logic;
signal \N__60155\ : std_logic;
signal \N__60152\ : std_logic;
signal \N__60149\ : std_logic;
signal \N__60148\ : std_logic;
signal \N__60143\ : std_logic;
signal \N__60140\ : std_logic;
signal \N__60135\ : std_logic;
signal \N__60132\ : std_logic;
signal \N__60131\ : std_logic;
signal \N__60128\ : std_logic;
signal \N__60125\ : std_logic;
signal \N__60120\ : std_logic;
signal \N__60117\ : std_logic;
signal \N__60116\ : std_logic;
signal \N__60113\ : std_logic;
signal \N__60110\ : std_logic;
signal \N__60107\ : std_logic;
signal \N__60102\ : std_logic;
signal \N__60099\ : std_logic;
signal \N__60096\ : std_logic;
signal \N__60093\ : std_logic;
signal \N__60090\ : std_logic;
signal \N__60087\ : std_logic;
signal \N__60084\ : std_logic;
signal \N__60081\ : std_logic;
signal \N__60080\ : std_logic;
signal \N__60077\ : std_logic;
signal \N__60074\ : std_logic;
signal \N__60071\ : std_logic;
signal \N__60068\ : std_logic;
signal \N__60063\ : std_logic;
signal \N__60062\ : std_logic;
signal \N__60061\ : std_logic;
signal \N__60060\ : std_logic;
signal \N__60057\ : std_logic;
signal \N__60054\ : std_logic;
signal \N__60049\ : std_logic;
signal \N__60048\ : std_logic;
signal \N__60045\ : std_logic;
signal \N__60040\ : std_logic;
signal \N__60037\ : std_logic;
signal \N__60030\ : std_logic;
signal \N__60029\ : std_logic;
signal \N__60026\ : std_logic;
signal \N__60023\ : std_logic;
signal \N__60020\ : std_logic;
signal \N__60017\ : std_logic;
signal \N__60012\ : std_logic;
signal \N__60009\ : std_logic;
signal \N__60006\ : std_logic;
signal \N__60003\ : std_logic;
signal \N__60000\ : std_logic;
signal \N__59997\ : std_logic;
signal \N__59994\ : std_logic;
signal \N__59991\ : std_logic;
signal \N__59988\ : std_logic;
signal \N__59985\ : std_logic;
signal \N__59982\ : std_logic;
signal \N__59979\ : std_logic;
signal \N__59976\ : std_logic;
signal \N__59973\ : std_logic;
signal \N__59970\ : std_logic;
signal \N__59967\ : std_logic;
signal \N__59964\ : std_logic;
signal \N__59961\ : std_logic;
signal \N__59958\ : std_logic;
signal \N__59955\ : std_logic;
signal \N__59952\ : std_logic;
signal \N__59949\ : std_logic;
signal \N__59946\ : std_logic;
signal \N__59943\ : std_logic;
signal \N__59940\ : std_logic;
signal \N__59937\ : std_logic;
signal \N__59934\ : std_logic;
signal \N__59931\ : std_logic;
signal \N__59928\ : std_logic;
signal \N__59925\ : std_logic;
signal \N__59922\ : std_logic;
signal \N__59919\ : std_logic;
signal \N__59916\ : std_logic;
signal \N__59913\ : std_logic;
signal \N__59912\ : std_logic;
signal \N__59909\ : std_logic;
signal \N__59906\ : std_logic;
signal \N__59901\ : std_logic;
signal \N__59898\ : std_logic;
signal \N__59897\ : std_logic;
signal \N__59896\ : std_logic;
signal \N__59893\ : std_logic;
signal \N__59890\ : std_logic;
signal \N__59887\ : std_logic;
signal \N__59880\ : std_logic;
signal \N__59877\ : std_logic;
signal \N__59876\ : std_logic;
signal \N__59875\ : std_logic;
signal \N__59872\ : std_logic;
signal \N__59869\ : std_logic;
signal \N__59868\ : std_logic;
signal \N__59867\ : std_logic;
signal \N__59864\ : std_logic;
signal \N__59861\ : std_logic;
signal \N__59858\ : std_logic;
signal \N__59853\ : std_logic;
signal \N__59850\ : std_logic;
signal \N__59845\ : std_logic;
signal \N__59838\ : std_logic;
signal \N__59835\ : std_logic;
signal \N__59832\ : std_logic;
signal \N__59829\ : std_logic;
signal \N__59826\ : std_logic;
signal \N__59823\ : std_logic;
signal \N__59820\ : std_logic;
signal \N__59817\ : std_logic;
signal \N__59814\ : std_logic;
signal \N__59811\ : std_logic;
signal \N__59808\ : std_logic;
signal \N__59805\ : std_logic;
signal \N__59802\ : std_logic;
signal \N__59799\ : std_logic;
signal \N__59796\ : std_logic;
signal \N__59793\ : std_logic;
signal \N__59790\ : std_logic;
signal \N__59787\ : std_logic;
signal \N__59786\ : std_logic;
signal \N__59783\ : std_logic;
signal \N__59782\ : std_logic;
signal \N__59777\ : std_logic;
signal \N__59774\ : std_logic;
signal \N__59771\ : std_logic;
signal \N__59768\ : std_logic;
signal \N__59763\ : std_logic;
signal \N__59760\ : std_logic;
signal \N__59757\ : std_logic;
signal \N__59754\ : std_logic;
signal \N__59751\ : std_logic;
signal \N__59748\ : std_logic;
signal \N__59745\ : std_logic;
signal \N__59742\ : std_logic;
signal \N__59739\ : std_logic;
signal \N__59738\ : std_logic;
signal \N__59735\ : std_logic;
signal \N__59732\ : std_logic;
signal \N__59731\ : std_logic;
signal \N__59730\ : std_logic;
signal \N__59725\ : std_logic;
signal \N__59724\ : std_logic;
signal \N__59721\ : std_logic;
signal \N__59720\ : std_logic;
signal \N__59717\ : std_logic;
signal \N__59714\ : std_logic;
signal \N__59711\ : std_logic;
signal \N__59706\ : std_logic;
signal \N__59703\ : std_logic;
signal \N__59702\ : std_logic;
signal \N__59699\ : std_logic;
signal \N__59692\ : std_logic;
signal \N__59689\ : std_logic;
signal \N__59686\ : std_logic;
signal \N__59683\ : std_logic;
signal \N__59676\ : std_logic;
signal \N__59673\ : std_logic;
signal \N__59670\ : std_logic;
signal \N__59667\ : std_logic;
signal \N__59664\ : std_logic;
signal \N__59663\ : std_logic;
signal \N__59660\ : std_logic;
signal \N__59657\ : std_logic;
signal \N__59654\ : std_logic;
signal \N__59651\ : std_logic;
signal \N__59648\ : std_logic;
signal \N__59645\ : std_logic;
signal \N__59640\ : std_logic;
signal \N__59637\ : std_logic;
signal \N__59636\ : std_logic;
signal \N__59633\ : std_logic;
signal \N__59630\ : std_logic;
signal \N__59629\ : std_logic;
signal \N__59628\ : std_logic;
signal \N__59625\ : std_logic;
signal \N__59622\ : std_logic;
signal \N__59619\ : std_logic;
signal \N__59616\ : std_logic;
signal \N__59613\ : std_logic;
signal \N__59610\ : std_logic;
signal \N__59607\ : std_logic;
signal \N__59604\ : std_logic;
signal \N__59601\ : std_logic;
signal \N__59598\ : std_logic;
signal \N__59589\ : std_logic;
signal \N__59588\ : std_logic;
signal \N__59587\ : std_logic;
signal \N__59582\ : std_logic;
signal \N__59579\ : std_logic;
signal \N__59578\ : std_logic;
signal \N__59575\ : std_logic;
signal \N__59570\ : std_logic;
signal \N__59567\ : std_logic;
signal \N__59562\ : std_logic;
signal \N__59561\ : std_logic;
signal \N__59558\ : std_logic;
signal \N__59557\ : std_logic;
signal \N__59556\ : std_logic;
signal \N__59553\ : std_logic;
signal \N__59550\ : std_logic;
signal \N__59545\ : std_logic;
signal \N__59542\ : std_logic;
signal \N__59539\ : std_logic;
signal \N__59532\ : std_logic;
signal \N__59529\ : std_logic;
signal \N__59526\ : std_logic;
signal \N__59525\ : std_logic;
signal \N__59524\ : std_logic;
signal \N__59521\ : std_logic;
signal \N__59516\ : std_logic;
signal \N__59513\ : std_logic;
signal \N__59508\ : std_logic;
signal \N__59505\ : std_logic;
signal \N__59502\ : std_logic;
signal \N__59499\ : std_logic;
signal \N__59496\ : std_logic;
signal \N__59493\ : std_logic;
signal \N__59490\ : std_logic;
signal \N__59487\ : std_logic;
signal \N__59484\ : std_logic;
signal \N__59481\ : std_logic;
signal \N__59480\ : std_logic;
signal \N__59479\ : std_logic;
signal \N__59476\ : std_logic;
signal \N__59471\ : std_logic;
signal \N__59468\ : std_logic;
signal \N__59463\ : std_logic;
signal \N__59460\ : std_logic;
signal \N__59457\ : std_logic;
signal \N__59456\ : std_logic;
signal \N__59453\ : std_logic;
signal \N__59450\ : std_logic;
signal \N__59445\ : std_logic;
signal \N__59442\ : std_logic;
signal \N__59441\ : std_logic;
signal \N__59440\ : std_logic;
signal \N__59435\ : std_logic;
signal \N__59434\ : std_logic;
signal \N__59433\ : std_logic;
signal \N__59430\ : std_logic;
signal \N__59427\ : std_logic;
signal \N__59424\ : std_logic;
signal \N__59421\ : std_logic;
signal \N__59418\ : std_logic;
signal \N__59415\ : std_logic;
signal \N__59412\ : std_logic;
signal \N__59403\ : std_logic;
signal \N__59400\ : std_logic;
signal \N__59397\ : std_logic;
signal \N__59394\ : std_logic;
signal \N__59391\ : std_logic;
signal \N__59388\ : std_logic;
signal \N__59385\ : std_logic;
signal \N__59382\ : std_logic;
signal \N__59379\ : std_logic;
signal \N__59376\ : std_logic;
signal \N__59373\ : std_logic;
signal \N__59370\ : std_logic;
signal \N__59367\ : std_logic;
signal \N__59366\ : std_logic;
signal \N__59363\ : std_logic;
signal \N__59360\ : std_logic;
signal \N__59355\ : std_logic;
signal \N__59352\ : std_logic;
signal \N__59349\ : std_logic;
signal \N__59348\ : std_logic;
signal \N__59345\ : std_logic;
signal \N__59342\ : std_logic;
signal \N__59339\ : std_logic;
signal \N__59334\ : std_logic;
signal \N__59333\ : std_logic;
signal \N__59330\ : std_logic;
signal \N__59329\ : std_logic;
signal \N__59326\ : std_logic;
signal \N__59321\ : std_logic;
signal \N__59316\ : std_logic;
signal \N__59313\ : std_logic;
signal \N__59310\ : std_logic;
signal \N__59307\ : std_logic;
signal \N__59304\ : std_logic;
signal \N__59301\ : std_logic;
signal \N__59300\ : std_logic;
signal \N__59297\ : std_logic;
signal \N__59294\ : std_logic;
signal \N__59289\ : std_logic;
signal \N__59286\ : std_logic;
signal \N__59283\ : std_logic;
signal \N__59282\ : std_logic;
signal \N__59281\ : std_logic;
signal \N__59280\ : std_logic;
signal \N__59277\ : std_logic;
signal \N__59270\ : std_logic;
signal \N__59265\ : std_logic;
signal \N__59262\ : std_logic;
signal \N__59261\ : std_logic;
signal \N__59260\ : std_logic;
signal \N__59259\ : std_logic;
signal \N__59256\ : std_logic;
signal \N__59253\ : std_logic;
signal \N__59250\ : std_logic;
signal \N__59247\ : std_logic;
signal \N__59244\ : std_logic;
signal \N__59243\ : std_logic;
signal \N__59240\ : std_logic;
signal \N__59237\ : std_logic;
signal \N__59232\ : std_logic;
signal \N__59231\ : std_logic;
signal \N__59228\ : std_logic;
signal \N__59225\ : std_logic;
signal \N__59220\ : std_logic;
signal \N__59215\ : std_logic;
signal \N__59208\ : std_logic;
signal \N__59207\ : std_logic;
signal \N__59206\ : std_logic;
signal \N__59205\ : std_logic;
signal \N__59202\ : std_logic;
signal \N__59199\ : std_logic;
signal \N__59198\ : std_logic;
signal \N__59197\ : std_logic;
signal \N__59194\ : std_logic;
signal \N__59191\ : std_logic;
signal \N__59190\ : std_logic;
signal \N__59187\ : std_logic;
signal \N__59184\ : std_logic;
signal \N__59179\ : std_logic;
signal \N__59176\ : std_logic;
signal \N__59173\ : std_logic;
signal \N__59170\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59162\ : std_logic;
signal \N__59157\ : std_logic;
signal \N__59154\ : std_logic;
signal \N__59149\ : std_logic;
signal \N__59148\ : std_logic;
signal \N__59143\ : std_logic;
signal \N__59140\ : std_logic;
signal \N__59137\ : std_logic;
signal \N__59130\ : std_logic;
signal \N__59129\ : std_logic;
signal \N__59126\ : std_logic;
signal \N__59125\ : std_logic;
signal \N__59122\ : std_logic;
signal \N__59119\ : std_logic;
signal \N__59116\ : std_logic;
signal \N__59109\ : std_logic;
signal \N__59106\ : std_logic;
signal \N__59105\ : std_logic;
signal \N__59102\ : std_logic;
signal \N__59099\ : std_logic;
signal \N__59096\ : std_logic;
signal \N__59093\ : std_logic;
signal \N__59088\ : std_logic;
signal \N__59085\ : std_logic;
signal \N__59082\ : std_logic;
signal \N__59081\ : std_logic;
signal \N__59078\ : std_logic;
signal \N__59075\ : std_logic;
signal \N__59072\ : std_logic;
signal \N__59069\ : std_logic;
signal \N__59064\ : std_logic;
signal \N__59061\ : std_logic;
signal \N__59058\ : std_logic;
signal \N__59057\ : std_logic;
signal \N__59054\ : std_logic;
signal \N__59053\ : std_logic;
signal \N__59050\ : std_logic;
signal \N__59047\ : std_logic;
signal \N__59044\ : std_logic;
signal \N__59039\ : std_logic;
signal \N__59034\ : std_logic;
signal \N__59031\ : std_logic;
signal \N__59028\ : std_logic;
signal \N__59025\ : std_logic;
signal \N__59022\ : std_logic;
signal \N__59019\ : std_logic;
signal \N__59018\ : std_logic;
signal \N__59015\ : std_logic;
signal \N__59012\ : std_logic;
signal \N__59011\ : std_logic;
signal \N__59010\ : std_logic;
signal \N__59005\ : std_logic;
signal \N__59002\ : std_logic;
signal \N__59001\ : std_logic;
signal \N__58998\ : std_logic;
signal \N__58995\ : std_logic;
signal \N__58990\ : std_logic;
signal \N__58983\ : std_logic;
signal \N__58980\ : std_logic;
signal \N__58979\ : std_logic;
signal \N__58974\ : std_logic;
signal \N__58971\ : std_logic;
signal \N__58968\ : std_logic;
signal \N__58967\ : std_logic;
signal \N__58966\ : std_logic;
signal \N__58963\ : std_logic;
signal \N__58960\ : std_logic;
signal \N__58957\ : std_logic;
signal \N__58952\ : std_logic;
signal \N__58949\ : std_logic;
signal \N__58946\ : std_logic;
signal \N__58943\ : std_logic;
signal \N__58938\ : std_logic;
signal \N__58937\ : std_logic;
signal \N__58934\ : std_logic;
signal \N__58931\ : std_logic;
signal \N__58930\ : std_logic;
signal \N__58927\ : std_logic;
signal \N__58924\ : std_logic;
signal \N__58921\ : std_logic;
signal \N__58918\ : std_logic;
signal \N__58915\ : std_logic;
signal \N__58912\ : std_logic;
signal \N__58907\ : std_logic;
signal \N__58902\ : std_logic;
signal \N__58899\ : std_logic;
signal \N__58896\ : std_logic;
signal \N__58893\ : std_logic;
signal \N__58892\ : std_logic;
signal \N__58891\ : std_logic;
signal \N__58890\ : std_logic;
signal \N__58887\ : std_logic;
signal \N__58884\ : std_logic;
signal \N__58879\ : std_logic;
signal \N__58872\ : std_logic;
signal \N__58871\ : std_logic;
signal \N__58868\ : std_logic;
signal \N__58865\ : std_logic;
signal \N__58862\ : std_logic;
signal \N__58859\ : std_logic;
signal \N__58854\ : std_logic;
signal \N__58851\ : std_logic;
signal \N__58848\ : std_logic;
signal \N__58847\ : std_logic;
signal \N__58844\ : std_logic;
signal \N__58843\ : std_logic;
signal \N__58836\ : std_logic;
signal \N__58833\ : std_logic;
signal \N__58830\ : std_logic;
signal \N__58829\ : std_logic;
signal \N__58828\ : std_logic;
signal \N__58825\ : std_logic;
signal \N__58822\ : std_logic;
signal \N__58821\ : std_logic;
signal \N__58818\ : std_logic;
signal \N__58815\ : std_logic;
signal \N__58810\ : std_logic;
signal \N__58803\ : std_logic;
signal \N__58800\ : std_logic;
signal \N__58797\ : std_logic;
signal \N__58794\ : std_logic;
signal \N__58791\ : std_logic;
signal \N__58788\ : std_logic;
signal \N__58785\ : std_logic;
signal \N__58782\ : std_logic;
signal \N__58779\ : std_logic;
signal \N__58778\ : std_logic;
signal \N__58777\ : std_logic;
signal \N__58776\ : std_logic;
signal \N__58775\ : std_logic;
signal \N__58768\ : std_logic;
signal \N__58767\ : std_logic;
signal \N__58764\ : std_logic;
signal \N__58761\ : std_logic;
signal \N__58758\ : std_logic;
signal \N__58755\ : std_logic;
signal \N__58752\ : std_logic;
signal \N__58751\ : std_logic;
signal \N__58748\ : std_logic;
signal \N__58743\ : std_logic;
signal \N__58740\ : std_logic;
signal \N__58737\ : std_logic;
signal \N__58732\ : std_logic;
signal \N__58725\ : std_logic;
signal \N__58722\ : std_logic;
signal \N__58719\ : std_logic;
signal \N__58716\ : std_logic;
signal \N__58715\ : std_logic;
signal \N__58712\ : std_logic;
signal \N__58709\ : std_logic;
signal \N__58704\ : std_logic;
signal \N__58701\ : std_logic;
signal \N__58700\ : std_logic;
signal \N__58697\ : std_logic;
signal \N__58694\ : std_logic;
signal \N__58689\ : std_logic;
signal \N__58686\ : std_logic;
signal \N__58683\ : std_logic;
signal \N__58680\ : std_logic;
signal \N__58677\ : std_logic;
signal \N__58674\ : std_logic;
signal \N__58671\ : std_logic;
signal \N__58670\ : std_logic;
signal \N__58669\ : std_logic;
signal \N__58666\ : std_logic;
signal \N__58663\ : std_logic;
signal \N__58662\ : std_logic;
signal \N__58659\ : std_logic;
signal \N__58656\ : std_logic;
signal \N__58651\ : std_logic;
signal \N__58646\ : std_logic;
signal \N__58643\ : std_logic;
signal \N__58638\ : std_logic;
signal \N__58635\ : std_logic;
signal \N__58632\ : std_logic;
signal \N__58629\ : std_logic;
signal \N__58626\ : std_logic;
signal \N__58623\ : std_logic;
signal \N__58620\ : std_logic;
signal \N__58619\ : std_logic;
signal \N__58618\ : std_logic;
signal \N__58615\ : std_logic;
signal \N__58614\ : std_logic;
signal \N__58611\ : std_logic;
signal \N__58608\ : std_logic;
signal \N__58605\ : std_logic;
signal \N__58602\ : std_logic;
signal \N__58599\ : std_logic;
signal \N__58594\ : std_logic;
signal \N__58587\ : std_logic;
signal \N__58584\ : std_logic;
signal \N__58581\ : std_logic;
signal \N__58578\ : std_logic;
signal \N__58575\ : std_logic;
signal \N__58572\ : std_logic;
signal \N__58569\ : std_logic;
signal \N__58566\ : std_logic;
signal \N__58563\ : std_logic;
signal \N__58560\ : std_logic;
signal \N__58557\ : std_logic;
signal \N__58554\ : std_logic;
signal \N__58551\ : std_logic;
signal \N__58548\ : std_logic;
signal \N__58545\ : std_logic;
signal \N__58544\ : std_logic;
signal \N__58541\ : std_logic;
signal \N__58538\ : std_logic;
signal \N__58535\ : std_logic;
signal \N__58532\ : std_logic;
signal \N__58527\ : std_logic;
signal \N__58524\ : std_logic;
signal \N__58523\ : std_logic;
signal \N__58520\ : std_logic;
signal \N__58517\ : std_logic;
signal \N__58514\ : std_logic;
signal \N__58511\ : std_logic;
signal \N__58506\ : std_logic;
signal \N__58503\ : std_logic;
signal \N__58500\ : std_logic;
signal \N__58497\ : std_logic;
signal \N__58496\ : std_logic;
signal \N__58493\ : std_logic;
signal \N__58490\ : std_logic;
signal \N__58485\ : std_logic;
signal \N__58482\ : std_logic;
signal \N__58479\ : std_logic;
signal \N__58476\ : std_logic;
signal \N__58473\ : std_logic;
signal \N__58472\ : std_logic;
signal \N__58469\ : std_logic;
signal \N__58466\ : std_logic;
signal \N__58461\ : std_logic;
signal \N__58458\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58451\ : std_logic;
signal \N__58448\ : std_logic;
signal \N__58447\ : std_logic;
signal \N__58444\ : std_logic;
signal \N__58441\ : std_logic;
signal \N__58438\ : std_logic;
signal \N__58435\ : std_logic;
signal \N__58430\ : std_logic;
signal \N__58425\ : std_logic;
signal \N__58422\ : std_logic;
signal \N__58419\ : std_logic;
signal \N__58416\ : std_logic;
signal \N__58413\ : std_logic;
signal \N__58410\ : std_logic;
signal \N__58407\ : std_logic;
signal \N__58404\ : std_logic;
signal \N__58403\ : std_logic;
signal \N__58400\ : std_logic;
signal \N__58399\ : std_logic;
signal \N__58396\ : std_logic;
signal \N__58395\ : std_logic;
signal \N__58392\ : std_logic;
signal \N__58387\ : std_logic;
signal \N__58384\ : std_logic;
signal \N__58377\ : std_logic;
signal \N__58374\ : std_logic;
signal \N__58373\ : std_logic;
signal \N__58372\ : std_logic;
signal \N__58369\ : std_logic;
signal \N__58366\ : std_logic;
signal \N__58363\ : std_logic;
signal \N__58360\ : std_logic;
signal \N__58355\ : std_logic;
signal \N__58350\ : std_logic;
signal \N__58347\ : std_logic;
signal \N__58344\ : std_logic;
signal \N__58341\ : std_logic;
signal \N__58338\ : std_logic;
signal \N__58335\ : std_logic;
signal \N__58332\ : std_logic;
signal \N__58331\ : std_logic;
signal \N__58326\ : std_logic;
signal \N__58323\ : std_logic;
signal \N__58320\ : std_logic;
signal \N__58317\ : std_logic;
signal \N__58314\ : std_logic;
signal \N__58313\ : std_logic;
signal \N__58308\ : std_logic;
signal \N__58305\ : std_logic;
signal \N__58304\ : std_logic;
signal \N__58301\ : std_logic;
signal \N__58298\ : std_logic;
signal \N__58295\ : std_logic;
signal \N__58292\ : std_logic;
signal \N__58289\ : std_logic;
signal \N__58284\ : std_logic;
signal \N__58281\ : std_logic;
signal \N__58280\ : std_logic;
signal \N__58279\ : std_logic;
signal \N__58274\ : std_logic;
signal \N__58271\ : std_logic;
signal \N__58268\ : std_logic;
signal \N__58263\ : std_logic;
signal \N__58260\ : std_logic;
signal \N__58257\ : std_logic;
signal \N__58254\ : std_logic;
signal \N__58253\ : std_logic;
signal \N__58250\ : std_logic;
signal \N__58247\ : std_logic;
signal \N__58242\ : std_logic;
signal \N__58239\ : std_logic;
signal \N__58236\ : std_logic;
signal \N__58233\ : std_logic;
signal \N__58230\ : std_logic;
signal \N__58227\ : std_logic;
signal \N__58224\ : std_logic;
signal \N__58221\ : std_logic;
signal \N__58218\ : std_logic;
signal \N__58215\ : std_logic;
signal \N__58212\ : std_logic;
signal \N__58209\ : std_logic;
signal \N__58206\ : std_logic;
signal \N__58203\ : std_logic;
signal \N__58200\ : std_logic;
signal \N__58199\ : std_logic;
signal \N__58196\ : std_logic;
signal \N__58193\ : std_logic;
signal \N__58190\ : std_logic;
signal \N__58187\ : std_logic;
signal \N__58184\ : std_logic;
signal \N__58181\ : std_logic;
signal \N__58178\ : std_logic;
signal \N__58173\ : std_logic;
signal \N__58170\ : std_logic;
signal \N__58169\ : std_logic;
signal \N__58166\ : std_logic;
signal \N__58163\ : std_logic;
signal \N__58162\ : std_logic;
signal \N__58159\ : std_logic;
signal \N__58156\ : std_logic;
signal \N__58155\ : std_logic;
signal \N__58152\ : std_logic;
signal \N__58147\ : std_logic;
signal \N__58144\ : std_logic;
signal \N__58137\ : std_logic;
signal \N__58136\ : std_logic;
signal \N__58133\ : std_logic;
signal \N__58132\ : std_logic;
signal \N__58129\ : std_logic;
signal \N__58128\ : std_logic;
signal \N__58125\ : std_logic;
signal \N__58122\ : std_logic;
signal \N__58119\ : std_logic;
signal \N__58116\ : std_logic;
signal \N__58113\ : std_logic;
signal \N__58108\ : std_logic;
signal \N__58101\ : std_logic;
signal \N__58098\ : std_logic;
signal \N__58097\ : std_logic;
signal \N__58094\ : std_logic;
signal \N__58091\ : std_logic;
signal \N__58090\ : std_logic;
signal \N__58087\ : std_logic;
signal \N__58084\ : std_logic;
signal \N__58081\ : std_logic;
signal \N__58080\ : std_logic;
signal \N__58079\ : std_logic;
signal \N__58078\ : std_logic;
signal \N__58075\ : std_logic;
signal \N__58072\ : std_logic;
signal \N__58063\ : std_logic;
signal \N__58056\ : std_logic;
signal \N__58055\ : std_logic;
signal \N__58054\ : std_logic;
signal \N__58053\ : std_logic;
signal \N__58052\ : std_logic;
signal \N__58051\ : std_logic;
signal \N__58050\ : std_logic;
signal \N__58049\ : std_logic;
signal \N__58048\ : std_logic;
signal \N__58047\ : std_logic;
signal \N__58044\ : std_logic;
signal \N__58043\ : std_logic;
signal \N__58040\ : std_logic;
signal \N__58037\ : std_logic;
signal \N__58026\ : std_logic;
signal \N__58021\ : std_logic;
signal \N__58018\ : std_logic;
signal \N__58015\ : std_logic;
signal \N__58014\ : std_logic;
signal \N__58013\ : std_logic;
signal \N__58012\ : std_logic;
signal \N__58009\ : std_logic;
signal \N__58002\ : std_logic;
signal \N__57999\ : std_logic;
signal \N__57996\ : std_logic;
signal \N__57993\ : std_logic;
signal \N__57988\ : std_logic;
signal \N__57983\ : std_logic;
signal \N__57972\ : std_logic;
signal \N__57969\ : std_logic;
signal \N__57966\ : std_logic;
signal \N__57963\ : std_logic;
signal \N__57960\ : std_logic;
signal \N__57959\ : std_logic;
signal \N__57958\ : std_logic;
signal \N__57957\ : std_logic;
signal \N__57952\ : std_logic;
signal \N__57951\ : std_logic;
signal \N__57950\ : std_logic;
signal \N__57949\ : std_logic;
signal \N__57946\ : std_logic;
signal \N__57943\ : std_logic;
signal \N__57942\ : std_logic;
signal \N__57939\ : std_logic;
signal \N__57934\ : std_logic;
signal \N__57931\ : std_logic;
signal \N__57930\ : std_logic;
signal \N__57925\ : std_logic;
signal \N__57922\ : std_logic;
signal \N__57917\ : std_logic;
signal \N__57912\ : std_logic;
signal \N__57909\ : std_logic;
signal \N__57900\ : std_logic;
signal \N__57897\ : std_logic;
signal \N__57894\ : std_logic;
signal \N__57891\ : std_logic;
signal \N__57888\ : std_logic;
signal \N__57887\ : std_logic;
signal \N__57886\ : std_logic;
signal \N__57883\ : std_logic;
signal \N__57878\ : std_logic;
signal \N__57875\ : std_logic;
signal \N__57872\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57864\ : std_logic;
signal \N__57861\ : std_logic;
signal \N__57858\ : std_logic;
signal \N__57855\ : std_logic;
signal \N__57852\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57846\ : std_logic;
signal \N__57843\ : std_logic;
signal \N__57840\ : std_logic;
signal \N__57837\ : std_logic;
signal \N__57834\ : std_logic;
signal \N__57831\ : std_logic;
signal \N__57828\ : std_logic;
signal \N__57825\ : std_logic;
signal \N__57822\ : std_logic;
signal \N__57819\ : std_logic;
signal \N__57816\ : std_logic;
signal \N__57813\ : std_logic;
signal \N__57810\ : std_logic;
signal \N__57807\ : std_logic;
signal \N__57804\ : std_logic;
signal \N__57801\ : std_logic;
signal \N__57800\ : std_logic;
signal \N__57797\ : std_logic;
signal \N__57794\ : std_logic;
signal \N__57791\ : std_logic;
signal \N__57788\ : std_logic;
signal \N__57783\ : std_logic;
signal \N__57782\ : std_logic;
signal \N__57779\ : std_logic;
signal \N__57776\ : std_logic;
signal \N__57773\ : std_logic;
signal \N__57768\ : std_logic;
signal \N__57765\ : std_logic;
signal \N__57762\ : std_logic;
signal \N__57759\ : std_logic;
signal \N__57756\ : std_logic;
signal \N__57753\ : std_logic;
signal \N__57750\ : std_logic;
signal \N__57747\ : std_logic;
signal \N__57744\ : std_logic;
signal \N__57741\ : std_logic;
signal \N__57738\ : std_logic;
signal \N__57735\ : std_logic;
signal \N__57732\ : std_logic;
signal \N__57731\ : std_logic;
signal \N__57730\ : std_logic;
signal \N__57729\ : std_logic;
signal \N__57728\ : std_logic;
signal \N__57725\ : std_logic;
signal \N__57722\ : std_logic;
signal \N__57721\ : std_logic;
signal \N__57714\ : std_logic;
signal \N__57711\ : std_logic;
signal \N__57708\ : std_logic;
signal \N__57705\ : std_logic;
signal \N__57702\ : std_logic;
signal \N__57699\ : std_logic;
signal \N__57694\ : std_logic;
signal \N__57691\ : std_logic;
signal \N__57684\ : std_logic;
signal \N__57683\ : std_logic;
signal \N__57678\ : std_logic;
signal \N__57675\ : std_logic;
signal \N__57672\ : std_logic;
signal \N__57671\ : std_logic;
signal \N__57668\ : std_logic;
signal \N__57667\ : std_logic;
signal \N__57664\ : std_logic;
signal \N__57663\ : std_logic;
signal \N__57662\ : std_logic;
signal \N__57661\ : std_logic;
signal \N__57658\ : std_logic;
signal \N__57655\ : std_logic;
signal \N__57650\ : std_logic;
signal \N__57647\ : std_logic;
signal \N__57644\ : std_logic;
signal \N__57639\ : std_logic;
signal \N__57638\ : std_logic;
signal \N__57637\ : std_logic;
signal \N__57636\ : std_logic;
signal \N__57633\ : std_logic;
signal \N__57628\ : std_logic;
signal \N__57625\ : std_logic;
signal \N__57620\ : std_logic;
signal \N__57617\ : std_logic;
signal \N__57606\ : std_logic;
signal \N__57603\ : std_logic;
signal \N__57600\ : std_logic;
signal \N__57597\ : std_logic;
signal \N__57594\ : std_logic;
signal \N__57593\ : std_logic;
signal \N__57592\ : std_logic;
signal \N__57589\ : std_logic;
signal \N__57584\ : std_logic;
signal \N__57579\ : std_logic;
signal \N__57576\ : std_logic;
signal \N__57573\ : std_logic;
signal \N__57570\ : std_logic;
signal \N__57567\ : std_logic;
signal \N__57564\ : std_logic;
signal \N__57563\ : std_logic;
signal \N__57562\ : std_logic;
signal \N__57559\ : std_logic;
signal \N__57554\ : std_logic;
signal \N__57551\ : std_logic;
signal \N__57548\ : std_logic;
signal \N__57545\ : std_logic;
signal \N__57542\ : std_logic;
signal \N__57537\ : std_logic;
signal \N__57536\ : std_logic;
signal \N__57535\ : std_logic;
signal \N__57532\ : std_logic;
signal \N__57529\ : std_logic;
signal \N__57526\ : std_logic;
signal \N__57523\ : std_logic;
signal \N__57520\ : std_logic;
signal \N__57517\ : std_logic;
signal \N__57510\ : std_logic;
signal \N__57507\ : std_logic;
signal \N__57504\ : std_logic;
signal \N__57501\ : std_logic;
signal \N__57498\ : std_logic;
signal \N__57495\ : std_logic;
signal \N__57494\ : std_logic;
signal \N__57489\ : std_logic;
signal \N__57488\ : std_logic;
signal \N__57485\ : std_logic;
signal \N__57484\ : std_logic;
signal \N__57483\ : std_logic;
signal \N__57480\ : std_logic;
signal \N__57477\ : std_logic;
signal \N__57474\ : std_logic;
signal \N__57469\ : std_logic;
signal \N__57462\ : std_logic;
signal \N__57461\ : std_logic;
signal \N__57460\ : std_logic;
signal \N__57457\ : std_logic;
signal \N__57450\ : std_logic;
signal \N__57447\ : std_logic;
signal \N__57444\ : std_logic;
signal \N__57441\ : std_logic;
signal \N__57438\ : std_logic;
signal \N__57435\ : std_logic;
signal \N__57432\ : std_logic;
signal \N__57429\ : std_logic;
signal \N__57428\ : std_logic;
signal \N__57425\ : std_logic;
signal \N__57422\ : std_logic;
signal \N__57417\ : std_logic;
signal \N__57416\ : std_logic;
signal \N__57413\ : std_logic;
signal \N__57410\ : std_logic;
signal \N__57409\ : std_logic;
signal \N__57406\ : std_logic;
signal \N__57403\ : std_logic;
signal \N__57400\ : std_logic;
signal \N__57399\ : std_logic;
signal \N__57396\ : std_logic;
signal \N__57393\ : std_logic;
signal \N__57388\ : std_logic;
signal \N__57381\ : std_logic;
signal \N__57378\ : std_logic;
signal \N__57377\ : std_logic;
signal \N__57376\ : std_logic;
signal \N__57373\ : std_logic;
signal \N__57370\ : std_logic;
signal \N__57367\ : std_logic;
signal \N__57366\ : std_logic;
signal \N__57365\ : std_logic;
signal \N__57362\ : std_logic;
signal \N__57359\ : std_logic;
signal \N__57356\ : std_logic;
signal \N__57355\ : std_logic;
signal \N__57352\ : std_logic;
signal \N__57349\ : std_logic;
signal \N__57346\ : std_logic;
signal \N__57343\ : std_logic;
signal \N__57340\ : std_logic;
signal \N__57337\ : std_logic;
signal \N__57324\ : std_logic;
signal \N__57323\ : std_logic;
signal \N__57322\ : std_logic;
signal \N__57319\ : std_logic;
signal \N__57314\ : std_logic;
signal \N__57309\ : std_logic;
signal \N__57308\ : std_logic;
signal \N__57305\ : std_logic;
signal \N__57302\ : std_logic;
signal \N__57299\ : std_logic;
signal \N__57298\ : std_logic;
signal \N__57297\ : std_logic;
signal \N__57294\ : std_logic;
signal \N__57291\ : std_logic;
signal \N__57286\ : std_logic;
signal \N__57283\ : std_logic;
signal \N__57280\ : std_logic;
signal \N__57277\ : std_logic;
signal \N__57270\ : std_logic;
signal \N__57267\ : std_logic;
signal \N__57264\ : std_logic;
signal \N__57263\ : std_logic;
signal \N__57260\ : std_logic;
signal \N__57257\ : std_logic;
signal \N__57254\ : std_logic;
signal \N__57251\ : std_logic;
signal \N__57246\ : std_logic;
signal \N__57245\ : std_logic;
signal \N__57244\ : std_logic;
signal \N__57243\ : std_logic;
signal \N__57240\ : std_logic;
signal \N__57237\ : std_logic;
signal \N__57236\ : std_logic;
signal \N__57235\ : std_logic;
signal \N__57234\ : std_logic;
signal \N__57233\ : std_logic;
signal \N__57232\ : std_logic;
signal \N__57229\ : std_logic;
signal \N__57228\ : std_logic;
signal \N__57225\ : std_logic;
signal \N__57220\ : std_logic;
signal \N__57213\ : std_logic;
signal \N__57208\ : std_logic;
signal \N__57203\ : std_logic;
signal \N__57192\ : std_logic;
signal \N__57189\ : std_logic;
signal \N__57186\ : std_logic;
signal \N__57183\ : std_logic;
signal \N__57180\ : std_logic;
signal \N__57177\ : std_logic;
signal \N__57174\ : std_logic;
signal \N__57171\ : std_logic;
signal \N__57168\ : std_logic;
signal \N__57165\ : std_logic;
signal \N__57162\ : std_logic;
signal \N__57159\ : std_logic;
signal \N__57156\ : std_logic;
signal \N__57155\ : std_logic;
signal \N__57152\ : std_logic;
signal \N__57149\ : std_logic;
signal \N__57146\ : std_logic;
signal \N__57143\ : std_logic;
signal \N__57140\ : std_logic;
signal \N__57137\ : std_logic;
signal \N__57134\ : std_logic;
signal \N__57129\ : std_logic;
signal \N__57126\ : std_logic;
signal \N__57123\ : std_logic;
signal \N__57120\ : std_logic;
signal \N__57117\ : std_logic;
signal \N__57114\ : std_logic;
signal \N__57113\ : std_logic;
signal \N__57112\ : std_logic;
signal \N__57109\ : std_logic;
signal \N__57106\ : std_logic;
signal \N__57103\ : std_logic;
signal \N__57102\ : std_logic;
signal \N__57099\ : std_logic;
signal \N__57096\ : std_logic;
signal \N__57091\ : std_logic;
signal \N__57088\ : std_logic;
signal \N__57081\ : std_logic;
signal \N__57080\ : std_logic;
signal \N__57077\ : std_logic;
signal \N__57076\ : std_logic;
signal \N__57073\ : std_logic;
signal \N__57072\ : std_logic;
signal \N__57069\ : std_logic;
signal \N__57066\ : std_logic;
signal \N__57063\ : std_logic;
signal \N__57060\ : std_logic;
signal \N__57053\ : std_logic;
signal \N__57048\ : std_logic;
signal \N__57045\ : std_logic;
signal \N__57042\ : std_logic;
signal \N__57039\ : std_logic;
signal \N__57036\ : std_logic;
signal \N__57033\ : std_logic;
signal \N__57030\ : std_logic;
signal \N__57027\ : std_logic;
signal \N__57024\ : std_logic;
signal \N__57021\ : std_logic;
signal \N__57018\ : std_logic;
signal \N__57017\ : std_logic;
signal \N__57016\ : std_logic;
signal \N__57015\ : std_logic;
signal \N__57014\ : std_logic;
signal \N__57011\ : std_logic;
signal \N__57002\ : std_logic;
signal \N__57001\ : std_logic;
signal \N__56998\ : std_logic;
signal \N__56995\ : std_logic;
signal \N__56994\ : std_logic;
signal \N__56991\ : std_logic;
signal \N__56988\ : std_logic;
signal \N__56985\ : std_logic;
signal \N__56980\ : std_logic;
signal \N__56973\ : std_logic;
signal \N__56970\ : std_logic;
signal \N__56967\ : std_logic;
signal \N__56964\ : std_logic;
signal \N__56961\ : std_logic;
signal \N__56958\ : std_logic;
signal \N__56955\ : std_logic;
signal \N__56952\ : std_logic;
signal \N__56949\ : std_logic;
signal \N__56946\ : std_logic;
signal \N__56943\ : std_logic;
signal \N__56940\ : std_logic;
signal \N__56937\ : std_logic;
signal \N__56934\ : std_logic;
signal \N__56931\ : std_logic;
signal \N__56928\ : std_logic;
signal \N__56925\ : std_logic;
signal \N__56922\ : std_logic;
signal \N__56919\ : std_logic;
signal \N__56916\ : std_logic;
signal \N__56913\ : std_logic;
signal \N__56910\ : std_logic;
signal \N__56907\ : std_logic;
signal \N__56904\ : std_logic;
signal \N__56903\ : std_logic;
signal \N__56898\ : std_logic;
signal \N__56895\ : std_logic;
signal \N__56894\ : std_logic;
signal \N__56893\ : std_logic;
signal \N__56890\ : std_logic;
signal \N__56887\ : std_logic;
signal \N__56886\ : std_logic;
signal \N__56883\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56872\ : std_logic;
signal \N__56869\ : std_logic;
signal \N__56862\ : std_logic;
signal \N__56859\ : std_logic;
signal \N__56858\ : std_logic;
signal \N__56855\ : std_logic;
signal \N__56854\ : std_logic;
signal \N__56853\ : std_logic;
signal \N__56850\ : std_logic;
signal \N__56847\ : std_logic;
signal \N__56844\ : std_logic;
signal \N__56841\ : std_logic;
signal \N__56836\ : std_logic;
signal \N__56833\ : std_logic;
signal \N__56830\ : std_logic;
signal \N__56827\ : std_logic;
signal \N__56824\ : std_logic;
signal \N__56817\ : std_logic;
signal \N__56816\ : std_logic;
signal \N__56815\ : std_logic;
signal \N__56814\ : std_logic;
signal \N__56811\ : std_logic;
signal \N__56808\ : std_logic;
signal \N__56805\ : std_logic;
signal \N__56802\ : std_logic;
signal \N__56799\ : std_logic;
signal \N__56798\ : std_logic;
signal \N__56797\ : std_logic;
signal \N__56794\ : std_logic;
signal \N__56791\ : std_logic;
signal \N__56788\ : std_logic;
signal \N__56785\ : std_logic;
signal \N__56780\ : std_logic;
signal \N__56773\ : std_logic;
signal \N__56766\ : std_logic;
signal \N__56763\ : std_logic;
signal \N__56760\ : std_logic;
signal \N__56757\ : std_logic;
signal \N__56754\ : std_logic;
signal \N__56753\ : std_logic;
signal \N__56752\ : std_logic;
signal \N__56751\ : std_logic;
signal \N__56748\ : std_logic;
signal \N__56745\ : std_logic;
signal \N__56742\ : std_logic;
signal \N__56739\ : std_logic;
signal \N__56738\ : std_logic;
signal \N__56737\ : std_logic;
signal \N__56736\ : std_logic;
signal \N__56733\ : std_logic;
signal \N__56726\ : std_logic;
signal \N__56719\ : std_logic;
signal \N__56712\ : std_logic;
signal \N__56709\ : std_logic;
signal \N__56706\ : std_logic;
signal \N__56705\ : std_logic;
signal \N__56702\ : std_logic;
signal \N__56699\ : std_logic;
signal \N__56696\ : std_logic;
signal \N__56691\ : std_logic;
signal \N__56688\ : std_logic;
signal \N__56685\ : std_logic;
signal \N__56684\ : std_logic;
signal \N__56681\ : std_logic;
signal \N__56678\ : std_logic;
signal \N__56675\ : std_logic;
signal \N__56670\ : std_logic;
signal \N__56669\ : std_logic;
signal \N__56666\ : std_logic;
signal \N__56663\ : std_logic;
signal \N__56658\ : std_logic;
signal \N__56655\ : std_logic;
signal \N__56652\ : std_logic;
signal \N__56651\ : std_logic;
signal \N__56650\ : std_logic;
signal \N__56649\ : std_logic;
signal \N__56642\ : std_logic;
signal \N__56639\ : std_logic;
signal \N__56636\ : std_logic;
signal \N__56633\ : std_logic;
signal \N__56632\ : std_logic;
signal \N__56629\ : std_logic;
signal \N__56626\ : std_logic;
signal \N__56623\ : std_logic;
signal \N__56620\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56610\ : std_logic;
signal \N__56607\ : std_logic;
signal \N__56604\ : std_logic;
signal \N__56601\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56595\ : std_logic;
signal \N__56594\ : std_logic;
signal \N__56589\ : std_logic;
signal \N__56588\ : std_logic;
signal \N__56585\ : std_logic;
signal \N__56582\ : std_logic;
signal \N__56579\ : std_logic;
signal \N__56574\ : std_logic;
signal \N__56573\ : std_logic;
signal \N__56572\ : std_logic;
signal \N__56569\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56561\ : std_logic;
signal \N__56560\ : std_logic;
signal \N__56557\ : std_logic;
signal \N__56554\ : std_logic;
signal \N__56551\ : std_logic;
signal \N__56548\ : std_logic;
signal \N__56545\ : std_logic;
signal \N__56542\ : std_logic;
signal \N__56539\ : std_logic;
signal \N__56536\ : std_logic;
signal \N__56529\ : std_logic;
signal \N__56526\ : std_logic;
signal \N__56523\ : std_logic;
signal \N__56522\ : std_logic;
signal \N__56519\ : std_logic;
signal \N__56516\ : std_logic;
signal \N__56515\ : std_logic;
signal \N__56512\ : std_logic;
signal \N__56509\ : std_logic;
signal \N__56506\ : std_logic;
signal \N__56499\ : std_logic;
signal \N__56496\ : std_logic;
signal \N__56493\ : std_logic;
signal \N__56490\ : std_logic;
signal \N__56487\ : std_logic;
signal \N__56484\ : std_logic;
signal \N__56483\ : std_logic;
signal \N__56482\ : std_logic;
signal \N__56481\ : std_logic;
signal \N__56480\ : std_logic;
signal \N__56479\ : std_logic;
signal \N__56476\ : std_logic;
signal \N__56471\ : std_logic;
signal \N__56468\ : std_logic;
signal \N__56465\ : std_logic;
signal \N__56462\ : std_logic;
signal \N__56461\ : std_logic;
signal \N__56456\ : std_logic;
signal \N__56453\ : std_logic;
signal \N__56450\ : std_logic;
signal \N__56445\ : std_logic;
signal \N__56438\ : std_logic;
signal \N__56435\ : std_logic;
signal \N__56432\ : std_logic;
signal \N__56427\ : std_logic;
signal \N__56424\ : std_logic;
signal \N__56421\ : std_logic;
signal \N__56418\ : std_logic;
signal \N__56415\ : std_logic;
signal \N__56412\ : std_logic;
signal \N__56411\ : std_logic;
signal \N__56408\ : std_logic;
signal \N__56407\ : std_logic;
signal \N__56406\ : std_logic;
signal \N__56403\ : std_logic;
signal \N__56400\ : std_logic;
signal \N__56397\ : std_logic;
signal \N__56396\ : std_logic;
signal \N__56393\ : std_logic;
signal \N__56390\ : std_logic;
signal \N__56387\ : std_logic;
signal \N__56382\ : std_logic;
signal \N__56373\ : std_logic;
signal \N__56372\ : std_logic;
signal \N__56371\ : std_logic;
signal \N__56370\ : std_logic;
signal \N__56369\ : std_logic;
signal \N__56366\ : std_logic;
signal \N__56361\ : std_logic;
signal \N__56358\ : std_logic;
signal \N__56355\ : std_logic;
signal \N__56354\ : std_logic;
signal \N__56351\ : std_logic;
signal \N__56348\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56342\ : std_logic;
signal \N__56339\ : std_logic;
signal \N__56334\ : std_logic;
signal \N__56325\ : std_logic;
signal \N__56324\ : std_logic;
signal \N__56323\ : std_logic;
signal \N__56322\ : std_logic;
signal \N__56317\ : std_logic;
signal \N__56312\ : std_logic;
signal \N__56309\ : std_logic;
signal \N__56306\ : std_logic;
signal \N__56303\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56295\ : std_logic;
signal \N__56292\ : std_logic;
signal \N__56289\ : std_logic;
signal \N__56286\ : std_logic;
signal \N__56283\ : std_logic;
signal \N__56280\ : std_logic;
signal \N__56277\ : std_logic;
signal \N__56276\ : std_logic;
signal \N__56273\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56269\ : std_logic;
signal \N__56268\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56262\ : std_logic;
signal \N__56259\ : std_logic;
signal \N__56256\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56244\ : std_logic;
signal \N__56241\ : std_logic;
signal \N__56240\ : std_logic;
signal \N__56239\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56223\ : std_logic;
signal \N__56220\ : std_logic;
signal \N__56217\ : std_logic;
signal \N__56214\ : std_logic;
signal \N__56211\ : std_logic;
signal \N__56208\ : std_logic;
signal \N__56203\ : std_logic;
signal \N__56196\ : std_logic;
signal \N__56193\ : std_logic;
signal \N__56192\ : std_logic;
signal \N__56189\ : std_logic;
signal \N__56186\ : std_logic;
signal \N__56185\ : std_logic;
signal \N__56182\ : std_logic;
signal \N__56179\ : std_logic;
signal \N__56176\ : std_logic;
signal \N__56171\ : std_logic;
signal \N__56166\ : std_logic;
signal \N__56163\ : std_logic;
signal \N__56160\ : std_logic;
signal \N__56159\ : std_logic;
signal \N__56156\ : std_logic;
signal \N__56153\ : std_logic;
signal \N__56148\ : std_logic;
signal \N__56147\ : std_logic;
signal \N__56144\ : std_logic;
signal \N__56143\ : std_logic;
signal \N__56140\ : std_logic;
signal \N__56139\ : std_logic;
signal \N__56136\ : std_logic;
signal \N__56133\ : std_logic;
signal \N__56130\ : std_logic;
signal \N__56127\ : std_logic;
signal \N__56124\ : std_logic;
signal \N__56119\ : std_logic;
signal \N__56112\ : std_logic;
signal \N__56109\ : std_logic;
signal \N__56106\ : std_logic;
signal \N__56103\ : std_logic;
signal \N__56100\ : std_logic;
signal \N__56097\ : std_logic;
signal \N__56094\ : std_logic;
signal \N__56091\ : std_logic;
signal \N__56088\ : std_logic;
signal \N__56085\ : std_logic;
signal \N__56084\ : std_logic;
signal \N__56079\ : std_logic;
signal \N__56076\ : std_logic;
signal \N__56073\ : std_logic;
signal \N__56072\ : std_logic;
signal \N__56069\ : std_logic;
signal \N__56066\ : std_logic;
signal \N__56063\ : std_logic;
signal \N__56060\ : std_logic;
signal \N__56057\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56051\ : std_logic;
signal \N__56048\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56039\ : std_logic;
signal \N__56038\ : std_logic;
signal \N__56035\ : std_logic;
signal \N__56030\ : std_logic;
signal \N__56027\ : std_logic;
signal \N__56022\ : std_logic;
signal \N__56019\ : std_logic;
signal \N__56016\ : std_logic;
signal \N__56013\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56009\ : std_logic;
signal \N__56006\ : std_logic;
signal \N__56005\ : std_logic;
signal \N__56002\ : std_logic;
signal \N__55999\ : std_logic;
signal \N__55994\ : std_logic;
signal \N__55991\ : std_logic;
signal \N__55988\ : std_logic;
signal \N__55983\ : std_logic;
signal \N__55980\ : std_logic;
signal \N__55977\ : std_logic;
signal \N__55976\ : std_logic;
signal \N__55973\ : std_logic;
signal \N__55972\ : std_logic;
signal \N__55969\ : std_logic;
signal \N__55966\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55962\ : std_logic;
signal \N__55959\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55953\ : std_logic;
signal \N__55944\ : std_logic;
signal \N__55943\ : std_logic;
signal \N__55938\ : std_logic;
signal \N__55935\ : std_logic;
signal \N__55932\ : std_logic;
signal \N__55931\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55923\ : std_logic;
signal \N__55920\ : std_logic;
signal \N__55919\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55913\ : std_logic;
signal \N__55910\ : std_logic;
signal \N__55905\ : std_logic;
signal \N__55902\ : std_logic;
signal \N__55901\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55899\ : std_logic;
signal \N__55898\ : std_logic;
signal \N__55889\ : std_logic;
signal \N__55886\ : std_logic;
signal \N__55883\ : std_logic;
signal \N__55882\ : std_logic;
signal \N__55879\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55866\ : std_logic;
signal \N__55863\ : std_logic;
signal \N__55860\ : std_logic;
signal \N__55857\ : std_logic;
signal \N__55854\ : std_logic;
signal \N__55851\ : std_logic;
signal \N__55848\ : std_logic;
signal \N__55845\ : std_logic;
signal \N__55842\ : std_logic;
signal \N__55839\ : std_logic;
signal \N__55838\ : std_logic;
signal \N__55835\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55827\ : std_logic;
signal \N__55824\ : std_logic;
signal \N__55823\ : std_logic;
signal \N__55820\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55814\ : std_logic;
signal \N__55811\ : std_logic;
signal \N__55808\ : std_logic;
signal \N__55803\ : std_logic;
signal \N__55800\ : std_logic;
signal \N__55799\ : std_logic;
signal \N__55798\ : std_logic;
signal \N__55797\ : std_logic;
signal \N__55790\ : std_logic;
signal \N__55787\ : std_logic;
signal \N__55782\ : std_logic;
signal \N__55779\ : std_logic;
signal \N__55776\ : std_logic;
signal \N__55775\ : std_logic;
signal \N__55770\ : std_logic;
signal \N__55767\ : std_logic;
signal \N__55766\ : std_logic;
signal \N__55761\ : std_logic;
signal \N__55760\ : std_logic;
signal \N__55757\ : std_logic;
signal \N__55754\ : std_logic;
signal \N__55751\ : std_logic;
signal \N__55746\ : std_logic;
signal \N__55743\ : std_logic;
signal \N__55742\ : std_logic;
signal \N__55741\ : std_logic;
signal \N__55740\ : std_logic;
signal \N__55737\ : std_logic;
signal \N__55734\ : std_logic;
signal \N__55731\ : std_logic;
signal \N__55728\ : std_logic;
signal \N__55727\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55721\ : std_logic;
signal \N__55718\ : std_logic;
signal \N__55715\ : std_logic;
signal \N__55712\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55704\ : std_logic;
signal \N__55701\ : std_logic;
signal \N__55698\ : std_logic;
signal \N__55695\ : std_logic;
signal \N__55686\ : std_logic;
signal \N__55683\ : std_logic;
signal \N__55682\ : std_logic;
signal \N__55679\ : std_logic;
signal \N__55676\ : std_logic;
signal \N__55673\ : std_logic;
signal \N__55670\ : std_logic;
signal \N__55665\ : std_logic;
signal \N__55664\ : std_logic;
signal \N__55661\ : std_logic;
signal \N__55658\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55647\ : std_logic;
signal \N__55644\ : std_logic;
signal \N__55641\ : std_logic;
signal \N__55638\ : std_logic;
signal \N__55635\ : std_logic;
signal \N__55632\ : std_logic;
signal \N__55631\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55627\ : std_logic;
signal \N__55624\ : std_logic;
signal \N__55621\ : std_logic;
signal \N__55618\ : std_logic;
signal \N__55615\ : std_logic;
signal \N__55612\ : std_logic;
signal \N__55611\ : std_logic;
signal \N__55604\ : std_logic;
signal \N__55601\ : std_logic;
signal \N__55598\ : std_logic;
signal \N__55593\ : std_logic;
signal \N__55590\ : std_logic;
signal \N__55587\ : std_logic;
signal \N__55584\ : std_logic;
signal \N__55581\ : std_logic;
signal \N__55578\ : std_logic;
signal \N__55575\ : std_logic;
signal \N__55572\ : std_logic;
signal \N__55569\ : std_logic;
signal \N__55566\ : std_logic;
signal \N__55565\ : std_logic;
signal \N__55564\ : std_logic;
signal \N__55561\ : std_logic;
signal \N__55558\ : std_logic;
signal \N__55555\ : std_logic;
signal \N__55552\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55546\ : std_logic;
signal \N__55543\ : std_logic;
signal \N__55538\ : std_logic;
signal \N__55533\ : std_logic;
signal \N__55530\ : std_logic;
signal \N__55527\ : std_logic;
signal \N__55524\ : std_logic;
signal \N__55523\ : std_logic;
signal \N__55520\ : std_logic;
signal \N__55517\ : std_logic;
signal \N__55514\ : std_logic;
signal \N__55513\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55509\ : std_logic;
signal \N__55508\ : std_logic;
signal \N__55505\ : std_logic;
signal \N__55500\ : std_logic;
signal \N__55497\ : std_logic;
signal \N__55494\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55482\ : std_logic;
signal \N__55479\ : std_logic;
signal \N__55478\ : std_logic;
signal \N__55475\ : std_logic;
signal \N__55472\ : std_logic;
signal \N__55469\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55463\ : std_logic;
signal \N__55460\ : std_logic;
signal \N__55455\ : std_logic;
signal \N__55454\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55442\ : std_logic;
signal \N__55439\ : std_logic;
signal \N__55434\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55429\ : std_logic;
signal \N__55426\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55415\ : std_logic;
signal \N__55410\ : std_logic;
signal \N__55407\ : std_logic;
signal \N__55404\ : std_logic;
signal \N__55401\ : std_logic;
signal \N__55398\ : std_logic;
signal \N__55395\ : std_logic;
signal \N__55392\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55386\ : std_logic;
signal \N__55383\ : std_logic;
signal \N__55380\ : std_logic;
signal \N__55377\ : std_logic;
signal \N__55374\ : std_logic;
signal \N__55371\ : std_logic;
signal \N__55368\ : std_logic;
signal \N__55365\ : std_logic;
signal \N__55362\ : std_logic;
signal \N__55359\ : std_logic;
signal \N__55356\ : std_logic;
signal \N__55353\ : std_logic;
signal \N__55350\ : std_logic;
signal \N__55347\ : std_logic;
signal \N__55344\ : std_logic;
signal \N__55341\ : std_logic;
signal \N__55338\ : std_logic;
signal \N__55335\ : std_logic;
signal \N__55332\ : std_logic;
signal \N__55331\ : std_logic;
signal \N__55330\ : std_logic;
signal \N__55329\ : std_logic;
signal \N__55326\ : std_logic;
signal \N__55323\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55316\ : std_logic;
signal \N__55311\ : std_logic;
signal \N__55308\ : std_logic;
signal \N__55305\ : std_logic;
signal \N__55302\ : std_logic;
signal \N__55297\ : std_logic;
signal \N__55290\ : std_logic;
signal \N__55287\ : std_logic;
signal \N__55284\ : std_logic;
signal \N__55281\ : std_logic;
signal \N__55278\ : std_logic;
signal \N__55275\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55269\ : std_logic;
signal \N__55266\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55260\ : std_logic;
signal \N__55257\ : std_logic;
signal \N__55254\ : std_logic;
signal \N__55251\ : std_logic;
signal \N__55248\ : std_logic;
signal \N__55245\ : std_logic;
signal \N__55242\ : std_logic;
signal \N__55241\ : std_logic;
signal \N__55238\ : std_logic;
signal \N__55235\ : std_logic;
signal \N__55232\ : std_logic;
signal \N__55229\ : std_logic;
signal \N__55226\ : std_logic;
signal \N__55221\ : std_logic;
signal \N__55220\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55214\ : std_logic;
signal \N__55211\ : std_logic;
signal \N__55208\ : std_logic;
signal \N__55207\ : std_logic;
signal \N__55206\ : std_logic;
signal \N__55203\ : std_logic;
signal \N__55200\ : std_logic;
signal \N__55195\ : std_logic;
signal \N__55188\ : std_logic;
signal \N__55187\ : std_logic;
signal \N__55186\ : std_logic;
signal \N__55185\ : std_logic;
signal \N__55184\ : std_logic;
signal \N__55179\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55171\ : std_logic;
signal \N__55168\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55162\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55152\ : std_logic;
signal \N__55149\ : std_logic;
signal \N__55146\ : std_logic;
signal \N__55143\ : std_logic;
signal \N__55140\ : std_logic;
signal \N__55137\ : std_logic;
signal \N__55134\ : std_logic;
signal \N__55133\ : std_logic;
signal \N__55128\ : std_logic;
signal \N__55125\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55121\ : std_logic;
signal \N__55118\ : std_logic;
signal \N__55115\ : std_logic;
signal \N__55114\ : std_logic;
signal \N__55113\ : std_logic;
signal \N__55110\ : std_logic;
signal \N__55107\ : std_logic;
signal \N__55104\ : std_logic;
signal \N__55101\ : std_logic;
signal \N__55100\ : std_logic;
signal \N__55097\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55087\ : std_logic;
signal \N__55080\ : std_logic;
signal \N__55077\ : std_logic;
signal \N__55074\ : std_logic;
signal \N__55071\ : std_logic;
signal \N__55070\ : std_logic;
signal \N__55069\ : std_logic;
signal \N__55066\ : std_logic;
signal \N__55063\ : std_logic;
signal \N__55060\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55050\ : std_logic;
signal \N__55049\ : std_logic;
signal \N__55046\ : std_logic;
signal \N__55045\ : std_logic;
signal \N__55040\ : std_logic;
signal \N__55037\ : std_logic;
signal \N__55034\ : std_logic;
signal \N__55031\ : std_logic;
signal \N__55028\ : std_logic;
signal \N__55023\ : std_logic;
signal \N__55022\ : std_logic;
signal \N__55021\ : std_logic;
signal \N__55020\ : std_logic;
signal \N__55017\ : std_logic;
signal \N__55014\ : std_logic;
signal \N__55009\ : std_logic;
signal \N__55006\ : std_logic;
signal \N__55003\ : std_logic;
signal \N__55000\ : std_logic;
signal \N__54995\ : std_logic;
signal \N__54992\ : std_logic;
signal \N__54987\ : std_logic;
signal \N__54984\ : std_logic;
signal \N__54981\ : std_logic;
signal \N__54978\ : std_logic;
signal \N__54975\ : std_logic;
signal \N__54972\ : std_logic;
signal \N__54969\ : std_logic;
signal \N__54968\ : std_logic;
signal \N__54963\ : std_logic;
signal \N__54960\ : std_logic;
signal \N__54957\ : std_logic;
signal \N__54954\ : std_logic;
signal \N__54951\ : std_logic;
signal \N__54950\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54944\ : std_logic;
signal \N__54943\ : std_logic;
signal \N__54940\ : std_logic;
signal \N__54937\ : std_logic;
signal \N__54936\ : std_logic;
signal \N__54933\ : std_logic;
signal \N__54930\ : std_logic;
signal \N__54927\ : std_logic;
signal \N__54924\ : std_logic;
signal \N__54921\ : std_logic;
signal \N__54918\ : std_logic;
signal \N__54909\ : std_logic;
signal \N__54906\ : std_logic;
signal \N__54903\ : std_logic;
signal \N__54900\ : std_logic;
signal \N__54897\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54891\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54883\ : std_logic;
signal \N__54882\ : std_logic;
signal \N__54881\ : std_logic;
signal \N__54880\ : std_logic;
signal \N__54879\ : std_logic;
signal \N__54872\ : std_logic;
signal \N__54863\ : std_logic;
signal \N__54862\ : std_logic;
signal \N__54861\ : std_logic;
signal \N__54860\ : std_logic;
signal \N__54859\ : std_logic;
signal \N__54858\ : std_logic;
signal \N__54857\ : std_logic;
signal \N__54856\ : std_logic;
signal \N__54855\ : std_logic;
signal \N__54854\ : std_logic;
signal \N__54853\ : std_logic;
signal \N__54852\ : std_logic;
signal \N__54851\ : std_logic;
signal \N__54850\ : std_logic;
signal \N__54849\ : std_logic;
signal \N__54848\ : std_logic;
signal \N__54847\ : std_logic;
signal \N__54846\ : std_logic;
signal \N__54845\ : std_logic;
signal \N__54844\ : std_logic;
signal \N__54843\ : std_logic;
signal \N__54842\ : std_logic;
signal \N__54841\ : std_logic;
signal \N__54840\ : std_logic;
signal \N__54839\ : std_logic;
signal \N__54838\ : std_logic;
signal \N__54837\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54834\ : std_logic;
signal \N__54833\ : std_logic;
signal \N__54832\ : std_logic;
signal \N__54831\ : std_logic;
signal \N__54830\ : std_logic;
signal \N__54829\ : std_logic;
signal \N__54828\ : std_logic;
signal \N__54827\ : std_logic;
signal \N__54822\ : std_logic;
signal \N__54815\ : std_logic;
signal \N__54806\ : std_logic;
signal \N__54799\ : std_logic;
signal \N__54790\ : std_logic;
signal \N__54783\ : std_logic;
signal \N__54774\ : std_logic;
signal \N__54767\ : std_logic;
signal \N__54758\ : std_logic;
signal \N__54755\ : std_logic;
signal \N__54754\ : std_logic;
signal \N__54751\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54746\ : std_logic;
signal \N__54743\ : std_logic;
signal \N__54742\ : std_logic;
signal \N__54741\ : std_logic;
signal \N__54740\ : std_logic;
signal \N__54739\ : std_logic;
signal \N__54738\ : std_logic;
signal \N__54737\ : std_logic;
signal \N__54736\ : std_logic;
signal \N__54733\ : std_logic;
signal \N__54732\ : std_logic;
signal \N__54729\ : std_logic;
signal \N__54728\ : std_logic;
signal \N__54725\ : std_logic;
signal \N__54724\ : std_logic;
signal \N__54721\ : std_logic;
signal \N__54720\ : std_logic;
signal \N__54719\ : std_logic;
signal \N__54718\ : std_logic;
signal \N__54717\ : std_logic;
signal \N__54716\ : std_logic;
signal \N__54715\ : std_logic;
signal \N__54714\ : std_logic;
signal \N__54695\ : std_logic;
signal \N__54680\ : std_logic;
signal \N__54673\ : std_logic;
signal \N__54664\ : std_logic;
signal \N__54649\ : std_logic;
signal \N__54642\ : std_logic;
signal \N__54633\ : std_logic;
signal \N__54632\ : std_logic;
signal \N__54631\ : std_logic;
signal \N__54630\ : std_logic;
signal \N__54615\ : std_logic;
signal \N__54614\ : std_logic;
signal \N__54613\ : std_logic;
signal \N__54612\ : std_logic;
signal \N__54611\ : std_logic;
signal \N__54610\ : std_logic;
signal \N__54609\ : std_logic;
signal \N__54608\ : std_logic;
signal \N__54607\ : std_logic;
signal \N__54606\ : std_logic;
signal \N__54605\ : std_logic;
signal \N__54604\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54602\ : std_logic;
signal \N__54601\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54599\ : std_logic;
signal \N__54598\ : std_logic;
signal \N__54597\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54595\ : std_logic;
signal \N__54594\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54590\ : std_logic;
signal \N__54589\ : std_logic;
signal \N__54586\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54582\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54579\ : std_logic;
signal \N__54578\ : std_logic;
signal \N__54577\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54575\ : std_logic;
signal \N__54574\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54572\ : std_logic;
signal \N__54571\ : std_logic;
signal \N__54570\ : std_logic;
signal \N__54569\ : std_logic;
signal \N__54566\ : std_logic;
signal \N__54559\ : std_logic;
signal \N__54550\ : std_logic;
signal \N__54543\ : std_logic;
signal \N__54534\ : std_logic;
signal \N__54527\ : std_logic;
signal \N__54518\ : std_logic;
signal \N__54517\ : std_logic;
signal \N__54516\ : std_logic;
signal \N__54515\ : std_logic;
signal \N__54514\ : std_logic;
signal \N__54513\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54510\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54508\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54506\ : std_logic;
signal \N__54505\ : std_logic;
signal \N__54504\ : std_logic;
signal \N__54503\ : std_logic;
signal \N__54502\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54500\ : std_logic;
signal \N__54499\ : std_logic;
signal \N__54498\ : std_logic;
signal \N__54497\ : std_logic;
signal \N__54496\ : std_logic;
signal \N__54495\ : std_logic;
signal \N__54494\ : std_logic;
signal \N__54493\ : std_logic;
signal \N__54492\ : std_logic;
signal \N__54491\ : std_logic;
signal \N__54490\ : std_logic;
signal \N__54475\ : std_logic;
signal \N__54474\ : std_logic;
signal \N__54471\ : std_logic;
signal \N__54470\ : std_logic;
signal \N__54467\ : std_logic;
signal \N__54466\ : std_logic;
signal \N__54463\ : std_logic;
signal \N__54462\ : std_logic;
signal \N__54461\ : std_logic;
signal \N__54458\ : std_logic;
signal \N__54457\ : std_logic;
signal \N__54454\ : std_logic;
signal \N__54453\ : std_logic;
signal \N__54450\ : std_logic;
signal \N__54449\ : std_logic;
signal \N__54448\ : std_logic;
signal \N__54445\ : std_logic;
signal \N__54444\ : std_logic;
signal \N__54441\ : std_logic;
signal \N__54440\ : std_logic;
signal \N__54437\ : std_logic;
signal \N__54436\ : std_logic;
signal \N__54435\ : std_logic;
signal \N__54432\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54428\ : std_logic;
signal \N__54427\ : std_logic;
signal \N__54424\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54421\ : std_logic;
signal \N__54420\ : std_logic;
signal \N__54419\ : std_logic;
signal \N__54418\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54386\ : std_logic;
signal \N__54379\ : std_logic;
signal \N__54370\ : std_logic;
signal \N__54363\ : std_logic;
signal \N__54354\ : std_logic;
signal \N__54347\ : std_logic;
signal \N__54338\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54336\ : std_logic;
signal \N__54335\ : std_logic;
signal \N__54334\ : std_logic;
signal \N__54333\ : std_logic;
signal \N__54332\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54330\ : std_logic;
signal \N__54329\ : std_logic;
signal \N__54328\ : std_logic;
signal \N__54327\ : std_logic;
signal \N__54326\ : std_logic;
signal \N__54325\ : std_logic;
signal \N__54324\ : std_logic;
signal \N__54323\ : std_logic;
signal \N__54322\ : std_logic;
signal \N__54321\ : std_logic;
signal \N__54320\ : std_logic;
signal \N__54319\ : std_logic;
signal \N__54318\ : std_logic;
signal \N__54317\ : std_logic;
signal \N__54316\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54314\ : std_logic;
signal \N__54313\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54311\ : std_logic;
signal \N__54310\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54307\ : std_logic;
signal \N__54304\ : std_logic;
signal \N__54289\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54259\ : std_logic;
signal \N__54244\ : std_logic;
signal \N__54243\ : std_logic;
signal \N__54240\ : std_logic;
signal \N__54239\ : std_logic;
signal \N__54236\ : std_logic;
signal \N__54235\ : std_logic;
signal \N__54232\ : std_logic;
signal \N__54231\ : std_logic;
signal \N__54230\ : std_logic;
signal \N__54227\ : std_logic;
signal \N__54226\ : std_logic;
signal \N__54223\ : std_logic;
signal \N__54222\ : std_logic;
signal \N__54219\ : std_logic;
signal \N__54218\ : std_logic;
signal \N__54199\ : std_logic;
signal \N__54192\ : std_logic;
signal \N__54183\ : std_logic;
signal \N__54176\ : std_logic;
signal \N__54167\ : std_logic;
signal \N__54160\ : std_logic;
signal \N__54151\ : std_logic;
signal \N__54150\ : std_logic;
signal \N__54147\ : std_logic;
signal \N__54146\ : std_logic;
signal \N__54143\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54139\ : std_logic;
signal \N__54138\ : std_logic;
signal \N__54137\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54135\ : std_logic;
signal \N__54134\ : std_logic;
signal \N__54133\ : std_logic;
signal \N__54132\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54124\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54103\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54073\ : std_logic;
signal \N__54058\ : std_logic;
signal \N__54043\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54027\ : std_logic;
signal \N__54026\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54024\ : std_logic;
signal \N__54023\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54021\ : std_logic;
signal \N__54020\ : std_logic;
signal \N__54015\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__54000\ : std_logic;
signal \N__53999\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53997\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53995\ : std_logic;
signal \N__53990\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53974\ : std_logic;
signal \N__53971\ : std_logic;
signal \N__53968\ : std_logic;
signal \N__53961\ : std_logic;
signal \N__53952\ : std_logic;
signal \N__53949\ : std_logic;
signal \N__53944\ : std_logic;
signal \N__53941\ : std_logic;
signal \N__53934\ : std_logic;
signal \N__53929\ : std_logic;
signal \N__53924\ : std_logic;
signal \N__53919\ : std_logic;
signal \N__53916\ : std_logic;
signal \N__53915\ : std_logic;
signal \N__53912\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53910\ : std_logic;
signal \N__53909\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53894\ : std_logic;
signal \N__53891\ : std_logic;
signal \N__53888\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53882\ : std_logic;
signal \N__53881\ : std_logic;
signal \N__53878\ : std_logic;
signal \N__53877\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53866\ : std_logic;
signal \N__53863\ : std_logic;
signal \N__53860\ : std_logic;
signal \N__53857\ : std_logic;
signal \N__53854\ : std_logic;
signal \N__53851\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53843\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53823\ : std_logic;
signal \N__53820\ : std_logic;
signal \N__53817\ : std_logic;
signal \N__53814\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53808\ : std_logic;
signal \N__53807\ : std_logic;
signal \N__53804\ : std_logic;
signal \N__53803\ : std_logic;
signal \N__53802\ : std_logic;
signal \N__53799\ : std_logic;
signal \N__53796\ : std_logic;
signal \N__53793\ : std_logic;
signal \N__53790\ : std_logic;
signal \N__53787\ : std_logic;
signal \N__53782\ : std_logic;
signal \N__53779\ : std_logic;
signal \N__53776\ : std_logic;
signal \N__53769\ : std_logic;
signal \N__53768\ : std_logic;
signal \N__53767\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53764\ : std_logic;
signal \N__53761\ : std_logic;
signal \N__53760\ : std_logic;
signal \N__53759\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53750\ : std_logic;
signal \N__53749\ : std_logic;
signal \N__53748\ : std_logic;
signal \N__53747\ : std_logic;
signal \N__53746\ : std_logic;
signal \N__53745\ : std_logic;
signal \N__53744\ : std_logic;
signal \N__53743\ : std_logic;
signal \N__53742\ : std_logic;
signal \N__53741\ : std_logic;
signal \N__53740\ : std_logic;
signal \N__53737\ : std_logic;
signal \N__53734\ : std_logic;
signal \N__53731\ : std_logic;
signal \N__53728\ : std_logic;
signal \N__53725\ : std_logic;
signal \N__53724\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53714\ : std_logic;
signal \N__53713\ : std_logic;
signal \N__53712\ : std_logic;
signal \N__53709\ : std_logic;
signal \N__53706\ : std_logic;
signal \N__53703\ : std_logic;
signal \N__53700\ : std_logic;
signal \N__53699\ : std_logic;
signal \N__53698\ : std_logic;
signal \N__53697\ : std_logic;
signal \N__53696\ : std_logic;
signal \N__53695\ : std_logic;
signal \N__53694\ : std_logic;
signal \N__53693\ : std_logic;
signal \N__53692\ : std_logic;
signal \N__53689\ : std_logic;
signal \N__53686\ : std_logic;
signal \N__53683\ : std_logic;
signal \N__53680\ : std_logic;
signal \N__53677\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53665\ : std_logic;
signal \N__53662\ : std_logic;
signal \N__53657\ : std_logic;
signal \N__53654\ : std_logic;
signal \N__53651\ : std_logic;
signal \N__53642\ : std_logic;
signal \N__53641\ : std_logic;
signal \N__53640\ : std_logic;
signal \N__53637\ : std_logic;
signal \N__53634\ : std_logic;
signal \N__53631\ : std_logic;
signal \N__53628\ : std_logic;
signal \N__53625\ : std_logic;
signal \N__53622\ : std_logic;
signal \N__53619\ : std_logic;
signal \N__53616\ : std_logic;
signal \N__53603\ : std_logic;
signal \N__53600\ : std_logic;
signal \N__53589\ : std_logic;
signal \N__53586\ : std_logic;
signal \N__53583\ : std_logic;
signal \N__53580\ : std_logic;
signal \N__53563\ : std_logic;
signal \N__53558\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53544\ : std_logic;
signal \N__53543\ : std_logic;
signal \N__53542\ : std_logic;
signal \N__53539\ : std_logic;
signal \N__53536\ : std_logic;
signal \N__53533\ : std_logic;
signal \N__53530\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53514\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53509\ : std_logic;
signal \N__53506\ : std_logic;
signal \N__53503\ : std_logic;
signal \N__53500\ : std_logic;
signal \N__53497\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53487\ : std_logic;
signal \N__53484\ : std_logic;
signal \N__53481\ : std_logic;
signal \N__53480\ : std_logic;
signal \N__53479\ : std_logic;
signal \N__53476\ : std_logic;
signal \N__53473\ : std_logic;
signal \N__53470\ : std_logic;
signal \N__53467\ : std_logic;
signal \N__53460\ : std_logic;
signal \N__53457\ : std_logic;
signal \N__53454\ : std_logic;
signal \N__53451\ : std_logic;
signal \N__53448\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53441\ : std_logic;
signal \N__53440\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53434\ : std_logic;
signal \N__53431\ : std_logic;
signal \N__53428\ : std_logic;
signal \N__53421\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53412\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53408\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53404\ : std_logic;
signal \N__53401\ : std_logic;
signal \N__53398\ : std_logic;
signal \N__53395\ : std_logic;
signal \N__53390\ : std_logic;
signal \N__53385\ : std_logic;
signal \N__53382\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53376\ : std_logic;
signal \N__53375\ : std_logic;
signal \N__53374\ : std_logic;
signal \N__53371\ : std_logic;
signal \N__53368\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53362\ : std_logic;
signal \N__53355\ : std_logic;
signal \N__53352\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53343\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53341\ : std_logic;
signal \N__53338\ : std_logic;
signal \N__53335\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53322\ : std_logic;
signal \N__53319\ : std_logic;
signal \N__53316\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53309\ : std_logic;
signal \N__53306\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53302\ : std_logic;
signal \N__53299\ : std_logic;
signal \N__53296\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53290\ : std_logic;
signal \N__53283\ : std_logic;
signal \N__53280\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53274\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53270\ : std_logic;
signal \N__53267\ : std_logic;
signal \N__53264\ : std_logic;
signal \N__53263\ : std_logic;
signal \N__53258\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53252\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53238\ : std_logic;
signal \N__53235\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53219\ : std_logic;
signal \N__53216\ : std_logic;
signal \N__53213\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53207\ : std_logic;
signal \N__53204\ : std_logic;
signal \N__53201\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53193\ : std_logic;
signal \N__53190\ : std_logic;
signal \N__53187\ : std_logic;
signal \N__53184\ : std_logic;
signal \N__53181\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53174\ : std_logic;
signal \N__53171\ : std_logic;
signal \N__53170\ : std_logic;
signal \N__53165\ : std_logic;
signal \N__53162\ : std_logic;
signal \N__53159\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53151\ : std_logic;
signal \N__53148\ : std_logic;
signal \N__53145\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53139\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53133\ : std_logic;
signal \N__53132\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53126\ : std_logic;
signal \N__53125\ : std_logic;
signal \N__53120\ : std_logic;
signal \N__53117\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53109\ : std_logic;
signal \N__53106\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53100\ : std_logic;
signal \N__53099\ : std_logic;
signal \N__53096\ : std_logic;
signal \N__53093\ : std_logic;
signal \N__53090\ : std_logic;
signal \N__53089\ : std_logic;
signal \N__53084\ : std_logic;
signal \N__53081\ : std_logic;
signal \N__53078\ : std_logic;
signal \N__53073\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53054\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53045\ : std_logic;
signal \N__53042\ : std_logic;
signal \N__53039\ : std_logic;
signal \N__53038\ : std_logic;
signal \N__53033\ : std_logic;
signal \N__53030\ : std_logic;
signal \N__53027\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53019\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53013\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53007\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52997\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52977\ : std_logic;
signal \N__52974\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52968\ : std_logic;
signal \N__52965\ : std_logic;
signal \N__52962\ : std_logic;
signal \N__52959\ : std_logic;
signal \N__52956\ : std_logic;
signal \N__52955\ : std_logic;
signal \N__52952\ : std_logic;
signal \N__52949\ : std_logic;
signal \N__52946\ : std_logic;
signal \N__52943\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52936\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52930\ : std_logic;
signal \N__52923\ : std_logic;
signal \N__52920\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52914\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52904\ : std_logic;
signal \N__52901\ : std_logic;
signal \N__52898\ : std_logic;
signal \N__52895\ : std_logic;
signal \N__52892\ : std_logic;
signal \N__52891\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52872\ : std_logic;
signal \N__52869\ : std_logic;
signal \N__52866\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52857\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52851\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52842\ : std_logic;
signal \N__52839\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52835\ : std_logic;
signal \N__52832\ : std_logic;
signal \N__52829\ : std_logic;
signal \N__52826\ : std_logic;
signal \N__52823\ : std_logic;
signal \N__52820\ : std_logic;
signal \N__52817\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52808\ : std_logic;
signal \N__52805\ : std_logic;
signal \N__52800\ : std_logic;
signal \N__52797\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52776\ : std_logic;
signal \N__52773\ : std_logic;
signal \N__52770\ : std_logic;
signal \N__52769\ : std_logic;
signal \N__52766\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52760\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52756\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52748\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52740\ : std_logic;
signal \N__52737\ : std_logic;
signal \N__52734\ : std_logic;
signal \N__52731\ : std_logic;
signal \N__52728\ : std_logic;
signal \N__52725\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52721\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52712\ : std_logic;
signal \N__52709\ : std_logic;
signal \N__52706\ : std_logic;
signal \N__52703\ : std_logic;
signal \N__52698\ : std_logic;
signal \N__52695\ : std_logic;
signal \N__52694\ : std_logic;
signal \N__52691\ : std_logic;
signal \N__52688\ : std_logic;
signal \N__52685\ : std_logic;
signal \N__52682\ : std_logic;
signal \N__52679\ : std_logic;
signal \N__52676\ : std_logic;
signal \N__52673\ : std_logic;
signal \N__52670\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52666\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52660\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52647\ : std_logic;
signal \N__52644\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52628\ : std_logic;
signal \N__52625\ : std_logic;
signal \N__52622\ : std_logic;
signal \N__52619\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52615\ : std_logic;
signal \N__52610\ : std_logic;
signal \N__52607\ : std_logic;
signal \N__52604\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52596\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52584\ : std_logic;
signal \N__52581\ : std_logic;
signal \N__52578\ : std_logic;
signal \N__52575\ : std_logic;
signal \N__52572\ : std_logic;
signal \N__52569\ : std_logic;
signal \N__52568\ : std_logic;
signal \N__52565\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52553\ : std_logic;
signal \N__52552\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52540\ : std_logic;
signal \N__52537\ : std_logic;
signal \N__52534\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52526\ : std_logic;
signal \N__52525\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52519\ : std_logic;
signal \N__52516\ : std_logic;
signal \N__52509\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52494\ : std_logic;
signal \N__52491\ : std_logic;
signal \N__52488\ : std_logic;
signal \N__52485\ : std_logic;
signal \N__52482\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52480\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52455\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52451\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52440\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52422\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52409\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52389\ : std_logic;
signal \N__52384\ : std_logic;
signal \N__52381\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52374\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52366\ : std_logic;
signal \N__52363\ : std_logic;
signal \N__52362\ : std_logic;
signal \N__52359\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52353\ : std_logic;
signal \N__52350\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52335\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52329\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52317\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52308\ : std_logic;
signal \N__52305\ : std_logic;
signal \N__52302\ : std_logic;
signal \N__52299\ : std_logic;
signal \N__52296\ : std_logic;
signal \N__52293\ : std_logic;
signal \N__52290\ : std_logic;
signal \N__52287\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52281\ : std_logic;
signal \N__52278\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52263\ : std_logic;
signal \N__52260\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52251\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52245\ : std_logic;
signal \N__52242\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52238\ : std_logic;
signal \N__52235\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52229\ : std_logic;
signal \N__52226\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52212\ : std_logic;
signal \N__52209\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52204\ : std_logic;
signal \N__52201\ : std_logic;
signal \N__52198\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52188\ : std_logic;
signal \N__52185\ : std_logic;
signal \N__52182\ : std_logic;
signal \N__52179\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52166\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52156\ : std_logic;
signal \N__52155\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52145\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52137\ : std_logic;
signal \N__52134\ : std_logic;
signal \N__52133\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52129\ : std_logic;
signal \N__52124\ : std_logic;
signal \N__52121\ : std_logic;
signal \N__52118\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52104\ : std_logic;
signal \N__52101\ : std_logic;
signal \N__52098\ : std_logic;
signal \N__52097\ : std_logic;
signal \N__52094\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52075\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52071\ : std_logic;
signal \N__52068\ : std_logic;
signal \N__52065\ : std_logic;
signal \N__52062\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52056\ : std_logic;
signal \N__52051\ : std_logic;
signal \N__52048\ : std_logic;
signal \N__52045\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52032\ : std_logic;
signal \N__52029\ : std_logic;
signal \N__52028\ : std_logic;
signal \N__52025\ : std_logic;
signal \N__52022\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52014\ : std_logic;
signal \N__52013\ : std_logic;
signal \N__52010\ : std_logic;
signal \N__52007\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51998\ : std_logic;
signal \N__51995\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51987\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51981\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51972\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51963\ : std_logic;
signal \N__51960\ : std_logic;
signal \N__51957\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51944\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51940\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51912\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51903\ : std_logic;
signal \N__51900\ : std_logic;
signal \N__51897\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51875\ : std_logic;
signal \N__51870\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51864\ : std_logic;
signal \N__51861\ : std_logic;
signal \N__51858\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51849\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51840\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51834\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51828\ : std_logic;
signal \N__51825\ : std_logic;
signal \N__51822\ : std_logic;
signal \N__51819\ : std_logic;
signal \N__51816\ : std_logic;
signal \N__51813\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51788\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51780\ : std_logic;
signal \N__51779\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51777\ : std_logic;
signal \N__51774\ : std_logic;
signal \N__51773\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51767\ : std_logic;
signal \N__51764\ : std_logic;
signal \N__51761\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51751\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51735\ : std_logic;
signal \N__51732\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51719\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51702\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51671\ : std_logic;
signal \N__51668\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51662\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51651\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51627\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51613\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51597\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51591\ : std_logic;
signal \N__51588\ : std_logic;
signal \N__51585\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51581\ : std_logic;
signal \N__51578\ : std_logic;
signal \N__51575\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51573\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51565\ : std_logic;
signal \N__51564\ : std_logic;
signal \N__51563\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51544\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51525\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51521\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51517\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51504\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51486\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51480\ : std_logic;
signal \N__51477\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51471\ : std_logic;
signal \N__51468\ : std_logic;
signal \N__51467\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51464\ : std_logic;
signal \N__51461\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51447\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51439\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51424\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51420\ : std_logic;
signal \N__51419\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51366\ : std_logic;
signal \N__51363\ : std_logic;
signal \N__51360\ : std_logic;
signal \N__51357\ : std_logic;
signal \N__51354\ : std_logic;
signal \N__51351\ : std_logic;
signal \N__51348\ : std_logic;
signal \N__51345\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51336\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51294\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51288\ : std_logic;
signal \N__51285\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51279\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51275\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51258\ : std_logic;
signal \N__51255\ : std_logic;
signal \N__51252\ : std_logic;
signal \N__51249\ : std_logic;
signal \N__51246\ : std_logic;
signal \N__51243\ : std_logic;
signal \N__51240\ : std_logic;
signal \N__51237\ : std_logic;
signal \N__51234\ : std_logic;
signal \N__51233\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51219\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51206\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51184\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51156\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51149\ : std_logic;
signal \N__51144\ : std_logic;
signal \N__51141\ : std_logic;
signal \N__51138\ : std_logic;
signal \N__51137\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51131\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51125\ : std_logic;
signal \N__51120\ : std_logic;
signal \N__51117\ : std_logic;
signal \N__51114\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51108\ : std_logic;
signal \N__51105\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51099\ : std_logic;
signal \N__51096\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51092\ : std_logic;
signal \N__51089\ : std_logic;
signal \N__51086\ : std_logic;
signal \N__51085\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51060\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51045\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51035\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51018\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51000\ : std_logic;
signal \N__50997\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50991\ : std_logic;
signal \N__50988\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50972\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50970\ : std_logic;
signal \N__50969\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50961\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50942\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50913\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50911\ : std_logic;
signal \N__50910\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50868\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50865\ : std_logic;
signal \N__50864\ : std_logic;
signal \N__50861\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50848\ : std_logic;
signal \N__50845\ : std_logic;
signal \N__50842\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50767\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50751\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50745\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50726\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50720\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50658\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50644\ : std_logic;
signal \N__50641\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50628\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50620\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50614\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50090\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50066\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50043\ : std_logic;
signal \N__50042\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49635\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49310\ : std_logic;
signal \N__49307\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49290\ : std_logic;
signal \N__49287\ : std_logic;
signal \N__49284\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49265\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49175\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48996\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48963\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48379\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48246\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47532\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44005\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal tx_enable : std_logic;
signal \LED_c\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \quad_counter0.n22_cascade_\ : std_logic;
signal \quad_counter0.n25_adj_4760_cascade_\ : std_logic;
signal \n12942_cascade_\ : std_logic;
signal \quad_counter0.n28_adj_4754\ : std_logic;
signal \quad_counter0.n26_adj_4755\ : std_logic;
signal \quad_counter0.n27_adj_4756_cascade_\ : std_logic;
signal \quad_counter0.n25_adj_4757\ : std_logic;
signal \n9809_cascade_\ : std_logic;
signal n9809 : std_logic;
signal \quad_counter1.n25_adj_4202_cascade_\ : std_logic;
signal n12940 : std_logic;
signal \PIN_13_c\ : std_logic;
signal \n12940_cascade_\ : std_logic;
signal \quadB_delayed_adj_4768\ : std_logic;
signal \n14425_cascade_\ : std_logic;
signal \quad_counter1.n26_adj_4200\ : std_logic;
signal b_delay_counter_0_adj_4766 : std_logic;
signal n187_adj_4771 : std_logic;
signal \bfn_5_17_0_\ : std_logic;
signal \quad_counter1.n19686\ : std_logic;
signal \quad_counter1.n19687\ : std_logic;
signal \quad_counter1.b_delay_counter_3\ : std_logic;
signal \quad_counter1.n19688\ : std_logic;
signal \quad_counter1.b_delay_counter_4\ : std_logic;
signal \quad_counter1.n19689\ : std_logic;
signal \quad_counter1.n19690\ : std_logic;
signal \quad_counter1.b_delay_counter_6\ : std_logic;
signal \quad_counter1.n19691\ : std_logic;
signal \quad_counter1.n19692\ : std_logic;
signal \quad_counter1.n19693\ : std_logic;
signal \quad_counter1.b_delay_counter_8\ : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal \quad_counter1.b_delay_counter_9\ : std_logic;
signal \quad_counter1.n19694\ : std_logic;
signal \quad_counter1.b_delay_counter_10\ : std_logic;
signal \quad_counter1.n19695\ : std_logic;
signal \quad_counter1.b_delay_counter_11\ : std_logic;
signal \quad_counter1.n19696\ : std_logic;
signal \quad_counter1.n19697\ : std_logic;
signal \quad_counter1.n19698\ : std_logic;
signal \quad_counter1.n19699\ : std_logic;
signal \quad_counter1.n19700\ : std_logic;
signal n14425 : std_logic;
signal \b_delay_counter_15__N_4140_adj_4773\ : std_logic;
signal b_delay_counter_0 : std_logic;
signal n187 : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \quad_counter0.b_delay_counter_1\ : std_logic;
signal \quad_counter0.n19656\ : std_logic;
signal \quad_counter0.b_delay_counter_2\ : std_logic;
signal \quad_counter0.n19657\ : std_logic;
signal \quad_counter0.b_delay_counter_3\ : std_logic;
signal \quad_counter0.n19658\ : std_logic;
signal \quad_counter0.b_delay_counter_4\ : std_logic;
signal \quad_counter0.n19659\ : std_logic;
signal \quad_counter0.n19660\ : std_logic;
signal \quad_counter0.b_delay_counter_6\ : std_logic;
signal \quad_counter0.n19661\ : std_logic;
signal \quad_counter0.n19662\ : std_logic;
signal \quad_counter0.n19663\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \quad_counter0.b_delay_counter_9\ : std_logic;
signal \quad_counter0.n19664\ : std_logic;
signal \quad_counter0.n19665\ : std_logic;
signal \quad_counter0.n19666\ : std_logic;
signal \quad_counter0.n19667\ : std_logic;
signal \quad_counter0.b_delay_counter_13\ : std_logic;
signal \quad_counter0.n19668\ : std_logic;
signal \quad_counter0.n19669\ : std_logic;
signal \quad_counter0.n19670\ : std_logic;
signal n14315 : std_logic;
signal \b_delay_counter_15__N_4140\ : std_logic;
signal \PIN_8_c\ : std_logic;
signal \quadB_delayed\ : std_logic;
signal n12942 : std_logic;
signal \quad_counter0.b_delay_counter_15\ : std_logic;
signal \quad_counter0.b_delay_counter_8\ : std_logic;
signal \quad_counter0.A_delayed\ : std_logic;
signal \quad_counter0.b_delay_counter_7\ : std_logic;
signal \quad_counter0.b_delay_counter_12\ : std_logic;
signal \quad_counter0.b_delay_counter_5\ : std_logic;
signal \quad_counter0.b_delay_counter_14\ : std_logic;
signal \quad_counter0.b_delay_counter_10\ : std_logic;
signal \quad_counter0.b_delay_counter_11\ : std_logic;
signal \quad_counter0.n24_adj_4758_cascade_\ : std_logic;
signal \quad_counter0.n18\ : std_logic;
signal \quad_counter0.n26_adj_4759\ : std_logic;
signal a_delay_counter_0 : std_logic;
signal n39 : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal \quad_counter0.a_delay_counter_1\ : std_logic;
signal \quad_counter0.n19671\ : std_logic;
signal \quad_counter0.a_delay_counter_2\ : std_logic;
signal \quad_counter0.n19672\ : std_logic;
signal \quad_counter0.a_delay_counter_3\ : std_logic;
signal \quad_counter0.n19673\ : std_logic;
signal \quad_counter0.a_delay_counter_4\ : std_logic;
signal \quad_counter0.n19674\ : std_logic;
signal \quad_counter0.a_delay_counter_5\ : std_logic;
signal \quad_counter0.n19675\ : std_logic;
signal \quad_counter0.a_delay_counter_6\ : std_logic;
signal \quad_counter0.n19676\ : std_logic;
signal \quad_counter0.a_delay_counter_7\ : std_logic;
signal \quad_counter0.n19677\ : std_logic;
signal \quad_counter0.n19678\ : std_logic;
signal \quad_counter0.a_delay_counter_8\ : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \quad_counter0.a_delay_counter_9\ : std_logic;
signal \quad_counter0.n19679\ : std_logic;
signal \quad_counter0.a_delay_counter_10\ : std_logic;
signal \quad_counter0.n19680\ : std_logic;
signal \quad_counter0.a_delay_counter_11\ : std_logic;
signal \quad_counter0.n19681\ : std_logic;
signal \quad_counter0.a_delay_counter_12\ : std_logic;
signal \quad_counter0.n19682\ : std_logic;
signal \quad_counter0.a_delay_counter_13\ : std_logic;
signal \quad_counter0.n19683\ : std_logic;
signal \quad_counter0.a_delay_counter_14\ : std_logic;
signal \quad_counter0.n19684\ : std_logic;
signal \quad_counter0.n19685\ : std_logic;
signal \quad_counter0.a_delay_counter_15\ : std_logic;
signal n14469 : std_logic;
signal \a_delay_counter_15__N_4123\ : std_logic;
signal \quad_counter1.b_delay_counter_13\ : std_logic;
signal \quad_counter1.b_delay_counter_1\ : std_logic;
signal \quad_counter1.b_delay_counter_2\ : std_logic;
signal \quad_counter1.b_delay_counter_5\ : std_logic;
signal \quad_counter1.n28_adj_4199\ : std_logic;
signal \PIN_7_c\ : std_logic;
signal \quadA_delayed\ : std_logic;
signal \quad_counter1.b_delay_counter_14\ : std_logic;
signal \quad_counter1.b_delay_counter_7\ : std_logic;
signal \quad_counter1.b_delay_counter_12\ : std_logic;
signal \quad_counter1.b_delay_counter_15\ : std_logic;
signal \quad_counter1.n27_adj_4201\ : std_logic;
signal \A_filtered\ : std_logic;
signal n8628 : std_logic;
signal \n9603_cascade_\ : std_logic;
signal \B_filtered\ : std_logic;
signal \quad_counter0.B_delayed\ : std_logic;
signal n10_adj_4777 : std_logic;
signal \c0.n25086_cascade_\ : std_logic;
signal data_out_frame_9_3 : std_logic;
signal \n24802_cascade_\ : std_logic;
signal \c0.n11_adj_4715_cascade_\ : std_logic;
signal n25010 : std_logic;
signal \c0.tx.n6_cascade_\ : std_logic;
signal \c0.n25089\ : std_logic;
signal n25018 : std_logic;
signal \c0.tx.n23980\ : std_logic;
signal \c0.n5_adj_4712_cascade_\ : std_logic;
signal \c0.n24800\ : std_logic;
signal \c0.tx.n5_adj_4207\ : std_logic;
signal \c0.n24949\ : std_logic;
signal \c0.n25104_cascade_\ : std_logic;
signal \c0.n25107\ : std_logic;
signal data_out_frame_5_7 : std_logic;
signal n25071 : std_logic;
signal \n3821_cascade_\ : std_logic;
signal data_out_frame_9_7 : std_logic;
signal \c0.rx.n24875\ : std_logic;
signal \c0.rx.n25068\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \quad_counter1.n19701\ : std_logic;
signal \quad_counter1.n19702\ : std_logic;
signal \quad_counter1.n19703\ : std_logic;
signal \quad_counter1.n19704\ : std_logic;
signal \quad_counter1.n19705\ : std_logic;
signal \quad_counter1.n19706\ : std_logic;
signal \quad_counter1.n19707\ : std_logic;
signal \quad_counter1.n19708\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \quad_counter1.n19709\ : std_logic;
signal \quad_counter1.n19710\ : std_logic;
signal \quad_counter1.n19711\ : std_logic;
signal \quad_counter1.n19712\ : std_logic;
signal \quad_counter1.n19713\ : std_logic;
signal \quad_counter1.n19714\ : std_logic;
signal \quad_counter1.n19715\ : std_logic;
signal \c0.tx.r_SM_Main_2\ : std_logic;
signal \r_SM_Main_2_N_3751_1\ : std_logic;
signal \c0.tx.n3843\ : std_logic;
signal \n3_cascade_\ : std_logic;
signal tx_o : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \c0.tx.n19492\ : std_logic;
signal \c0.tx.n22949\ : std_logic;
signal \c0.tx.n19492_cascade_\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \c0.tx.n25080\ : std_logic;
signal \c0.tx.n25083_cascade_\ : std_logic;
signal \c0.tx.o_Tx_Serial_N_3782\ : std_logic;
signal n10 : std_logic;
signal \c0.tx.r_Bit_Index_2\ : std_logic;
signal \c0.tx.n17832\ : std_logic;
signal \n10_adj_4776_cascade_\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \c0.tx.n25077\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \c0.tx.r_Bit_Index_0\ : std_logic;
signal \c0.tx.r_Bit_Index_1\ : std_logic;
signal \c0.tx.n25074\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \c0.n24960_cascade_\ : std_logic;
signal \c0.n24806_cascade_\ : std_logic;
signal n24757 : std_logic;
signal \c0.n26_adj_4645\ : std_logic;
signal n24808 : std_logic;
signal n10_adj_4779 : std_logic;
signal \c0.tx.n5_cascade_\ : std_logic;
signal \c0.tx.n17904\ : std_logic;
signal \c0.tx.n25051\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_1\ : std_logic;
signal \c0.tx.n19723\ : std_logic;
signal \c0.tx.r_Clock_Count_2\ : std_logic;
signal \c0.tx.n19724\ : std_logic;
signal \c0.tx.r_Clock_Count_3\ : std_logic;
signal \c0.tx.n19725\ : std_logic;
signal \c0.tx.r_Clock_Count_4\ : std_logic;
signal \c0.tx.n19726\ : std_logic;
signal \c0.tx.r_Clock_Count_5\ : std_logic;
signal \c0.tx.n19727\ : std_logic;
signal \c0.tx.r_Clock_Count_6\ : std_logic;
signal \c0.tx.n19728\ : std_logic;
signal \c0.tx.r_Clock_Count_7\ : std_logic;
signal \c0.tx.n19729\ : std_logic;
signal \c0.tx.n19730\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_8\ : std_logic;
signal \c0.tx.n17199\ : std_logic;
signal \c0.tx.n4\ : std_logic;
signal \c0.tx.n14290_cascade_\ : std_logic;
signal data_out_frame_6_7 : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal data_out_frame_5_2 : std_logic;
signal n17951 : std_logic;
signal \r_SM_Main_1_adj_4774\ : std_logic;
signal n25006 : std_logic;
signal \c0.n11_adj_4663\ : std_logic;
signal data_out_frame_5_1 : std_logic;
signal data_out_frame_13_3 : std_logic;
signal data_out_frame_8_7 : std_logic;
signal data_out_frame_12_6 : std_logic;
signal \c0.n5_adj_4334\ : std_logic;
signal \c0.n4_adj_4332\ : std_logic;
signal \c0.n26_adj_4662\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \c0.n19795\ : std_logic;
signal \c0.n19796\ : std_logic;
signal \c0.n19797\ : std_logic;
signal \c0.n19798\ : std_logic;
signal \c0.n19799\ : std_logic;
signal \c0.byte_transmit_counter_6\ : std_logic;
signal \c0.n19800\ : std_logic;
signal \c0.n19801\ : std_logic;
signal \c0.byte_transmit_counter_7\ : std_logic;
signal \c0.n21611\ : std_logic;
signal \c0.FRAME_MATCHER_state_13\ : std_logic;
signal \c0.n21573\ : std_logic;
signal \c0.n21581\ : std_logic;
signal \c0.n21575\ : std_logic;
signal \c0.FRAME_MATCHER_state_14\ : std_logic;
signal \c0.n21577\ : std_logic;
signal \n9806_cascade_\ : std_logic;
signal \PIN_12_c\ : std_logic;
signal \quadA_delayed_adj_4767\ : std_logic;
signal n9806 : std_logic;
signal n14345 : std_logic;
signal \a_delay_counter_15__N_4123_adj_4772\ : std_logic;
signal \n14345_cascade_\ : std_logic;
signal n39_adj_4770 : std_logic;
signal \quad_counter1.a_delay_counter_5\ : std_logic;
signal \quad_counter1.a_delay_counter_11\ : std_logic;
signal \quad_counter1.a_delay_counter_4\ : std_logic;
signal a_delay_counter_0_adj_4765 : std_logic;
signal \quad_counter1.n25\ : std_logic;
signal \quad_counter1.a_delay_counter_9\ : std_logic;
signal \quad_counter1.a_delay_counter_6\ : std_logic;
signal \quad_counter1.a_delay_counter_12\ : std_logic;
signal \quad_counter1.a_delay_counter_13\ : std_logic;
signal \quad_counter1.n26\ : std_logic;
signal \quad_counter1.a_delay_counter_8\ : std_logic;
signal \quad_counter1.a_delay_counter_1\ : std_logic;
signal \quad_counter1.a_delay_counter_2\ : std_logic;
signal \quad_counter1.a_delay_counter_3\ : std_logic;
signal \quad_counter1.n28\ : std_logic;
signal \quad_counter1.a_delay_counter_14\ : std_logic;
signal \quad_counter1.a_delay_counter_7\ : std_logic;
signal \quad_counter1.a_delay_counter_10\ : std_logic;
signal \quad_counter1.a_delay_counter_15\ : std_logic;
signal \quad_counter1.n27\ : std_logic;
signal \B_filtered_adj_4764\ : std_logic;
signal \quad_counter1.A_delayed\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \c0.n21391_cascade_\ : std_logic;
signal \c0.n21362_cascade_\ : std_logic;
signal \c0.n21244_cascade_\ : std_logic;
signal \c0.n22163\ : std_logic;
signal \c0.n6_adj_4297_cascade_\ : std_logic;
signal \c0.data_out_frame_28_4\ : std_logic;
signal \n26_cascade_\ : std_logic;
signal n25021 : std_logic;
signal n25022 : std_logic;
signal \c0.n24033_cascade_\ : std_logic;
signal \n21307_cascade_\ : std_logic;
signal \c0.n7_cascade_\ : std_logic;
signal \c0.n23918\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \c0.n20341_cascade_\ : std_logic;
signal data_out_frame_13_7 : std_logic;
signal data_out_frame_10_7 : std_logic;
signal n9603 : std_logic;
signal byte_transmit_counter_5 : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal data_out_frame_13_6 : std_logic;
signal data_out_frame_8_3 : std_logic;
signal n24796 : std_logic;
signal data_out_frame_7_7 : std_logic;
signal \n24805_cascade_\ : std_logic;
signal n10_adj_4780 : std_logic;
signal data_out_frame_11_5 : std_logic;
signal \c0.n25092_cascade_\ : std_logic;
signal \c0.n25095_cascade_\ : std_logic;
signal n25014 : std_logic;
signal data_out_frame_9_5 : std_logic;
signal n25008 : std_logic;
signal \c0.n11_adj_4681\ : std_logic;
signal \c0.n24897\ : std_logic;
signal data_out_frame_5_0 : std_logic;
signal data_out_frame_0_2 : std_logic;
signal data_out_frame_12_5 : std_logic;
signal \c0.n24900\ : std_logic;
signal \n14247_cascade_\ : std_logic;
signal data_out_frame_0_3 : std_logic;
signal \c0.n8_adj_4740_cascade_\ : std_logic;
signal \c0.n22952_cascade_\ : std_logic;
signal \c0.n14380\ : std_logic;
signal \c0.n14380_cascade_\ : std_logic;
signal \c0.n14942\ : std_logic;
signal \c0.n4728\ : std_logic;
signal \c0.n4728_cascade_\ : std_logic;
signal \c0.n58_adj_4742\ : std_logic;
signal \c0.n22952\ : std_logic;
signal \c0.r_SM_Main_2_N_3754_0\ : std_logic;
signal \c0.tx_active\ : std_logic;
signal \c0.n5_cascade_\ : std_logic;
signal \c0.n21585\ : std_logic;
signal \c0.n3\ : std_logic;
signal \c0.n21597\ : std_logic;
signal \c0.n21587\ : std_logic;
signal \c0.n10_adj_4303_cascade_\ : std_logic;
signal \c0.data_out_frame_29__7__N_849\ : std_logic;
signal \c0.n22246_cascade_\ : std_logic;
signal \c0.n22846\ : std_logic;
signal \c0.n20379_cascade_\ : std_logic;
signal \A_filtered_adj_4763\ : std_logic;
signal \quad_counter1.B_delayed\ : std_logic;
signal \c0.n6_adj_4456\ : std_logic;
signal \n21484_cascade_\ : std_logic;
signal \c0.n22246\ : std_logic;
signal data_out_frame_7_3 : std_logic;
signal \c0.n10_adj_4313\ : std_logic;
signal data_out_frame_11_3 : std_logic;
signal \c0.n22534\ : std_logic;
signal \c0.n22534_cascade_\ : std_logic;
signal \c0.n20415_cascade_\ : std_logic;
signal \c0.n20384\ : std_logic;
signal \c0.n22544\ : std_logic;
signal \c0.data_out_frame_28_5\ : std_logic;
signal \c0.n26_adj_4680\ : std_logic;
signal \c0.n22478\ : std_logic;
signal n22735 : std_logic;
signal \n22735_cascade_\ : std_logic;
signal \c0.n22757\ : std_logic;
signal \c0.n20_adj_4699_cascade_\ : std_logic;
signal n22285 : std_logic;
signal \c0.n6_adj_4210\ : std_logic;
signal \c0.n13683\ : std_logic;
signal data_out_frame_10_3 : std_logic;
signal \c0.n21362\ : std_logic;
signal \c0.n11_adj_4572\ : std_logic;
signal data_out_frame_13_0 : std_logic;
signal data_out_frame_6_2 : std_logic;
signal \c0.n5_adj_4650_cascade_\ : std_logic;
signal \c0.n6_adj_4649\ : std_logic;
signal \c0.n24953\ : std_logic;
signal \c0.n24803\ : std_logic;
signal data_out_frame_8_2 : std_logic;
signal \c0.n25059_cascade_\ : std_logic;
signal \n25004_cascade_\ : std_logic;
signal n10_adj_4778 : std_logic;
signal \c0.n24809\ : std_logic;
signal n24811 : std_logic;
signal n24904 : std_logic;
signal data_out_frame_28_3 : std_logic;
signal \c0.n25110_cascade_\ : std_logic;
signal \c0.n25113\ : std_logic;
signal \c0.n25056\ : std_logic;
signal data_out_frame_10_2 : std_logic;
signal data_out_frame_11_0 : std_logic;
signal \c0.n11_adj_4703\ : std_logic;
signal \c0.n24945_cascade_\ : std_logic;
signal n24682 : std_logic;
signal \c0.n24797_cascade_\ : std_logic;
signal byte_transmit_counter_4 : std_logic;
signal byte_transmit_counter_3 : std_logic;
signal \n24799_cascade_\ : std_logic;
signal n25012 : std_logic;
signal n10_adj_4775 : std_logic;
signal data_out_frame_11_6 : std_logic;
signal \c0.n25098_cascade_\ : std_logic;
signal \c0.n25101\ : std_logic;
signal data_out_frame_6_5 : std_logic;
signal data_out_frame_5_5 : std_logic;
signal \c0.n5_adj_4679\ : std_logic;
signal \c0.n25016_cascade_\ : std_logic;
signal \c0.n24794\ : std_logic;
signal \c0.n5_adj_4700\ : std_logic;
signal \c0.n24255\ : std_logic;
signal \c0.n21583\ : std_logic;
signal \c0.FRAME_MATCHER_state_26\ : std_logic;
signal \c0.FRAME_MATCHER_state_17\ : std_logic;
signal \c0.n14530_cascade_\ : std_logic;
signal \c0.rx.n9_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_30\ : std_logic;
signal \c0.rx.n17531_cascade_\ : std_logic;
signal \c0.rx.n17590\ : std_logic;
signal \c0.rx.n17848\ : std_logic;
signal \c0.rx.n14\ : std_logic;
signal \c0.rx.n24697_cascade_\ : std_logic;
signal \c0.rx.n24914_cascade_\ : std_logic;
signal \n14895_cascade_\ : std_logic;
signal \n24921_cascade_\ : std_logic;
signal n24922 : std_logic;
signal \c0.rx.n24916\ : std_logic;
signal \c0.rx.n8\ : std_logic;
signal \r_Clock_Count_0\ : std_logic;
signal n226 : std_logic;
signal \bfn_11_26_0_\ : std_logic;
signal \c0.rx.r_Clock_Count_1\ : std_logic;
signal \c0.rx.n19716\ : std_logic;
signal \c0.rx.r_Clock_Count_2\ : std_logic;
signal \c0.rx.n19717\ : std_logic;
signal \c0.rx.r_Clock_Count_3\ : std_logic;
signal \c0.rx.n19718\ : std_logic;
signal \c0.rx.r_Clock_Count_4\ : std_logic;
signal \c0.rx.n19719\ : std_logic;
signal \c0.rx.r_Clock_Count_5\ : std_logic;
signal \c0.rx.n19720\ : std_logic;
signal \c0.rx.r_Clock_Count_6\ : std_logic;
signal \c0.rx.n19721\ : std_logic;
signal \c0.rx.n19722\ : std_logic;
signal \c0.rx.r_Clock_Count_7\ : std_logic;
signal n14895 : std_logic;
signal \c0.n21645\ : std_logic;
signal \c0.n22638_cascade_\ : std_logic;
signal \c0.n21323_cascade_\ : std_logic;
signal \c0.n14_adj_4368\ : std_logic;
signal \c0.n12488_cascade_\ : std_logic;
signal \c0.n20379\ : std_logic;
signal \c0.n13531_cascade_\ : std_logic;
signal \c0.n22294\ : std_logic;
signal \c0.n13741\ : std_logic;
signal \c0.n14_adj_4317_cascade_\ : std_logic;
signal \c0.n15_adj_4318\ : std_logic;
signal \c0.n6_adj_4330\ : std_logic;
signal \c0.n20367\ : std_logic;
signal \c0.n6_adj_4336\ : std_logic;
signal \c0.n22531\ : std_logic;
signal n25065 : std_logic;
signal \c0.n13531\ : std_logic;
signal \c0.n20415\ : std_logic;
signal \c0.n22452\ : std_logic;
signal \c0.n9_adj_4562\ : std_logic;
signal \c0.n10_adj_4690_cascade_\ : std_logic;
signal \c0.n22710\ : std_logic;
signal \c0.n22710_cascade_\ : std_logic;
signal \c0.n12539\ : std_logic;
signal \c0.n21309\ : std_logic;
signal \c0.n6_adj_4683_cascade_\ : std_logic;
signal \c0.n13938\ : std_logic;
signal \c0.n12_adj_4688\ : std_logic;
signal \c0.n20360\ : std_logic;
signal \c0.n22668\ : std_logic;
signal \c0.n20360_cascade_\ : std_logic;
signal \c0.data_out_frame_29_7\ : std_logic;
signal \c0.n26_adj_4713\ : std_logic;
signal data_out_frame_7_0 : std_logic;
signal \c0.n5_adj_4567\ : std_logic;
signal data_out_frame_13_1 : std_logic;
signal \c0.n11_adj_4646\ : std_logic;
signal \c0.n5_adj_4644\ : std_logic;
signal \c0.n11_adj_4652\ : std_logic;
signal \c0.data_out_frame_28_2\ : std_logic;
signal \c0.n26_adj_4651\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \quad_counter1.count_direction\ : std_logic;
signal n2291 : std_logic;
signal \quad_counter1.n19731\ : std_logic;
signal n2290 : std_logic;
signal \quad_counter1.n19732\ : std_logic;
signal n2289 : std_logic;
signal \quad_counter1.n19733\ : std_logic;
signal n2288 : std_logic;
signal \quad_counter1.n19734\ : std_logic;
signal n2287 : std_logic;
signal \quad_counter1.n19735\ : std_logic;
signal n2286 : std_logic;
signal \quad_counter1.n19736\ : std_logic;
signal n2285 : std_logic;
signal \quad_counter1.n19737\ : std_logic;
signal \quad_counter1.n19738\ : std_logic;
signal n2284 : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \quad_counter1.n19739\ : std_logic;
signal n2282 : std_logic;
signal \quad_counter1.n19740\ : std_logic;
signal \quad_counter1.n19741\ : std_logic;
signal n2280 : std_logic;
signal \quad_counter1.n19742\ : std_logic;
signal n2279 : std_logic;
signal \quad_counter1.n19743\ : std_logic;
signal encoder1_position_13 : std_logic;
signal n2278 : std_logic;
signal \quad_counter1.n19744\ : std_logic;
signal n2277 : std_logic;
signal \quad_counter1.n19745\ : std_logic;
signal \quad_counter1.n19746\ : std_logic;
signal n2276 : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \quad_counter1.n19747\ : std_logic;
signal \quad_counter1.n19748\ : std_logic;
signal \quad_counter1.n19749\ : std_logic;
signal encoder1_position_19 : std_logic;
signal n2272 : std_logic;
signal \quad_counter1.n19750\ : std_logic;
signal n2271 : std_logic;
signal \quad_counter1.n19751\ : std_logic;
signal \quad_counter1.n19752\ : std_logic;
signal n2269 : std_logic;
signal \quad_counter1.n19753\ : std_logic;
signal \quad_counter1.n19754\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \quad_counter1.n19755\ : std_logic;
signal n2266 : std_logic;
signal \quad_counter1.n19756\ : std_logic;
signal \quad_counter1.n19757\ : std_logic;
signal \quad_counter1.n19758\ : std_logic;
signal \quad_counter1.n19759\ : std_logic;
signal \quad_counter1.n19760\ : std_logic;
signal \quad_counter1.n19761\ : std_logic;
signal \quad_counter1.n19762\ : std_logic;
signal \quad_counter1.n2226\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \c0.n24784_cascade_\ : std_logic;
signal n25019 : std_logic;
signal data_out_frame_11_2 : std_logic;
signal n2273 : std_logic;
signal encoder1_position_18 : std_logic;
signal n2275 : std_logic;
signal data_out_frame_10_0 : std_logic;
signal data_out_frame_10_4 : std_logic;
signal \c0.n24783\ : std_logic;
signal data_out_frame_6_0 : std_logic;
signal \c0.tx_transmit_N_3650\ : std_logic;
signal \c0.n24888\ : std_logic;
signal data_out_frame_12_0 : std_logic;
signal data_out_frame_12_1 : std_logic;
signal data_out_frame_9_6 : std_logic;
signal data_out_frame_6_6 : std_logic;
signal n14247 : std_logic;
signal data_out_frame_0_4 : std_logic;
signal data_out_frame_9_2 : std_logic;
signal data_out_frame_11_4 : std_logic;
signal data_out_frame_13_2 : std_logic;
signal \c0.n12976\ : std_logic;
signal \c0.n12976_cascade_\ : std_logic;
signal \c0.data_out_frame_29_7_N_1482_0_cascade_\ : std_logic;
signal \c0.n6_adj_4495\ : std_logic;
signal \c0.n14784\ : std_logic;
signal \c0.n9706_cascade_\ : std_logic;
signal \c0.n6_cascade_\ : std_logic;
signal \c0.n21579\ : std_logic;
signal \c0.n4_adj_4678\ : std_logic;
signal \c0.FRAME_MATCHER_state_28\ : std_logic;
signal \c0.n22131\ : std_logic;
signal \c0.FRAME_MATCHER_state_9\ : std_logic;
signal \c0.FRAME_MATCHER_state_5\ : std_logic;
signal \c0.n21625\ : std_logic;
signal \c0.n8_adj_4561\ : std_logic;
signal \c0.FRAME_MATCHER_state_8\ : std_logic;
signal \c0.n8_adj_4558\ : std_logic;
signal \c0.n21637\ : std_logic;
signal \c0.n22638\ : std_logic;
signal \c0.n22831_cascade_\ : std_logic;
signal \c0.n20_adj_4321\ : std_logic;
signal \c0.n13_adj_4320_cascade_\ : std_logic;
signal \c0.n14_adj_4319\ : std_logic;
signal \c0.n28_adj_4322_cascade_\ : std_logic;
signal \c0.n12488\ : std_logic;
signal encoder1_position_14 : std_logic;
signal \c0.n20318_cascade_\ : std_logic;
signal encoder1_position_16 : std_logic;
signal \c0.n20449\ : std_logic;
signal \c0.n10_adj_4374\ : std_logic;
signal \c0.data_out_frame_29__7__N_855\ : std_logic;
signal \c0.n13384\ : std_logic;
signal encoder1_position_0 : std_logic;
signal \c0.n22611\ : std_logic;
signal \c0.n10_adj_4274\ : std_logic;
signal \c0.n22791\ : std_logic;
signal \c0.n22466\ : std_logic;
signal \c0.n13121\ : std_logic;
signal \c0.n34_adj_4328\ : std_logic;
signal \c0.n30_adj_4326_cascade_\ : std_logic;
signal \c0.n29_adj_4329\ : std_logic;
signal encoder1_position_20 : std_logic;
signal \c0.n22788\ : std_logic;
signal \c0.n22788_cascade_\ : std_logic;
signal n2274 : std_logic;
signal n2283 : std_logic;
signal \c0.n22656\ : std_logic;
signal \c0.n22800\ : std_logic;
signal \c0.n10_adj_4339\ : std_logic;
signal \c0.n14_adj_4338_cascade_\ : std_logic;
signal \c0.n20461_cascade_\ : std_logic;
signal \c0.n20388\ : std_logic;
signal \c0.n22408\ : std_logic;
signal \c0.n22268\ : std_logic;
signal \c0.n5_adj_4660\ : std_logic;
signal \c0.n6_adj_4659\ : std_logic;
signal \c0.n24755\ : std_logic;
signal \c0.n22330\ : std_logic;
signal \c0.n19_adj_4693_cascade_\ : std_logic;
signal \c0.n6_adj_4691_cascade_\ : std_logic;
signal \c0.n21_adj_4692\ : std_logic;
signal \c0.n21457\ : std_logic;
signal \c0.n21489\ : std_logic;
signal encoder1_position_6 : std_logic;
signal \c0.n20461\ : std_logic;
signal \c0.n21330_cascade_\ : std_logic;
signal \c0.n6_adj_4331\ : std_logic;
signal \c0.n22414\ : std_logic;
signal n21307 : std_logic;
signal \c0.n6_adj_4215_cascade_\ : std_logic;
signal \c0.data_out_frame_29_0\ : std_logic;
signal \c0.data_out_frame_28_0\ : std_logic;
signal \c0.n26_adj_4570\ : std_logic;
signal \c0.n10529_cascade_\ : std_logic;
signal \c0.n22489_cascade_\ : std_logic;
signal \c0.n21416_cascade_\ : std_logic;
signal \c0.n24530\ : std_logic;
signal \c0.n22671_cascade_\ : std_logic;
signal \c0.n20230\ : std_logic;
signal \c0.n20230_cascade_\ : std_logic;
signal \c0.data_out_frame_29_5\ : std_logic;
signal data_out_frame_7_1 : std_logic;
signal n2270 : std_logic;
signal \c0.n13395\ : std_logic;
signal encoder1_position_1 : std_logic;
signal data_out_frame_9_0 : std_logic;
signal data_out_frame_5_4 : std_logic;
signal encoder1_position_22 : std_logic;
signal encoder1_position_7 : std_logic;
signal data_out_frame_7_2 : std_logic;
signal encoder1_position_11 : std_logic;
signal data_out_frame_12_3 : std_logic;
signal data_out_frame_12_2 : std_logic;
signal n2281 : std_logic;
signal encoder1_position_10 : std_logic;
signal data_out_frame_5_6 : std_logic;
signal encoder1_position_15 : std_logic;
signal data_out_frame_12_7 : std_logic;
signal n2263 : std_logic;
signal n2264 : std_logic;
signal encoder1_position_27 : std_logic;
signal data_out_frame_5_3 : std_logic;
signal n2262 : std_logic;
signal data_out_frame_10_6 : std_logic;
signal encoder1_position_4 : std_logic;
signal data_out_frame_8_0 : std_logic;
signal encoder1_position_17 : std_logic;
signal \c0.n16_adj_4233\ : std_logic;
signal data_out_frame_11_7 : std_logic;
signal data_out_frame_13_5 : std_logic;
signal data_out_frame_13_4 : std_logic;
signal \c0.n11_adj_4669\ : std_logic;
signal data_out_frame_8_5 : std_logic;
signal data_out_frame_7_5 : std_logic;
signal encoder1_position_25 : std_logic;
signal \c0.n7570_cascade_\ : std_logic;
signal data_out_frame_6_4 : std_logic;
signal data_out_frame_7_4 : std_logic;
signal \c0.n13055_cascade_\ : std_logic;
signal \n13058_cascade_\ : std_logic;
signal data_out_frame_7_6 : std_logic;
signal \c0.FRAME_MATCHER_state_3\ : std_logic;
signal \c0.n5_adj_4477\ : std_logic;
signal \c0.data_out_frame_29_7_N_1482_2\ : std_logic;
signal \c0.n14_adj_4727_cascade_\ : std_logic;
signal \c0.n13056\ : std_logic;
signal \c0.n63_adj_4235\ : std_logic;
signal \c0.n63_adj_4238\ : std_logic;
signal \c0.n2004_cascade_\ : std_logic;
signal \c0.n28_adj_4565\ : std_logic;
signal \c0.FRAME_MATCHER_state_16\ : std_logic;
signal \c0.n6_adj_4583\ : std_logic;
signal \c0.FRAME_MATCHER_state_6\ : std_logic;
signal \c0.n14_adj_4520\ : std_logic;
signal \c0.FRAME_MATCHER_state_4\ : std_logic;
signal \c0.n9_adj_4522\ : std_logic;
signal \c0.n20_adj_4265\ : std_logic;
signal \c0.n16919\ : std_logic;
signal \c0.n20_adj_4265_cascade_\ : std_logic;
signal \c0.n22148\ : std_logic;
signal \c0.n22145\ : std_logic;
signal \c0.n6_adj_4264\ : std_logic;
signal \c0.FRAME_MATCHER_state_22\ : std_logic;
signal \c0.n14721\ : std_logic;
signal \c0.n14530\ : std_logic;
signal \c0.n7_adj_4741\ : std_logic;
signal \c0.n9683\ : std_logic;
signal \c0.n9587\ : std_logic;
signal \c0.n9683_cascade_\ : std_logic;
signal \c0.n10\ : std_logic;
signal \c0.FRAME_MATCHER_state_25\ : std_logic;
signal \c0.n21653\ : std_logic;
signal \c0.FRAME_MATCHER_state_29\ : std_logic;
signal \c0.n21649\ : std_logic;
signal \c0.FRAME_MATCHER_state_24\ : std_logic;
signal \c0.n21595\ : std_logic;
signal \c0.n21643\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal encoder0_position_0 : std_logic;
signal \quad_counter0.count_direction\ : std_logic;
signal n2357 : std_logic;
signal \quad_counter0.n19763\ : std_logic;
signal encoder0_position_1 : std_logic;
signal n2356 : std_logic;
signal \quad_counter0.n19764\ : std_logic;
signal n2355 : std_logic;
signal \quad_counter0.n19765\ : std_logic;
signal n2354 : std_logic;
signal \quad_counter0.n19766\ : std_logic;
signal n2353 : std_logic;
signal \quad_counter0.n19767\ : std_logic;
signal \quad_counter0.n19768\ : std_logic;
signal n2351 : std_logic;
signal \quad_counter0.n19769\ : std_logic;
signal \quad_counter0.n19770\ : std_logic;
signal encoder0_position_7 : std_logic;
signal n2350 : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \quad_counter0.n19771\ : std_logic;
signal \quad_counter0.n19772\ : std_logic;
signal encoder0_position_10 : std_logic;
signal n2347 : std_logic;
signal \quad_counter0.n19773\ : std_logic;
signal encoder0_position_11 : std_logic;
signal n2346 : std_logic;
signal \quad_counter0.n19774\ : std_logic;
signal encoder0_position_12 : std_logic;
signal n2345 : std_logic;
signal \quad_counter0.n19775\ : std_logic;
signal \quad_counter0.n19776\ : std_logic;
signal \quad_counter0.n19777\ : std_logic;
signal \quad_counter0.n19778\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal encoder0_position_16 : std_logic;
signal n2341 : std_logic;
signal \quad_counter0.n19779\ : std_logic;
signal \quad_counter0.n19780\ : std_logic;
signal \quad_counter0.n19781\ : std_logic;
signal \quad_counter0.n19782\ : std_logic;
signal \quad_counter0.n19783\ : std_logic;
signal \quad_counter0.n19784\ : std_logic;
signal \quad_counter0.n19785\ : std_logic;
signal \quad_counter0.n19786\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal n2333 : std_logic;
signal \quad_counter0.n19787\ : std_logic;
signal n2332 : std_logic;
signal \quad_counter0.n19788\ : std_logic;
signal encoder0_position_26 : std_logic;
signal n2331 : std_logic;
signal \quad_counter0.n19789\ : std_logic;
signal n2330 : std_logic;
signal \quad_counter0.n19790\ : std_logic;
signal encoder0_position_28 : std_logic;
signal n2329 : std_logic;
signal \quad_counter0.n19791\ : std_logic;
signal encoder0_position_29 : std_logic;
signal n2328 : std_logic;
signal \quad_counter0.n19792\ : std_logic;
signal n2327 : std_logic;
signal \quad_counter0.n19793\ : std_logic;
signal \quad_counter0.n19794\ : std_logic;
signal \quad_counter0.n2313\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \n2326_cascade_\ : std_logic;
signal \c0.n22218\ : std_logic;
signal \c0.n21323\ : std_logic;
signal \c0.n22671\ : std_logic;
signal \c0.n20_adj_4694\ : std_logic;
signal \c0.n20348\ : std_logic;
signal \c0.n21330\ : std_logic;
signal \c0.n21355_cascade_\ : std_logic;
signal \c0.n12464\ : std_logic;
signal \c0.n20404\ : std_logic;
signal \c0.n20766\ : std_logic;
signal n2335 : std_logic;
signal \c0.n10427\ : std_logic;
signal \c0.n21360_cascade_\ : std_logic;
signal \c0.n10504\ : std_logic;
signal \c0.n22366\ : std_logic;
signal \c0.n10504_cascade_\ : std_logic;
signal \c0.n22327\ : std_logic;
signal n21484 : std_logic;
signal \c0.n28_adj_4698\ : std_logic;
signal \c0.n25_adj_4695_cascade_\ : std_logic;
signal \c0.data_out_frame_29_1\ : std_logic;
signal \c0.n22489\ : std_logic;
signal \c0.n21393\ : std_logic;
signal \c0.n22797\ : std_logic;
signal \c0.n26_adj_4697\ : std_logic;
signal \c0.n22475\ : std_logic;
signal \c0.data_out_frame_29__7__N_1143\ : std_logic;
signal \c0.n10_adj_4214\ : std_logic;
signal \c0.data_out_frame_28_1\ : std_logic;
signal \c0.n24033\ : std_logic;
signal \c0.n27_adj_4696\ : std_logic;
signal data_in_0_0 : std_logic;
signal data_in_0_4 : std_logic;
signal \c0.n15_adj_4242_cascade_\ : std_logic;
signal \c0.n22291\ : std_logic;
signal \c0.n20333\ : std_logic;
signal \c0.data_out_frame_29__7__N_1148\ : std_logic;
signal \c0.n21464\ : std_logic;
signal n2267 : std_logic;
signal encoder1_position_24 : std_logic;
signal \c0.n10_adj_4367\ : std_logic;
signal \c0.n10_adj_4239\ : std_logic;
signal \c0.n13049\ : std_logic;
signal data_in_2_4 : std_logic;
signal \c0.n13049_cascade_\ : std_logic;
signal \c0.n18_adj_4236_cascade_\ : std_logic;
signal \c0.n20_adj_4237\ : std_logic;
signal data_in_1_4 : std_logic;
signal \c0.n14_adj_4241\ : std_logic;
signal \c0.n17_adj_4234\ : std_logic;
signal n2268 : std_logic;
signal encoder1_position_23 : std_logic;
signal n2344 : std_logic;
signal \c0.n10_adj_4240\ : std_logic;
signal n14374 : std_logic;
signal \c0.tx.n24889\ : std_logic;
signal \c0.tx.r_Clock_Count_0\ : std_logic;
signal n2265 : std_logic;
signal encoder1_position_26 : std_logic;
signal data_out_frame_10_1 : std_logic;
signal data_out_frame_11_1 : std_logic;
signal \c0.n25116_cascade_\ : std_logic;
signal data_out_frame_9_1 : std_logic;
signal \c0.n25119\ : std_logic;
signal data_in_2_2 : std_logic;
signal data_out_frame_8_1 : std_logic;
signal encoder1_position_29 : std_logic;
signal data_out_frame_10_5 : std_logic;
signal \c0.n13046\ : std_logic;
signal \c0.n12898\ : std_logic;
signal \c0.n20_adj_4308_cascade_\ : std_logic;
signal \c0.n19_adj_4307\ : std_logic;
signal \c0.n16_adj_4231_cascade_\ : std_logic;
signal \c0.n12986\ : std_logic;
signal \c0.n24745\ : std_logic;
signal data_in_2_6 : std_logic;
signal data_in_0_5 : std_logic;
signal \c0.n17_adj_4232\ : std_logic;
signal n2261 : std_logic;
signal encoder1_position_30 : std_logic;
signal data_in_3_7 : std_logic;
signal data_in_3_5 : std_logic;
signal \c0.n13063\ : std_logic;
signal \c0.n13063_cascade_\ : std_logic;
signal \c0.n6_adj_4263\ : std_logic;
signal \c0.n9706\ : std_logic;
signal \c0.n3325\ : std_logic;
signal data_in_2_7 : std_logic;
signal data_in_1_7 : std_logic;
signal \c0.n17682\ : std_logic;
signal \c0.n1\ : std_logic;
signal \c0.n17846\ : std_logic;
signal \c0.n4_adj_4654\ : std_logic;
signal \c0.n17533\ : std_logic;
signal \c0.n22907\ : std_logic;
signal \c0.n24422\ : std_logic;
signal \c0.n24596_cascade_\ : std_logic;
signal \c0.n2004\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_3686_0\ : std_logic;
signal \c0.rx.n6_cascade_\ : std_logic;
signal n14439 : std_logic;
signal \c0.n7570\ : std_logic;
signal \c0.n24386\ : std_logic;
signal \c0.n24302_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_10\ : std_logic;
signal \c0.n8_adj_4556\ : std_logic;
signal \c0.FRAME_MATCHER_state_18\ : std_logic;
signal \c0.n21639\ : std_logic;
signal \c0.FRAME_MATCHER_state_12\ : std_logic;
signal \c0.n8_adj_4555\ : std_logic;
signal \c0.n21641\ : std_logic;
signal encoder0_position_30 : std_logic;
signal n2342 : std_logic;
signal encoder0_position_15 : std_logic;
signal n2352 : std_logic;
signal \c0.n30_adj_4730_cascade_\ : std_logic;
signal \c0.n17539\ : std_logic;
signal \c0.n22372\ : std_logic;
signal encoder1_position_28 : std_logic;
signal \c0.n31_adj_4325\ : std_logic;
signal \c0.n22775\ : std_logic;
signal n2348 : std_logic;
signal n2336 : std_logic;
signal \c0.n22608\ : std_logic;
signal encoder0_position_2 : std_logic;
signal \c0.n22785\ : std_logic;
signal \c0.n13630\ : std_logic;
signal n2340 : std_logic;
signal \c0.byte_transmit_counter_2\ : std_logic;
signal \c0.n5_adj_4217\ : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal \c0.n24901\ : std_logic;
signal \c0.n25062\ : std_logic;
signal n2260 : std_logic;
signal count_enable_adj_4769 : std_logic;
signal encoder1_position_31 : std_logic;
signal n2338 : std_logic;
signal encoder1_position_21 : std_logic;
signal encoder0_position_17 : std_logic;
signal encoder1_position_8 : std_logic;
signal \c0.n22593\ : std_logic;
signal encoder1_position_9 : std_logic;
signal \c0.n6_adj_4276\ : std_logic;
signal \c0.n21441\ : std_logic;
signal encoder0_position_25 : std_logic;
signal data_out_frame_6_1 : std_logic;
signal data_out_frame_29_2 : std_logic;
signal \c0.n12_adj_4312\ : std_logic;
signal \c0.n24113_cascade_\ : std_logic;
signal \c0.n10529\ : std_logic;
signal encoder1_position_5 : std_logic;
signal \c0.n21364\ : std_logic;
signal \c0.n24113\ : std_logic;
signal \c0.n21311_cascade_\ : std_logic;
signal \c0.n21244\ : std_logic;
signal \c0.n21496\ : std_logic;
signal \c0.n21273_cascade_\ : std_logic;
signal \c0.data_out_frame_29_6\ : std_logic;
signal \c0.data_out_frame_28_6\ : std_logic;
signal \c0.n26_adj_4702\ : std_logic;
signal \c0.n22617\ : std_logic;
signal \c0.n20341\ : std_logic;
signal \c0.n18_adj_4684_cascade_\ : std_logic;
signal \c0.n13268\ : std_logic;
signal \c0.n15_adj_4686\ : std_logic;
signal \c0.n20_adj_4685_cascade_\ : std_logic;
signal \c0.n21475\ : std_logic;
signal \c0.data_out_frame_28_7\ : std_logic;
signal \c0.n22461\ : std_logic;
signal \c0.n21358\ : std_logic;
signal \c0.n22461_cascade_\ : std_logic;
signal \c0.n21406\ : std_logic;
signal \c0.n24028\ : std_logic;
signal \c0.n14_adj_4478_cascade_\ : std_logic;
signal \c0.n22193\ : std_logic;
signal \c0.n13422\ : std_logic;
signal \c0.n22722\ : std_logic;
signal \data_out_frame_29__2__N_1748\ : std_logic;
signal \c0.n19_adj_4720\ : std_logic;
signal data_in_2_1 : std_logic;
signal data_out_frame_29_3 : std_logic;
signal encoder1_position_12 : std_logic;
signal data_out_frame_12_4 : std_logic;
signal data_in_0_3 : std_logic;
signal \c0.n15\ : std_logic;
signal data_in_3_4 : std_logic;
signal n2334 : std_logic;
signal data_in_1_0 : std_logic;
signal n2349 : std_logic;
signal \c0.rx.r_SM_Main_2_N_3680_2\ : std_logic;
signal encoder0_position_19 : std_logic;
signal \c0.n22199_cascade_\ : std_logic;
signal \c0.n22834\ : std_logic;
signal encoder0_position_13 : std_logic;
signal encoder0_position_22 : std_logic;
signal \c0.n6_adj_4366\ : std_logic;
signal data_in_2_0 : std_logic;
signal \c0.n22635\ : std_logic;
signal \c0.n22256_cascade_\ : std_logic;
signal \c0.n22772\ : std_logic;
signal data_in_1_3 : std_logic;
signal control_mode_4 : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal data_out_frame_9_4 : std_logic;
signal data_out_frame_8_4 : std_logic;
signal \c0.n24782\ : std_logic;
signal encoder0_position_8 : std_logic;
signal \c0.n22423\ : std_logic;
signal encoder0_position_6 : std_logic;
signal \c0.n6_adj_4293\ : std_logic;
signal encoder0_position_23 : std_logic;
signal encoder0_position_9 : std_logic;
signal control_mode_7 : std_logic;
signal \c0.n22385_cascade_\ : std_logic;
signal encoder0_position_24 : std_logic;
signal \c0.n20325\ : std_logic;
signal data_in_2_5 : std_logic;
signal data_in_1_5 : std_logic;
signal control_mode_6 : std_logic;
signal data_in_1_1 : std_logic;
signal data_in_0_1 : std_logic;
signal data_in_3_2 : std_logic;
signal \c0.n74_adj_4525\ : std_logic;
signal \c0.n4_adj_4212\ : std_logic;
signal \c0.n22098_cascade_\ : std_logic;
signal \c0.n4_adj_4306\ : std_logic;
signal \c0.n63_adj_4305_cascade_\ : std_logic;
signal \c0.n13001\ : std_logic;
signal \c0.FRAME_MATCHER_state_0\ : std_logic;
signal \c0.n9248\ : std_logic;
signal \c0.n13055\ : std_logic;
signal \c0.data_out_frame_29_7_N_1482_0\ : std_logic;
signal \data_out_frame_29_7_N_2878_2\ : std_logic;
signal \c0.n9_adj_4549\ : std_logic;
signal n63 : std_logic;
signal \c0.n3844\ : std_logic;
signal \c0.n58_adj_4706\ : std_logic;
signal \c0.n24591_cascade_\ : std_logic;
signal \c0.n6_adj_4728\ : std_logic;
signal \c0.FRAME_MATCHER_state_2\ : std_logic;
signal \c0.FRAME_MATCHER_state_15\ : std_logic;
signal \c0.n21659\ : std_logic;
signal \c0.n4_adj_4721\ : std_logic;
signal \c0.n937\ : std_logic;
signal \c0.data_out_frame_29_7_N_1482_1\ : std_logic;
signal \c0.FRAME_MATCHER_state_1\ : std_logic;
signal \c0.FRAME_MATCHER_state_20\ : std_logic;
signal \c0.n8_adj_4553\ : std_logic;
signal data_in_1_6 : std_logic;
signal data_in_0_6 : std_logic;
signal data_in_3_6 : std_logic;
signal \c0.n20_adj_4726\ : std_logic;
signal \c0.n27_adj_4735\ : std_logic;
signal \c0.data_out_frame_29__7__N_735\ : std_logic;
signal \c0.n13665\ : std_logic;
signal \c0.n22754\ : std_logic;
signal \c0.n13558\ : std_logic;
signal \c0.n22754_cascade_\ : std_logic;
signal \c0.n22243\ : std_logic;
signal \c0.n22580\ : std_logic;
signal \c0.n10477\ : std_logic;
signal n2339 : std_logic;
signal encoder0_position_18 : std_logic;
signal \c0.n22583\ : std_logic;
signal \c0.n22149\ : std_logic;
signal encoder0_position_3 : std_logic;
signal \c0.n22583_cascade_\ : std_logic;
signal encoder0_position_31 : std_logic;
signal \c0.n13872\ : std_logic;
signal n2337 : std_logic;
signal n17571 : std_logic;
signal encoder0_position_21 : std_logic;
signal \c0.n22252\ : std_logic;
signal encoder0_position_27 : std_logic;
signal data_out_frame_6_3 : std_logic;
signal encoder1_position_3 : std_logic;
signal \c0.n20455\ : std_logic;
signal encoder0_position_5 : std_logic;
signal encoder0_position_20 : std_logic;
signal \c0.n22689\ : std_logic;
signal \c0.n22641\ : std_logic;
signal encoder0_position_4 : std_logic;
signal \c0.n22689_cascade_\ : std_logic;
signal control_mode_0 : std_logic;
signal \c0.n10455\ : std_logic;
signal \c0.n20312\ : std_logic;
signal \c0.n20312_cascade_\ : std_logic;
signal \c0.n22522\ : std_logic;
signal \c0.n6_adj_4674_cascade_\ : std_logic;
signal \c0.data_out_frame_29_4\ : std_logic;
signal \c0.n8162\ : std_logic;
signal \c0.n21355\ : std_logic;
signal \c0.n12604\ : std_logic;
signal \c0.n20786\ : std_logic;
signal \c0.n20786_cascade_\ : std_logic;
signal \c0.n9_adj_4494\ : std_logic;
signal \c0.n10497\ : std_logic;
signal \c0.n21433\ : std_logic;
signal \c0.n21311\ : std_logic;
signal \c0.n12590\ : std_logic;
signal \c0.n21399\ : std_logic;
signal \c0.n22553\ : std_logic;
signal encoder1_position_2 : std_logic;
signal \c0.n21416\ : std_logic;
signal \c0.n10531\ : std_logic;
signal \c0.n20511\ : std_logic;
signal \c0.n10531_cascade_\ : std_logic;
signal \c0.n21451\ : std_logic;
signal \c0.n21437\ : std_logic;
signal \c0.n21451_cascade_\ : std_logic;
signal n13058 : std_logic;
signal data_out_frame_8_6 : std_logic;
signal \c0.n10467\ : std_logic;
signal \c0.n10500\ : std_logic;
signal \c0.n21349\ : std_logic;
signal \c0.n4_adj_4271\ : std_logic;
signal \c0.data_out_frame_29__6__N_1538\ : std_logic;
signal \c0.n21327\ : std_logic;
signal \c0.n4_adj_4271_cascade_\ : std_logic;
signal \c0.data_out_frame_29__3__N_1730\ : std_logic;
signal \data_out_frame_29__3__N_1661\ : std_logic;
signal \c0.rx.n12909\ : std_logic;
signal \c0.n22112_cascade_\ : std_logic;
signal data_in_2_3 : std_logic;
signal \c0.n82_cascade_\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \c0.rx.n17834_cascade_\ : std_logic;
signal n14484 : std_logic;
signal n14988 : std_logic;
signal control_mode_5 : std_logic;
signal control_mode_1 : std_logic;
signal control_mode_3 : std_logic;
signal count_enable : std_logic;
signal n2343 : std_logic;
signal encoder0_position_14 : std_logic;
signal n4_adj_4761 : std_logic;
signal \c0.data_in_frame_29_3\ : std_logic;
signal \c0.n17_adj_4483\ : std_logic;
signal \c0.n26_adj_4480_cascade_\ : std_logic;
signal \c0.n63_adj_4249\ : std_logic;
signal \c0.n34_adj_4546_cascade_\ : std_logic;
signal n24622 : std_logic;
signal \n24622_cascade_\ : std_logic;
signal control_mode_2 : std_logic;
signal \c0.n24539\ : std_logic;
signal \c0.n24733\ : std_logic;
signal \c0.n18_adj_4485\ : std_logic;
signal \c0.n22134_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_11\ : std_logic;
signal \c0.n21633\ : std_logic;
signal \c0.n6\ : std_logic;
signal \c0.n4_adj_4266\ : std_logic;
signal \c0.n5024\ : std_logic;
signal \c0.n12992\ : std_logic;
signal \c0.n13052\ : std_logic;
signal \c0.n24736\ : std_logic;
signal \c0.FRAME_MATCHER_state_31\ : std_logic;
signal \c0.n21651\ : std_logic;
signal \FRAME_MATCHER_state_31_N_2975_2\ : std_logic;
signal \c0.n22_adj_4643_cascade_\ : std_logic;
signal \c0.n10_adj_4639_cascade_\ : std_logic;
signal \c0.n13_adj_4640\ : std_logic;
signal \c0.n20_adj_4642\ : std_logic;
signal \c0.n14_adj_4607_cascade_\ : std_logic;
signal \c0.n22626\ : std_logic;
signal \c0.data_out_frame_0__7__N_2626_cascade_\ : std_logic;
signal \c0.n30_adj_4585\ : std_logic;
signal \c0.n6_adj_4254_cascade_\ : std_logic;
signal \c0.n28_adj_4731\ : std_logic;
signal data_in_3_3 : std_logic;
signal data_in_0_7 : std_logic;
signal \c0.n14\ : std_logic;
signal \c0.n20_adj_4729\ : std_logic;
signal \c0.n6_adj_4704\ : std_logic;
signal \c0.n14016_cascade_\ : std_logic;
signal \c0.n20_cascade_\ : std_logic;
signal data_in_frame_5_6 : std_logic;
signal \c0.data_in_frame_7_7\ : std_logic;
signal \c0.FRAME_MATCHER_state_7\ : std_logic;
signal \c0.n21629\ : std_logic;
signal \c0.n25_adj_4723\ : std_logic;
signal \c0.FRAME_MATCHER_state_19\ : std_logic;
signal \c0.FRAME_MATCHER_state_23\ : std_logic;
signal \c0.FRAME_MATCHER_state_21\ : std_logic;
signal \c0.n22049\ : std_logic;
signal \c0.n5\ : std_logic;
signal \c0.FRAME_MATCHER_state_27\ : std_logic;
signal \c0.n21647\ : std_logic;
signal data_in_1_2 : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.n10_adj_4732\ : std_logic;
signal \c0.n26_adj_4733_cascade_\ : std_logic;
signal \c0.n20409_cascade_\ : std_logic;
signal \c0.n22716_cascade_\ : std_logic;
signal \c0.n8_adj_4248\ : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_3_0 : std_logic;
signal n12981 : std_logic;
signal n4_adj_4762 : std_logic;
signal \c0.n22716\ : std_logic;
signal \c0.n5_adj_4302\ : std_logic;
signal \c0.n12_adj_4348_cascade_\ : std_logic;
signal \c0.n8_adj_4526\ : std_logic;
signal \c0.n8_adj_4526_cascade_\ : std_logic;
signal \c0.n9_adj_4536\ : std_logic;
signal \c0.n14_adj_4528\ : std_logic;
signal \c0.n14_adj_4576\ : std_logic;
signal \c0.data_in_frame_29_5\ : std_logic;
signal \c0.n24098_cascade_\ : std_logic;
signal \c0.n10_adj_4484\ : std_logic;
signal \c0.n52_cascade_\ : std_logic;
signal \c0.n47_adj_4537_cascade_\ : std_logic;
signal \c0.n24581\ : std_logic;
signal \c0.data_in_frame_29_1\ : std_logic;
signal \c0.data_in_frame_29_6\ : std_logic;
signal \c0.n20793\ : std_logic;
signal \c0.n20793_cascade_\ : std_logic;
signal \c0.n12927\ : std_logic;
signal \c0.n39_adj_4295\ : std_logic;
signal \c0.n13043\ : std_logic;
signal \c0.n23912\ : std_logic;
signal \c0.n35\ : std_logic;
signal \c0.n22885\ : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal n4 : std_logic;
signal \r_Rx_Data\ : std_logic;
signal \n4_cascade_\ : std_logic;
signal n12904 : std_logic;
signal \c0.rx.n14277\ : std_logic;
signal \c0.n12514\ : std_logic;
signal \c0.n20641\ : std_logic;
signal \c0.n21391\ : std_logic;
signal \c0.n21360\ : std_logic;
signal \c0.n21_adj_4719\ : std_logic;
signal rx_data_ready : std_logic;
signal \c0.FRAME_MATCHER_rx_data_ready_prev\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \c0.rx.r_SM_Main_0\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \c0.rx.n22094\ : std_logic;
signal \c0.n46_adj_4739\ : std_logic;
signal \c0.n39_adj_4737\ : std_logic;
signal \c0.n38_adj_4736\ : std_logic;
signal \c0.n23562\ : std_logic;
signal \c0.n23562_cascade_\ : std_logic;
signal data_in_frame_5_5 : std_logic;
signal \c0.data_in_frame_3_4\ : std_logic;
signal \c0.n12_adj_4657\ : std_logic;
signal \c0.n23_adj_4648\ : std_logic;
signal \c0.n38_adj_4285_cascade_\ : std_logic;
signal \c0.n26_adj_4289\ : std_logic;
signal \c0.n26_adj_4289_cascade_\ : std_logic;
signal \c0.data_out_frame_0__7__N_2626\ : std_logic;
signal \c0.n20_adj_4290\ : std_logic;
signal \c0.n20_adj_4290_cascade_\ : std_logic;
signal data_in_frame_1_1 : std_logic;
signal \c0.n51\ : std_logic;
signal \c0.n29\ : std_logic;
signal \c0.n51_cascade_\ : std_logic;
signal \c0.n22_adj_4647\ : std_logic;
signal \c0.n102_cascade_\ : std_logic;
signal \c0.n32\ : std_logic;
signal \c0.n16_adj_4256_cascade_\ : std_logic;
signal \c0.n9_adj_4279\ : std_logic;
signal \c0.n13141\ : std_logic;
signal \c0.n9_adj_4279_cascade_\ : std_logic;
signal \c0.n23574_cascade_\ : std_logic;
signal \c0.n11_adj_4257\ : std_logic;
signal \c0.n7_adj_4337\ : std_logic;
signal \c0.n38_adj_4573_cascade_\ : std_logic;
signal \c0.n44_adj_4744\ : std_logic;
signal \c0.n43_adj_4574_cascade_\ : std_logic;
signal \c0.n41_adj_4745\ : std_logic;
signal \c0.n24048\ : std_logic;
signal \c0.n24048_cascade_\ : std_logic;
signal \c0.n109\ : std_logic;
signal \c0.n23_adj_4590\ : std_logic;
signal \c0.n29_adj_4734\ : std_logic;
signal \c0.n7_adj_4221\ : std_logic;
signal \c0.n16_adj_4641\ : std_logic;
signal \c0.n23116_cascade_\ : std_logic;
signal \c0.n23116\ : std_logic;
signal \c0.n128\ : std_logic;
signal \c0.n129_cascade_\ : std_logic;
signal \c0.n11_adj_4614\ : std_logic;
signal \c0.n16_adj_4613_cascade_\ : std_logic;
signal data_in_frame_1_3 : std_logic;
signal \c0.n126\ : std_logic;
signal \c0.n123\ : std_logic;
signal \c0.n144_cascade_\ : std_logic;
signal \c0.n154\ : std_logic;
signal \c0.n15_adj_4301\ : std_logic;
signal \c0.n21_adj_4605\ : std_logic;
signal \c0.n19_adj_4604\ : std_logic;
signal \c0.n16_adj_4256\ : std_logic;
signal \c0.n22\ : std_logic;
signal \c0.n13280\ : std_logic;
signal \c0.n13_cascade_\ : std_logic;
signal \c0.n20_adj_4222\ : std_logic;
signal \c0.data_in_frame_3_5\ : std_logic;
signal \c0.n22_adj_4223_cascade_\ : std_logic;
signal \c0.n21_adj_4225_cascade_\ : std_logic;
signal \c0.n10_adj_4277_cascade_\ : std_logic;
signal \c0.n10_adj_4591_cascade_\ : std_logic;
signal \c0.n10_adj_4591\ : std_logic;
signal data_in_frame_21_2 : std_logic;
signal \c0.n12_adj_4606_cascade_\ : std_logic;
signal \c0.n21325_cascade_\ : std_logic;
signal \c0.n24384\ : std_logic;
signal \c0.n4_adj_4464_cascade_\ : std_logic;
signal \c0.n21428_cascade_\ : std_logic;
signal \c0.n24_adj_4593\ : std_logic;
signal \c0.n23_adj_4598\ : std_logic;
signal \c0.n4_adj_4352\ : std_logic;
signal \c0.n23_adj_4353\ : std_logic;
signal \c0.n23_adj_4353_cascade_\ : std_logic;
signal \c0.n15_adj_4344\ : std_logic;
signal \c0.n21428\ : std_logic;
signal \c0.n11_adj_4438_cascade_\ : std_logic;
signal \c0.n16_adj_4437\ : std_logic;
signal \c0.n22420\ : std_logic;
signal \c0.data_in_frame_28_0\ : std_logic;
signal \c0.n21491\ : std_logic;
signal \c0.n23187_cascade_\ : std_logic;
signal \c0.n10_adj_4439_cascade_\ : std_logic;
signal \c0.n20_adj_4441\ : std_logic;
signal \c0.n13_adj_4442_cascade_\ : std_logic;
signal \c0.n24528_cascade_\ : std_logic;
signal \c0.n23718\ : std_logic;
signal \c0.n12_adj_4506\ : std_logic;
signal \c0.n20_adj_4512\ : std_logic;
signal \c0.n24_adj_4509\ : std_logic;
signal \c0.n22_adj_4507\ : std_logic;
signal \c0.n23627\ : std_logic;
signal \c0.n23627_cascade_\ : std_logic;
signal \c0.n24528\ : std_logic;
signal \c0.n10_adj_4575\ : std_logic;
signal \c0.data_in_frame_24_7\ : std_logic;
signal \c0.n25467\ : std_logic;
signal \c0.n24098\ : std_logic;
signal \c0.data_in_frame_29_4\ : std_logic;
signal \c0.n23533\ : std_logic;
signal \c0.n5_adj_4370\ : std_logic;
signal \c0.n10_adj_4371\ : std_logic;
signal \c0.n5_adj_4349\ : std_logic;
signal \c0.n10_adj_4371_cascade_\ : std_logic;
signal \c0.n12_adj_4372\ : std_logic;
signal \c0.n12_adj_4671_cascade_\ : std_logic;
signal \c0.data_in_frame_28_7\ : std_logic;
signal \c0.n45_adj_4298\ : std_logic;
signal \c0.data_in_frame_25_3\ : std_logic;
signal \c0.data_in_frame_25_2\ : std_logic;
signal \c0.n40_adj_4294\ : std_logic;
signal \c0.n41_adj_4292\ : std_logic;
signal \c0.n42_adj_4272_cascade_\ : std_logic;
signal \c0.n44_adj_4270\ : std_logic;
signal \c0.n50_adj_4296\ : std_logic;
signal \c0.n43_adj_4275\ : std_logic;
signal \c0.n161\ : std_logic;
signal \bfn_19_1_0_\ : std_logic;
signal \c0.n19625\ : std_logic;
signal \c0.n19625_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19625_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19625_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19625_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19625_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19625_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19625_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_2_0_\ : std_logic;
signal \c0.n3_adj_4434\ : std_logic;
signal \c0.n19626\ : std_logic;
signal \c0.n19626_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19626_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19626_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19626_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19626_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19626_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19626_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_3_0_\ : std_logic;
signal \c0.n3_adj_4432\ : std_logic;
signal \c0.n19627\ : std_logic;
signal \c0.n19627_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19627_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19627_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19627_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19627_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19627_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19627_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_4_0_\ : std_logic;
signal \c0.n19628\ : std_logic;
signal \c0.n19628_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19628_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19628_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19628_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19628_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19628_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19628_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_4\ : std_logic;
signal \bfn_19_5_0_\ : std_logic;
signal \c0.n3_adj_4428\ : std_logic;
signal \c0.n19629\ : std_logic;
signal \c0.n19629_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19629_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19629_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19629_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19629_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19629_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19629_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_5\ : std_logic;
signal \bfn_19_6_0_\ : std_logic;
signal \c0.n3_adj_4426\ : std_logic;
signal \c0.n19630\ : std_logic;
signal \c0.n19630_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19630_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19630_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19630_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19630_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19630_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19630_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_6\ : std_logic;
signal \bfn_19_7_0_\ : std_logic;
signal \c0.n3_adj_4424\ : std_logic;
signal \c0.n19631\ : std_logic;
signal \c0.n19631_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19631_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19631_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19631_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19631_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19631_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19631_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_7\ : std_logic;
signal \bfn_19_8_0_\ : std_logic;
signal \c0.n3_adj_4422\ : std_logic;
signal \c0.n19632\ : std_logic;
signal \c0.n19632_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19632_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19632_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19632_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19632_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19632_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19632_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_8\ : std_logic;
signal \bfn_19_9_0_\ : std_logic;
signal \c0.n3_adj_4420\ : std_logic;
signal \c0.n19633\ : std_logic;
signal \c0.n19633_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19633_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19633_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19633_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19633_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19633_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19633_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_9\ : std_logic;
signal \bfn_19_10_0_\ : std_logic;
signal \c0.n3_adj_4418\ : std_logic;
signal \c0.n19634\ : std_logic;
signal \c0.n19634_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19634_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19634_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19634_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19634_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19634_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19634_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_10\ : std_logic;
signal \bfn_19_11_0_\ : std_logic;
signal \c0.n3_adj_4416\ : std_logic;
signal \c0.n19635\ : std_logic;
signal \c0.n19635_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19635_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19635_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19635_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19635_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19635_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19635_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_11\ : std_logic;
signal \bfn_19_12_0_\ : std_logic;
signal \c0.n3_adj_4414\ : std_logic;
signal \c0.n19636\ : std_logic;
signal \c0.n19636_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19636_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19636_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19636_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19636_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19636_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19636_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_12\ : std_logic;
signal \bfn_19_13_0_\ : std_logic;
signal \c0.n3_adj_4412\ : std_logic;
signal \c0.n19637\ : std_logic;
signal \c0.n19637_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19637_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19637_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19637_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19637_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19637_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19637_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_14_0_\ : std_logic;
signal \c0.n19638\ : std_logic;
signal \c0.n19638_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19638_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19638_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19638_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19638_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19638_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19638_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_14\ : std_logic;
signal \bfn_19_15_0_\ : std_logic;
signal \c0.n3_adj_4408\ : std_logic;
signal \c0.n19639\ : std_logic;
signal \c0.n19639_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19639_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19639_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19639_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19639_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19639_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19639_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_15\ : std_logic;
signal \bfn_19_16_0_\ : std_logic;
signal \c0.n3_adj_4406\ : std_logic;
signal \c0.n19640\ : std_logic;
signal \c0.n19640_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19640_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19640_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19640_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19640_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19640_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19640_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_16\ : std_logic;
signal \bfn_19_17_0_\ : std_logic;
signal \c0.n3_adj_4404\ : std_logic;
signal \c0.n19641\ : std_logic;
signal \c0.n19641_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19641_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19641_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19641_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19641_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19641_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19641_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_17\ : std_logic;
signal \bfn_19_18_0_\ : std_logic;
signal \c0.n3_adj_4402\ : std_logic;
signal \c0.n19642\ : std_logic;
signal \c0.n19642_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19642_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19642_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19642_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19642_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19642_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19642_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_19_0_\ : std_logic;
signal \c0.n19643\ : std_logic;
signal \c0.n19643_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19643_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19643_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19643_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19643_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19643_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19643_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_19\ : std_logic;
signal \bfn_19_20_0_\ : std_logic;
signal \c0.n3_adj_4398\ : std_logic;
signal \c0.n19644\ : std_logic;
signal \c0.n19644_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19644_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19644_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19644_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19644_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19644_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19644_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_20\ : std_logic;
signal \bfn_19_21_0_\ : std_logic;
signal \c0.n3_adj_4396\ : std_logic;
signal \c0.n19645\ : std_logic;
signal \c0.n19645_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19645_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19645_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19645_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19645_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19645_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19645_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_21\ : std_logic;
signal \bfn_19_22_0_\ : std_logic;
signal \c0.n3_adj_4394\ : std_logic;
signal \c0.n19646\ : std_logic;
signal \c0.n19646_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19646_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19646_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19646_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19646_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19646_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19646_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_22\ : std_logic;
signal \bfn_19_23_0_\ : std_logic;
signal \c0.n3_adj_4392\ : std_logic;
signal \c0.n19647\ : std_logic;
signal \c0.n19647_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19647_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19647_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19647_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19647_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19647_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19647_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_23\ : std_logic;
signal \bfn_19_24_0_\ : std_logic;
signal \c0.n3_adj_4390\ : std_logic;
signal \c0.n19648\ : std_logic;
signal \c0.n19648_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19648_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19648_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19648_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19648_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19648_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19648_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_24\ : std_logic;
signal \bfn_19_25_0_\ : std_logic;
signal \c0.n3_adj_4388\ : std_logic;
signal \c0.n19649\ : std_logic;
signal \c0.n19649_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19649_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19649_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19649_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19649_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19649_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19649_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_25\ : std_logic;
signal \bfn_19_26_0_\ : std_logic;
signal \c0.n3_adj_4386\ : std_logic;
signal \c0.n19650\ : std_logic;
signal \c0.n19650_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19650_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19650_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19650_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19650_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19650_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19650_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_26\ : std_logic;
signal \bfn_19_27_0_\ : std_logic;
signal \c0.n3_adj_4384\ : std_logic;
signal \c0.n19651\ : std_logic;
signal \c0.n19651_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19651_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19651_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19651_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19651_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19651_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19651_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_27\ : std_logic;
signal \bfn_19_28_0_\ : std_logic;
signal \c0.n3_adj_4382\ : std_logic;
signal \c0.n19652\ : std_logic;
signal \c0.n19652_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19652_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19652_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19652_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19652_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19652_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19652_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_28\ : std_logic;
signal \bfn_19_29_0_\ : std_logic;
signal \c0.n3_adj_4380\ : std_logic;
signal \c0.n19653\ : std_logic;
signal \c0.n19653_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19653_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19653_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19653_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19653_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19653_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19653_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_29\ : std_logic;
signal \bfn_19_30_0_\ : std_logic;
signal \c0.n3_adj_4378\ : std_logic;
signal \c0.n19654\ : std_logic;
signal \c0.n19654_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19654_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19654_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19654_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19654_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19654_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19654_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_30\ : std_logic;
signal \bfn_19_31_0_\ : std_logic;
signal \c0.n3_adj_4376\ : std_logic;
signal \c0.n19655\ : std_logic;
signal \c0.n19655_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19655_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19655_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19655_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19655_THRU_CRY_4_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.n19655_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19655_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_32_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31\ : std_logic;
signal \c0.n3_adj_4373\ : std_logic;
signal \c0.n17856\ : std_logic;
signal \c0.n1306\ : std_logic;
signal \c0.n3_adj_4436\ : std_logic;
signal \c0.n22196_cascade_\ : std_logic;
signal \c0.n12_adj_4258\ : std_logic;
signal \c0.data_in_frame_3_0\ : std_logic;
signal \c0.n10_adj_4615\ : std_logic;
signal \c0.data_in_frame_3_1\ : std_logic;
signal \c0.n7_adj_4300\ : std_logic;
signal \c0.n12_adj_4299\ : std_logic;
signal \c0.n7_adj_4300_cascade_\ : std_logic;
signal \c0.n11_adj_4280\ : std_logic;
signal \c0.n23251\ : std_logic;
signal \c0.n23305\ : std_logic;
signal \c0.n23251_cascade_\ : std_logic;
signal \c0.n23574\ : std_logic;
signal \c0.n7_adj_4282_cascade_\ : std_logic;
signal \c0.n10_adj_4283\ : std_logic;
signal \c0.data_in_frame_8_1\ : std_logic;
signal \c0.n13_adj_4638_cascade_\ : std_logic;
signal \c0.data_in_frame_10_1\ : std_logic;
signal \c0.data_in_frame_10_2\ : std_logic;
signal \c0.data_in_frame_9_7\ : std_logic;
signal \c0.n5_adj_4268\ : std_logic;
signal \c0.n4_adj_4267\ : std_logic;
signal \c0.n4_adj_4269\ : std_logic;
signal \c0.n22196\ : std_logic;
signal \c0.n4_adj_4269_cascade_\ : std_logic;
signal \c0.n68\ : std_logic;
signal \c0.n89_cascade_\ : std_logic;
signal \c0.n23_cascade_\ : std_logic;
signal \c0.n26\ : std_logic;
signal \c0.n13075_cascade_\ : std_logic;
signal \c0.n93_cascade_\ : std_logic;
signal data_in_frame_14_1 : std_logic;
signal \c0.n102\ : std_logic;
signal \c0.n147_cascade_\ : std_logic;
signal \c0.n134\ : std_logic;
signal \c0.n131\ : std_logic;
signal \c0.n31_adj_4284\ : std_logic;
signal \c0.n36_adj_4447\ : std_logic;
signal \c0.n41_adj_4452_cascade_\ : std_logic;
signal \c0.data_in_frame_11_7\ : std_logic;
signal \c0.n39_adj_4453\ : std_logic;
signal \c0.n40_adj_4451\ : std_logic;
signal \c0.n14016\ : std_logic;
signal \c0.n13223\ : std_logic;
signal \c0.n16_adj_4608\ : std_logic;
signal \c0.n21\ : std_logic;
signal \c0.n20\ : std_logic;
signal \c0.n13_adj_4610\ : std_logic;
signal \c0.data_in_frame_4_1\ : std_logic;
signal \c0.data_in_frame_10_4\ : std_logic;
signal \c0.n22455\ : std_logic;
signal \c0.data_in_frame_12_5\ : std_logic;
signal \c0.n42\ : std_logic;
signal \c0.n58\ : std_logic;
signal \c0.n127\ : std_logic;
signal \c0.n5_adj_4311\ : std_logic;
signal \c0.n5_adj_4311_cascade_\ : std_logic;
signal \c0.data_in_frame_10_3\ : std_logic;
signal \c0.n23677\ : std_logic;
signal data_in_frame_14_4 : std_logic;
signal \c0.data_in_frame_8_2\ : std_logic;
signal \c0.n120_cascade_\ : std_logic;
signal \c0.n142\ : std_logic;
signal \c0.n152_cascade_\ : std_logic;
signal \c0.n158\ : std_logic;
signal \c0.n22472\ : std_logic;
signal data_in_frame_14_3 : std_logic;
signal \c0.n30_adj_4571_cascade_\ : std_logic;
signal \c0.n33\ : std_logic;
signal \c0.n34_adj_4600_cascade_\ : std_logic;
signal \c0.n38_adj_4573\ : std_logic;
signal \c0.n24333_cascade_\ : std_logic;
signal \c0.n23661\ : std_logic;
signal \c0.data_in_frame_18_5\ : std_logic;
signal \c0.data_in_frame_16_3\ : std_logic;
signal \c0.n155\ : std_logic;
signal \c0.n160\ : std_logic;
signal \c0.n12989\ : std_logic;
signal \c0.n22104_cascade_\ : std_logic;
signal \c0.data_in_frame_19_4\ : std_logic;
signal \c0.n22347_cascade_\ : std_logic;
signal \c0.n24520\ : std_logic;
signal \c0.data_in_frame_20_5\ : std_logic;
signal \c0.n22_adj_4350\ : std_logic;
signal \c0.n22_adj_4350_cascade_\ : std_logic;
signal \c0.data_in_frame_20_6\ : std_logic;
signal \c0.data_in_frame_20_7\ : std_logic;
signal \c0.n21_adj_4225\ : std_logic;
signal \c0.n22227\ : std_logic;
signal \c0.n23863\ : std_logic;
signal \c0.n9_adj_4521\ : std_logic;
signal \c0.n20_adj_4596\ : std_logic;
signal \c0.n23733_cascade_\ : std_logic;
signal \c0.data_in_frame_26_0\ : std_logic;
signal \c0.data_in_frame_27_7\ : std_logic;
signal \c0.n20314_cascade_\ : std_logic;
signal \c0.n21325\ : std_logic;
signal \c0.n20314\ : std_logic;
signal \c0.n22_adj_4597\ : std_logic;
signal \c0.n12_adj_4671\ : std_logic;
signal \c0.data_in_frame_29_7\ : std_logic;
signal \c0.data_in_frame_27_5\ : std_logic;
signal \c0.data_in_frame_27_6\ : std_logic;
signal \c0.data_in_frame_25_5\ : std_logic;
signal \c0.n12_adj_4466\ : std_logic;
signal \c0.n11_adj_4474_cascade_\ : std_logic;
signal \c0.n21280\ : std_logic;
signal \c0.data_in_frame_29_2\ : std_logic;
signal \c0.n25446\ : std_logic;
signal \c0.data_in_frame_29_0\ : std_logic;
signal \c0.n10874\ : std_logic;
signal \c0.n43_adj_4463_cascade_\ : std_logic;
signal \c0.n21389\ : std_logic;
signal \c0.data_in_frame_25_0\ : std_logic;
signal \c0.n64_adj_4539\ : std_logic;
signal \c0.n10_adj_4544\ : std_logic;
signal \c0.n13911\ : std_logic;
signal \c0.n23921_cascade_\ : std_logic;
signal \c0.n21_adj_4547\ : std_logic;
signal \c0.n23975\ : std_logic;
signal \c0.n32_adj_4533\ : std_logic;
signal \c0.n74\ : std_logic;
signal \c0.n70_adj_4514\ : std_logic;
signal \c0.n71_cascade_\ : std_logic;
signal \c0.n17537\ : std_logic;
signal \c0.n81_cascade_\ : std_logic;
signal \c0.n82_adj_4517\ : std_logic;
signal \c0.n28_adj_4523\ : std_logic;
signal \c0.data_in_frame_27_3\ : std_logic;
signal \c0.data_in_frame_27_4\ : std_logic;
signal \c0.n23_adj_4532_cascade_\ : std_logic;
signal \c0.n31_adj_4542\ : std_logic;
signal \c0.n38_adj_4535_cascade_\ : std_logic;
signal \c0.n32_adj_4534\ : std_logic;
signal \c0.n8_adj_4677\ : std_logic;
signal \c0.data_in_frame_9_6\ : std_logic;
signal data_in_frame_5_3 : std_logic;
signal data_in_frame_5_2 : std_logic;
signal \c0.data_in_frame_7_6\ : std_logic;
signal data_in_frame_1_2 : std_logic;
signal \c0.n12_adj_4612\ : std_logic;
signal \c0.n15_adj_4444\ : std_logic;
signal \c0.n15_adj_4444_cascade_\ : std_logic;
signal \c0.n11_adj_4656\ : std_logic;
signal \c0.data_in_frame_3_2\ : std_logic;
signal data_in_frame_5_4 : std_logic;
signal \c0.n6_adj_4611\ : std_logic;
signal \c0.n6_adj_4611_cascade_\ : std_logic;
signal \c0.n91\ : std_logic;
signal \c0.n13453\ : std_logic;
signal \c0.n13_adj_4584\ : std_logic;
signal \c0.n102_adj_4445\ : std_logic;
signal \c0.n101\ : std_logic;
signal \c0.n103\ : std_logic;
signal \c0.n98\ : std_logic;
signal \c0.n97\ : std_logic;
signal \c0.n110_cascade_\ : std_logic;
signal \c0.n24465\ : std_logic;
signal \c0.data_out_frame_0__7__N_2579\ : std_logic;
signal \c0.n15_adj_4450\ : std_logic;
signal \c0.n87\ : std_logic;
signal \c0.n85\ : std_logic;
signal \c0.n88\ : std_logic;
signal \c0.n87_cascade_\ : std_logic;
signal \c0.n106\ : std_logic;
signal \c0.n22160\ : std_logic;
signal \c0.n7_adj_4304\ : std_logic;
signal \c0.n7_adj_4304_cascade_\ : std_logic;
signal data_in_frame_5_7 : std_logic;
signal data_in_frame_6_0 : std_logic;
signal \c0.n27_adj_4725\ : std_logic;
signal \c0.n17_adj_4224\ : std_logic;
signal \c0.n130\ : std_logic;
signal \c0.n14_adj_4707\ : std_logic;
signal \c0.n15_adj_4710\ : std_logic;
signal \c0.n22511\ : std_logic;
signal \c0.n22_adj_4259\ : std_logic;
signal data_in_frame_6_1 : std_logic;
signal \c0.n18_adj_4314_cascade_\ : std_logic;
signal \c0.data_in_frame_3_7\ : std_logic;
signal data_in_frame_1_6 : std_logic;
signal \c0.n38_adj_4448\ : std_logic;
signal \c0.n42_adj_4449\ : std_logic;
signal \c0.data_in_frame_3_3\ : std_logic;
signal \c0.n24_adj_4689\ : std_logic;
signal \c0.n13_adj_4281\ : std_logic;
signal \c0.n31\ : std_logic;
signal \c0.n31_cascade_\ : std_logic;
signal \c0.data_in_frame_10_0\ : std_logic;
signal \c0.n28\ : std_logic;
signal \c0.n24\ : std_logic;
signal \c0.n16\ : std_logic;
signal data_in_frame_14_2 : std_logic;
signal \c0.n8_adj_4673\ : std_logic;
signal data_in_frame_6_2 : std_logic;
signal \c0.data_in_frame_13_0\ : std_logic;
signal \c0.n22205_cascade_\ : std_logic;
signal \c0.n23491\ : std_logic;
signal \c0.n23598_cascade_\ : std_logic;
signal \c0.n23611\ : std_logic;
signal \c0.n9_adj_4208_cascade_\ : std_logic;
signal \c0.n22304\ : std_logic;
signal \c0.n13892_cascade_\ : std_logic;
signal \c0.data_in_frame_11_6\ : std_logic;
signal \c0.n13892\ : std_logic;
signal \c0.data_in_frame_17_2\ : std_logic;
signal \c0.n22_adj_4622\ : std_logic;
signal \c0.n22825_cascade_\ : std_logic;
signal data_in_frame_14_0 : std_logic;
signal \c0.n136\ : std_logic;
signal \c0.n22751_cascade_\ : std_logic;
signal \c0.n107\ : std_logic;
signal \c0.n149\ : std_logic;
signal \c0.n140\ : std_logic;
signal \c0.n22843\ : std_logic;
signal \c0.n22_adj_4245\ : std_logic;
signal \c0.n22514_cascade_\ : std_logic;
signal \c0.data_in_frame_16_1\ : std_logic;
signal \c0.n14_adj_4566\ : std_logic;
signal \c0.n14165_cascade_\ : std_logic;
signal \c0.data_in_frame_12_4\ : std_logic;
signal \c0.n4_adj_4658_cascade_\ : std_logic;
signal \c0.n24433\ : std_logic;
signal \c0.data_in_frame_16_6\ : std_logic;
signal \c0.n12_adj_4682_cascade_\ : std_logic;
signal \c0.n23390\ : std_logic;
signal \c0.n22249\ : std_logic;
signal \c0.n10_adj_4315\ : std_logic;
signal \c0.n24534\ : std_logic;
signal \c0.data_in_frame_17_3\ : std_logic;
signal \c0.n4_adj_4345\ : std_logic;
signal \c0.n24534_cascade_\ : std_logic;
signal \c0.n12_adj_4346\ : std_logic;
signal \c0.n13329\ : std_logic;
signal \c0.n4_adj_4621\ : std_logic;
signal \c0.n12_adj_4500\ : std_logic;
signal \c0.n9_adj_4208\ : std_logic;
signal \c0.n6_adj_4587_cascade_\ : std_logic;
signal \c0.n13461\ : std_logic;
signal \c0.n13756\ : std_logic;
signal \c0.n13461_cascade_\ : std_logic;
signal \c0.n6227_cascade_\ : std_logic;
signal \c0.n22173\ : std_logic;
signal \c0.n19_adj_4291\ : std_logic;
signal data_in_frame_14_6 : std_logic;
signal n22118 : std_logic;
signal \c0.data_in_frame_19_3\ : std_logic;
signal \c0.n14088\ : std_logic;
signal \c0.n23300\ : std_logic;
signal \c0.n6_adj_4577\ : std_logic;
signal \c0.n22662\ : std_logic;
signal \c0.n23300_cascade_\ : std_logic;
signal \c0.n21_adj_4594\ : std_logic;
signal \c0.n4_adj_4347\ : std_logic;
signal \c0.data_in_frame_23_4\ : std_logic;
signal \c0.n4_adj_4347_cascade_\ : std_logic;
signal \c0.data_in_frame_23_1\ : std_logic;
signal \c0.n30_adj_4357_cascade_\ : std_logic;
signal \c0.n14_adj_4356\ : std_logic;
signal \c0.n40_adj_4359\ : std_logic;
signal \c0.n42_adj_4358_cascade_\ : std_logic;
signal \c0.n41_adj_4360\ : std_logic;
signal \c0.n37_adj_4458\ : std_logic;
signal \c0.n34_adj_4361_cascade_\ : std_logic;
signal \c0.n14148\ : std_logic;
signal \c0.data_in_frame_20_4\ : std_logic;
signal \c0.n30_adj_4357\ : std_logic;
signal \c0.n22334\ : std_logic;
signal \c0.data_in_frame_25_6\ : std_logic;
signal \c0.data_in_frame_24_3\ : std_logic;
signal \c0.n24547\ : std_logic;
signal \c0.n21353\ : std_logic;
signal \c0.n66_cascade_\ : std_logic;
signal \c0.n75\ : std_logic;
signal \c0.n46_adj_4461\ : std_logic;
signal \c0.n10_adj_4513\ : std_logic;
signal \c0.n15_adj_4497\ : std_logic;
signal \c0.data_in_frame_25_4\ : std_logic;
signal \c0.n23_adj_4551\ : std_logic;
signal \c0.n26_adj_4548\ : std_logic;
signal \c0.n24_adj_4550_cascade_\ : std_logic;
signal \c0.n21010_cascade_\ : std_logic;
signal \c0.n53_adj_4538\ : std_logic;
signal \c0.n61_adj_4543\ : std_logic;
signal \c0.n42_adj_4540\ : std_logic;
signal \c0.n62_adj_4541\ : std_logic;
signal \c0.n13_adj_4492\ : std_logic;
signal \c0.n18_adj_4493\ : std_logic;
signal \c0.n22_adj_4498\ : std_logic;
signal \c0.n26_adj_4499_cascade_\ : std_logic;
signal \c0.n24441_cascade_\ : std_logic;
signal \c0.n30_adj_4545\ : std_logic;
signal \c0.n72\ : std_logic;
signal \c0.n24559\ : std_logic;
signal \c0.n42_adj_4510\ : std_logic;
signal \c0.n20_adj_4518\ : std_logic;
signal \c0.n24751\ : std_logic;
signal \c0.n14_adj_4676_cascade_\ : std_logic;
signal \c0.data_out_frame_0__7__N_2777\ : std_logic;
signal \c0.data_in_frame_0_6\ : std_logic;
signal \c0.n24016\ : std_logic;
signal \c0.n24749\ : std_logic;
signal data_in_frame_1_4 : std_logic;
signal data_in_frame_1_5 : std_logic;
signal \c0.n37_adj_4738\ : std_logic;
signal \c0.data_in_frame_0_5\ : std_logic;
signal \c0.data_in_frame_0_7\ : std_logic;
signal \c0.n22316\ : std_logic;
signal \c0.n23554\ : std_logic;
signal \c0.n34_cascade_\ : std_logic;
signal \c0.n23655\ : std_logic;
signal \c0.n53\ : std_logic;
signal \c0.n54_cascade_\ : std_logic;
signal \c0.n56\ : std_logic;
signal \c0.n13821\ : std_logic;
signal \c0.n48\ : std_logic;
signal \c0.n37_cascade_\ : std_logic;
signal \c0.n22647_cascade_\ : std_logic;
signal \c0.data_in_frame_2_6\ : std_logic;
signal \c0.n24747\ : std_logic;
signal \c0.n10_adj_4722\ : std_logic;
signal \c0.n14_adj_4616_cascade_\ : std_logic;
signal \c0.n23666\ : std_logic;
signal \c0.n37\ : std_logic;
signal \c0.n55\ : std_logic;
signal \c0.n18_adj_4314\ : std_logic;
signal \c0.n24_adj_4724\ : std_logic;
signal data_in_frame_1_0 : std_logic;
signal \c0.n5_adj_4711\ : std_logic;
signal \c0.n16_adj_4716\ : std_logic;
signal \c0.n28_adj_4718_cascade_\ : std_logic;
signal \c0.n24_adj_4717\ : std_logic;
signal \c0.n23_adj_4599\ : std_logic;
signal \c0.n4_adj_4446\ : std_logic;
signal \c0.n4_adj_4446_cascade_\ : std_logic;
signal \c0.n26_adj_4714\ : std_logic;
signal \c0.data_in_frame_4_0\ : std_logic;
signal \c0.data_in_frame_3_6\ : std_logic;
signal \c0.n23597\ : std_logic;
signal \c0.data_in_frame_2_0\ : std_logic;
signal \c0.n22230\ : std_logic;
signal \c0.data_in_frame_9_4\ : std_logic;
signal \c0.n150\ : std_logic;
signal \c0.n13651\ : std_logic;
signal \c0.n18_adj_4228\ : std_logic;
signal \c0.n27_cascade_\ : std_logic;
signal \c0.n19\ : std_logic;
signal \c0.n23528_cascade_\ : std_logic;
signal \c0.n34_adj_4278_cascade_\ : std_logic;
signal \c0.n36\ : std_logic;
signal \c0.n48_adj_4227\ : std_logic;
signal \c0.n30_adj_4705_cascade_\ : std_logic;
signal \c0.n23523_cascade_\ : std_logic;
signal \c0.n30\ : std_logic;
signal \c0.n13075\ : std_logic;
signal \c0.n7_adj_4634_cascade_\ : std_logic;
signal \c0.data_in_frame_10_5\ : std_logic;
signal \c0.n96_cascade_\ : std_logic;
signal \c0.data_in_frame_8_0\ : std_logic;
signal \c0.n104\ : std_logic;
signal \c0.n7_adj_4253\ : std_logic;
signal \c0.n5_adj_4252\ : std_logic;
signal \c0.n5_adj_4443\ : std_logic;
signal \c0.n13734_cascade_\ : std_logic;
signal \c0.n17734\ : std_logic;
signal \c0.n12973\ : std_logic;
signal \c0.n13128\ : std_logic;
signal \c0.n7_adj_4603\ : std_logic;
signal \c0.n22589\ : std_logic;
signal \c0.n13738_cascade_\ : std_logic;
signal \c0.data_in_frame_10_6\ : std_logic;
signal \c0.data_in_frame_10_7\ : std_logic;
signal \c0.n13734\ : std_logic;
signal \c0.n39_adj_4708_cascade_\ : std_logic;
signal \c0.n63\ : std_logic;
signal \c0.n64_cascade_\ : std_logic;
signal \c0.n13721\ : std_logic;
signal \c0.n55_adj_4709\ : std_logic;
signal \c0.n13186\ : std_logic;
signal \c0.n124\ : std_logic;
signal \c0.n10_adj_4247\ : std_logic;
signal \c0.n22547\ : std_logic;
signal \c0.n13998\ : std_logic;
signal \c0.n23156\ : std_logic;
signal \c0.n65\ : std_logic;
signal \c0.n60\ : std_logic;
signal \c0.n59_cascade_\ : std_logic;
signal \c0.n70\ : std_logic;
signal \c0.n24444_cascade_\ : std_logic;
signal \c0.n21282\ : std_logic;
signal \c0.data_in_frame_15_7\ : std_logic;
signal \c0.n22514\ : std_logic;
signal \c0.n23224_cascade_\ : std_logic;
signal \c0.n21409\ : std_logic;
signal \c0.data_in_frame_18_6\ : std_logic;
signal \c0.n22540\ : std_logic;
signal \c0.n24333\ : std_logic;
signal \c0.n22822\ : std_logic;
signal data_in_frame_14_7 : std_logic;
signal \c0.n12_adj_4246_cascade_\ : std_logic;
signal \c0.n23691_cascade_\ : std_logic;
signal \c0.n20543\ : std_logic;
signal \c0.data_in_frame_16_5\ : std_logic;
signal \c0.n10_adj_4602\ : std_logic;
signal \c0.n22644\ : std_logic;
signal \c0.data_in_frame_15_1\ : std_logic;
signal \c0.n14165\ : std_logic;
signal data_in_frame_14_5 : std_logic;
signal \c0.n24444\ : std_logic;
signal \c0.n7_adj_4581\ : std_logic;
signal \c0.FRAME_MATCHER_i_3\ : std_logic;
signal \c0.n3_adj_4430\ : std_logic;
signal \c0.n20467\ : std_logic;
signal \c0.n20467_cascade_\ : std_logic;
signal \c0.n6404\ : std_logic;
signal \c0.n17_adj_4354_cascade_\ : std_logic;
signal \c0.n10_adj_4630\ : std_logic;
signal \c0.n23523\ : std_logic;
signal \c0.n6_adj_4209\ : std_logic;
signal \c0.data_in_frame_13_7\ : std_logic;
signal \c0.data_in_frame_12_6\ : std_logic;
signal \c0.n22782\ : std_logic;
signal \c0.n12_adj_4246\ : std_logic;
signal \c0.n23453\ : std_logic;
signal \c0.data_in_frame_12_7\ : std_logic;
signal \c0.n25_adj_4579\ : std_logic;
signal \c0.n25_adj_4579_cascade_\ : std_logic;
signal \c0.n23433_cascade_\ : std_logic;
signal \c0.n18_adj_4580\ : std_logic;
signal \c0.n24_adj_4655\ : std_logic;
signal \c0.n41_adj_4592\ : std_logic;
signal \c0.n43_adj_4661\ : std_logic;
signal \c0.n44_adj_4588\ : std_logic;
signal \c0.n39_adj_4341\ : std_logic;
signal \c0.n22205\ : std_logic;
signal \c0.n50_adj_4340_cascade_\ : std_logic;
signal \c0.n5_adj_4486\ : std_logic;
signal \c0.n12559_cascade_\ : std_logic;
signal \c0.n22375\ : std_logic;
signal \c0.n24451\ : std_logic;
signal \c0.data_in_frame_19_1\ : std_logic;
signal \c0.n6215\ : std_logic;
signal \c0.data_in_frame_19_2\ : std_logic;
signal \c0.n21275\ : std_logic;
signal \c0.n21275_cascade_\ : std_logic;
signal \c0.n14_adj_4440\ : std_logic;
signal \c0.n63_adj_4516\ : std_logic;
signal \c0.n14189\ : std_logic;
signal \c0.n46\ : std_logic;
signal \c0.n46_cascade_\ : std_logic;
signal \c0.n34_adj_4361\ : std_logic;
signal \c0.n57_cascade_\ : std_logic;
signal \c0.n48_adj_4365\ : std_logic;
signal \c0.n21426_cascade_\ : std_logic;
signal \c0.n23032\ : std_logic;
signal \c0.n23032_cascade_\ : std_logic;
signal \c0.n25456\ : std_logic;
signal \c0.n23209_cascade_\ : std_logic;
signal \c0.n56_adj_4479\ : std_logic;
signal \c0.n21299\ : std_logic;
signal data_in_frame_22_6 : std_logic;
signal data_in_frame_22_0 : std_logic;
signal \c0.data_in_frame_23_7\ : std_logic;
signal \c0.n7_adj_4364_cascade_\ : std_logic;
signal \c0.n21426\ : std_logic;
signal \c0.n23031_cascade_\ : std_logic;
signal \c0.data_in_frame_25_7\ : std_logic;
signal \c0.data_in_frame_26_5\ : std_logic;
signal \c0.n24482\ : std_logic;
signal \c0.n23031\ : std_logic;
signal \c0.data_in_frame_28_2\ : std_logic;
signal \c0.n36_adj_4460_cascade_\ : std_logic;
signal \c0.n41_adj_4511\ : std_logic;
signal \c0.n6_adj_4459\ : std_logic;
signal \c0.n22426\ : std_logic;
signal \c0.data_in_frame_26_1\ : std_logic;
signal \c0.n22340\ : std_logic;
signal \c0.n5_adj_4472_cascade_\ : std_logic;
signal \c0.n21010\ : std_logic;
signal \c0.n24_adj_4496\ : std_logic;
signal \c0.data_in_frame_24_1\ : std_logic;
signal \c0.data_in_frame_27_1\ : std_logic;
signal \c0.n39_adj_4515\ : std_logic;
signal \c0.n10_adj_4675\ : std_logic;
signal \c0.data_in_frame_11_0\ : std_logic;
signal \c0.data_in_frame_4_6\ : std_logic;
signal \c0.n4_adj_4211\ : std_logic;
signal \c0.n22647\ : std_logic;
signal \c0.n13904_cascade_\ : std_logic;
signal \c0.n21_adj_4327\ : std_logic;
signal \c0.n19_adj_4324_cascade_\ : std_logic;
signal \c0.n22417\ : std_logic;
signal \c0.data_in_frame_7_5\ : std_logic;
signal \c0.n22417_cascade_\ : std_logic;
signal \c0.n4_adj_4333\ : std_logic;
signal \c0.n86\ : std_logic;
signal \c0.n13085\ : std_logic;
signal \c0.n7_adj_4282\ : std_logic;
signal \c0.n50\ : std_logic;
signal \n22121_cascade_\ : std_logic;
signal data_in_frame_6_6 : std_logic;
signal \c0.data_in_frame_2_2\ : std_logic;
signal data_in_frame_6_7 : std_logic;
signal \c0.data_in_frame_4_7\ : std_logic;
signal \c0.data_in_frame_2_7\ : std_logic;
signal \c0.n49\ : std_logic;
signal \c0.n23528\ : std_logic;
signal \c0.n7_adj_4229\ : std_logic;
signal \c0.data_out_frame_0__7__N_2743\ : std_logic;
signal \c0.n13523\ : std_logic;
signal \c0.n47\ : std_logic;
signal \c0.n10_adj_4664\ : std_logic;
signal \c0.data_in_frame_9_2\ : std_logic;
signal \c0.data_in_frame_7_0\ : std_logic;
signal \c0.n23406\ : std_logic;
signal data_in_frame_6_4 : std_logic;
signal \c0.n14_adj_4609_cascade_\ : std_logic;
signal \c0.n10_adj_4617\ : std_logic;
signal \c0.n17\ : std_logic;
signal \c0.n8_adj_4216\ : std_logic;
signal \c0.n12_cascade_\ : std_logic;
signal \c0.data_in_frame_4_2\ : std_logic;
signal \c0.data_in_frame_12_2\ : std_logic;
signal \c0.n13809\ : std_logic;
signal \c0.data_in_frame_11_5\ : std_logic;
signal \c0.n22751\ : std_logic;
signal \c0.n23_adj_4665\ : std_logic;
signal \c0.data_in_frame_15_2\ : std_logic;
signal \c0.data_in_frame_8_5\ : std_logic;
signal \c0.data_in_frame_11_1\ : std_logic;
signal \c0.n22176\ : std_logic;
signal \c0.n28_adj_4637_cascade_\ : std_logic;
signal \c0.n24_adj_4636\ : std_logic;
signal \c0.n7_adj_4634\ : std_logic;
signal \c0.n16_adj_4635\ : std_logic;
signal \c0.data_in_frame_4_5\ : std_logic;
signal \c0.n23283\ : std_logic;
signal \c0.data_in_frame_8_7\ : std_logic;
signal \c0.n20_adj_4260\ : std_logic;
signal \c0.n22803\ : std_logic;
signal \c0.n4_adj_4261\ : std_logic;
signal \c0.n31_adj_4743\ : std_logic;
signal \c0.n5813\ : std_logic;
signal \c0.n22602\ : std_logic;
signal \c0.n11\ : std_logic;
signal \c0.n17_adj_4219\ : std_logic;
signal \c0.n16_adj_4218_cascade_\ : std_logic;
signal \c0.n13767_cascade_\ : std_logic;
signal \c0.n5965\ : std_logic;
signal \c0.n6_adj_4454\ : std_logic;
signal \c0.data_in_frame_15_3\ : std_logic;
signal \c0.n12_adj_4455\ : std_logic;
signal \c0.n22463\ : std_logic;
signal \c0.n24540\ : std_logic;
signal \c0.n23507\ : std_logic;
signal data_in_frame_21_0 : std_logic;
signal \c0.data_in_frame_17_0\ : std_logic;
signal \c0.n23313\ : std_logic;
signal \c0.n26_adj_4578\ : std_logic;
signal \c0.data_in_frame_13_5\ : std_logic;
signal \c0.data_in_frame_17_7\ : std_logic;
signal \c0.data_in_frame_16_2\ : std_logic;
signal \c0.n24527\ : std_logic;
signal data_in_frame_21_3 : std_logic;
signal \c0.n21344\ : std_logic;
signal \c0.n42_adj_4589\ : std_logic;
signal \c0.n22_adj_4243\ : std_logic;
signal \c0.n13738\ : std_logic;
signal \c0.n10_adj_4230\ : std_logic;
signal \c0.n5_adj_4310\ : std_logic;
signal \c0.n13604\ : std_logic;
signal \c0.n7_adj_4251_cascade_\ : std_logic;
signal \c0.n23224\ : std_logic;
signal \c0.n7_adj_4251\ : std_logic;
signal data_in_frame_22_7 : std_logic;
signal \c0.n22825\ : std_logic;
signal \c0.data_in_frame_15_4\ : std_logic;
signal \c0.data_in_frame_18_2\ : std_logic;
signal \c0.data_in_frame_18_4\ : std_logic;
signal \c0.data_in_frame_18_3\ : std_logic;
signal \c0.n5_adj_4335\ : std_logic;
signal \c0.n4_adj_4568\ : std_logic;
signal \c0.n15_adj_4569\ : std_logic;
signal \c0.data_in_frame_18_7\ : std_logic;
signal data_in_frame_22_5 : std_logic;
signal \c0.data_in_frame_17_5\ : std_logic;
signal \c0.n22748\ : std_logic;
signal \c0.n14_adj_4623_cascade_\ : std_logic;
signal \c0.n15_adj_4624\ : std_logic;
signal data_in_frame_21_1 : std_logic;
signal \c0.n13963_cascade_\ : std_logic;
signal \c0.n22508\ : std_logic;
signal \c0.n40_adj_4342\ : std_logic;
signal \c0.data_in_frame_24_6\ : std_logic;
signal \c0.n22495\ : std_logic;
signal \c0.data_in_frame_20_1\ : std_logic;
signal \c0.n58_adj_4355\ : std_logic;
signal \c0.n59_adj_4351\ : std_logic;
signal \c0.n28_adj_4363\ : std_logic;
signal \c0.n23691\ : std_logic;
signal \c0.n22577\ : std_logic;
signal \c0.n21414\ : std_logic;
signal \c0.n10_adj_4524_cascade_\ : std_logic;
signal \c0.n13797\ : std_logic;
signal \c0.n24576\ : std_logic;
signal \c0.data_in_frame_26_2\ : std_logic;
signal \c0.n24576_cascade_\ : std_logic;
signal \c0.n14_adj_4519\ : std_logic;
signal data_in_frame_21_4 : std_logic;
signal \c0.n23733\ : std_logic;
signal \c0.n22686\ : std_logic;
signal \c0.n5_adj_4472\ : std_logic;
signal \c0.n22686_cascade_\ : std_logic;
signal \c0.n21316\ : std_logic;
signal \c0.n39_adj_4487\ : std_logic;
signal \c0.n30_adj_4489_cascade_\ : std_logic;
signal \c0.n23209\ : std_logic;
signal \c0.n45_adj_4490_cascade_\ : std_logic;
signal \c0.n44_adj_4501\ : std_logic;
signal \c0.n11_adj_4505\ : std_logic;
signal \c0.n48_adj_4503_cascade_\ : std_logic;
signal \c0.n28_adj_4504\ : std_logic;
signal \c0.n24573\ : std_logic;
signal \c0.n41_adj_4488\ : std_logic;
signal \c0.n17_adj_4354\ : std_logic;
signal \c0.n28_adj_4343\ : std_logic;
signal \c0.n27_adj_4502\ : std_logic;
signal \c0.data_in_frame_26_7\ : std_logic;
signal \c0.data_in_frame_24_4\ : std_logic;
signal data_in_frame_21_6 : std_logic;
signal \c0.n21301\ : std_logic;
signal \c0.n23_adj_4582\ : std_logic;
signal \c0.data_in_frame_27_2\ : std_logic;
signal \c0.n25_adj_4469\ : std_logic;
signal \c0.n26_adj_4470\ : std_logic;
signal \c0.n39_adj_4467\ : std_logic;
signal \c0.n38_adj_4468\ : std_logic;
signal \c0.n37_adj_4473\ : std_logic;
signal \c0.n44_adj_4471_cascade_\ : std_logic;
signal \c0.n45_adj_4476\ : std_logic;
signal \c0.n14_adj_4529\ : std_logic;
signal \c0.n15_adj_4508\ : std_logic;
signal \c0.n24362_cascade_\ : std_logic;
signal \c0.n18_adj_4475\ : std_logic;
signal \c0.n26_adj_4530\ : std_logic;
signal n22103 : std_logic;
signal \c0.n22632\ : std_logic;
signal \c0.n22632_cascade_\ : std_logic;
signal \c0.data_in_frame_24_2\ : std_logic;
signal \c0.data_in_frame_26_3\ : std_logic;
signal \c0.n22362_cascade_\ : std_logic;
signal \c0.n12559\ : std_logic;
signal \c0.n13_adj_4527\ : std_logic;
signal \c0.n20802\ : std_logic;
signal \c0.n20358\ : std_logic;
signal \c0.n12_adj_4491\ : std_logic;
signal \c0.data_in_frame_28_6\ : std_logic;
signal \c0.data_in_frame_28_4\ : std_logic;
signal \c0.n13904\ : std_logic;
signal \c0.n28_adj_4286\ : std_logic;
signal data_in_frame_5_0 : std_logic;
signal \c0.n23302\ : std_logic;
signal \c0.data_in_frame_0_3\ : std_logic;
signal \c0.data_in_frame_2_4\ : std_logic;
signal \c0.n42_adj_4746\ : std_logic;
signal \c0.data_in_frame_7_1\ : std_logic;
signal \c0.data_in_frame_2_5\ : std_logic;
signal \c0.data_in_frame_4_3\ : std_logic;
signal \c0.n6_adj_4687_cascade_\ : std_logic;
signal \c0.n23274\ : std_logic;
signal \c0.n23282\ : std_logic;
signal \c0.n23274_cascade_\ : std_logic;
signal \c0.n20_adj_4316\ : std_logic;
signal \c0.n29_adj_4287\ : std_logic;
signal \c0.data_in_frame_0_2\ : std_logic;
signal \c0.data_in_frame_2_3\ : std_logic;
signal \c0.data_in_frame_0_1\ : std_logic;
signal \c0.data_in_frame_4_4\ : std_logic;
signal \c0.n23276\ : std_logic;
signal \c0.n22322\ : std_logic;
signal \c0.n23276_cascade_\ : std_logic;
signal \c0.n25\ : std_logic;
signal \c0.n24_adj_4213\ : std_logic;
signal \c0.n8_cascade_\ : std_logic;
signal \c0.data_in_frame_0_4\ : std_logic;
signal n22121 : std_logic;
signal \c0.data_in_frame_0_0\ : std_logic;
signal \c0.n22701\ : std_logic;
signal \c0.n5_adj_4323\ : std_logic;
signal n22101 : std_logic;
signal \c0.n9_cascade_\ : std_logic;
signal \c0.data_in_frame_9_1\ : std_logic;
signal \c0.data_in_frame_8_6\ : std_logic;
signal \c0.data_in_frame_18_0\ : std_logic;
signal data_in_frame_6_5 : std_logic;
signal \c0.n19_adj_4620\ : std_logic;
signal \c0.n9\ : std_logic;
signal \c0.n22392\ : std_logic;
signal \c0.data_in_frame_9_5\ : std_logic;
signal \c0.FRAME_MATCHER_i_13\ : std_logic;
signal \c0.n3_adj_4410\ : std_logic;
signal \c0.data_in_frame_7_4\ : std_logic;
signal data_in_frame_5_1 : std_logic;
signal \c0.n40_adj_4288\ : std_logic;
signal \c0.n22120\ : std_logic;
signal \c0.data_in_frame_7_3\ : std_logic;
signal \c0.data_in_frame_12_0\ : std_logic;
signal \c0.data_in_frame_12_1\ : std_logic;
signal \c0.n39\ : std_logic;
signal \c0.n61\ : std_logic;
signal \c0.n13253\ : std_logic;
signal \c0.n13253_cascade_\ : std_logic;
signal \c0.n22518\ : std_logic;
signal \c0.n22828\ : std_logic;
signal \c0.data_in_frame_11_4\ : std_logic;
signal \c0.data_in_frame_7_2\ : std_logic;
signal \c0.n9_adj_4220\ : std_logic;
signal \c0.n7_adj_4226\ : std_logic;
signal \c0.n27_adj_4748\ : std_logic;
signal \c0.data_in_frame_11_3\ : std_logic;
signal \c0.data_in_frame_9_0\ : std_logic;
signal \c0.n4\ : std_logic;
signal \c0.data_in_frame_28_3\ : std_logic;
signal \c0.data_in_frame_12_3\ : std_logic;
signal \c0.data_in_frame_15_6\ : std_logic;
signal \c0.n22379\ : std_logic;
signal \c0.n6_adj_4559\ : std_logic;
signal \c0.data_in_frame_17_6\ : std_logic;
signal \c0.data_in_frame_15_5\ : std_logic;
signal \c0.n31_adj_4701\ : std_logic;
signal \c0.n13474\ : std_logic;
signal \c0.n22650\ : std_logic;
signal data_in_frame_1_7 : std_logic;
signal \c0.n30_adj_4747\ : std_logic;
signal \c0.n6_adj_4632\ : std_logic;
signal \c0.n5_adj_4631\ : std_logic;
signal \c0.n23343\ : std_logic;
signal \c0.n25_adj_4633\ : std_logic;
signal \c0.data_in_frame_9_3\ : std_logic;
signal \c0.data_in_frame_11_2\ : std_logic;
signal \c0.data_in_frame_28_1\ : std_logic;
signal \c0.data_in_frame_8_3\ : std_logic;
signal \c0.data_in_frame_17_4\ : std_logic;
signal \c0.data_in_frame_13_3\ : std_logic;
signal \c0.n22319\ : std_logic;
signal \c0.n4_adj_4586\ : std_logic;
signal \c0.data_in_frame_16_0\ : std_logic;
signal \c0.data_in_frame_13_6\ : std_logic;
signal \c0.data_in_frame_18_1\ : std_logic;
signal \c0.n14081\ : std_logic;
signal \c0.n10_adj_4250\ : std_logic;
signal \c0.data_in_frame_16_4\ : std_logic;
signal rx_data_4 : std_logic;
signal \c0.data_in_frame_13_4\ : std_logic;
signal \c0.data_in_frame_19_5\ : std_logic;
signal \c0.FRAME_MATCHER_i_18\ : std_logic;
signal \c0.n2119\ : std_logic;
signal \c0.n3_adj_4400\ : std_logic;
signal \c0.n22112\ : std_logic;
signal \c0.data_in_frame_15_0\ : std_logic;
signal rx_data_6 : std_logic;
signal data_in_frame_22_1 : std_logic;
signal \c0.data_in_frame_20_2\ : std_logic;
signal \c0.data_in_frame_23_5\ : std_logic;
signal \c0.n9_adj_4563\ : std_logic;
signal \c0.data_in_frame_16_7\ : std_logic;
signal \c0.n22_adj_4244\ : std_logic;
signal \c0.n24_adj_4618\ : std_logic;
signal \c0.n14_adj_4619\ : std_logic;
signal \c0.data_in_frame_2_1\ : std_logic;
signal \c0.n22288\ : std_logic;
signal \c0.data_in_frame_13_2\ : std_logic;
signal \c0.n22288_cascade_\ : std_logic;
signal \c0.n5807\ : std_logic;
signal \c0.n14160\ : std_logic;
signal \c0.data_in_frame_17_1\ : std_logic;
signal \c0.FRAME_MATCHER_i_2\ : std_logic;
signal \c0.FRAME_MATCHER_i_1\ : std_logic;
signal \c0.FRAME_MATCHER_i_0\ : std_logic;
signal \c0.n9_adj_4601\ : std_logic;
signal \c0.data_in_frame_25_1\ : std_logic;
signal \c0.data_in_frame_20_0\ : std_logic;
signal \c0.data_in_frame_19_0\ : std_logic;
signal \c0.n12_adj_4564\ : std_logic;
signal \c0.n21404\ : std_logic;
signal \c0.n6_adj_4462_cascade_\ : std_logic;
signal \c0.n22562\ : std_logic;
signal data_in_frame_22_3 : std_logic;
signal \c0.data_in_frame_26_6\ : std_logic;
signal \c0.n22769\ : std_logic;
signal data_in_frame_21_5 : std_logic;
signal \c0.n22698\ : std_logic;
signal \c0.data_in_frame_23_6\ : std_logic;
signal \c0.n4_adj_4464\ : std_logic;
signal \c0.n14_adj_4465\ : std_logic;
signal \c0.data_in_frame_20_3\ : std_logic;
signal \c0.n21412\ : std_logic;
signal \c0.n4_adj_4369\ : std_logic;
signal \c0.data_in_frame_27_0\ : std_logic;
signal \c0.n73\ : std_logic;
signal \c0.n20409\ : std_logic;
signal data_in_frame_22_4 : std_logic;
signal \c0.n12_adj_4672\ : std_logic;
signal \c0.n22099\ : std_logic;
signal rx_data_1 : std_logic;
signal \c0.data_in_frame_13_1\ : std_logic;
signal \c0.n13490\ : std_logic;
signal \c0.data_in_frame_24_5\ : std_logic;
signal \c0.n22505\ : std_logic;
signal \c0.n6718\ : std_logic;
signal \c0.n13963\ : std_logic;
signal \c0.n21295\ : std_logic;
signal \c0.n20239\ : std_logic;
signal \c0.n13468\ : std_logic;
signal \c0.n20239_cascade_\ : std_logic;
signal \c0.data_in_frame_26_4\ : std_logic;
signal \c0.n10_adj_4457\ : std_logic;
signal \c0.n6_adj_4668\ : std_logic;
signal \c0.data_in_frame_23_2\ : std_logic;
signal \c0.n13314\ : std_logic;
signal \c0.n6227\ : std_logic;
signal data_in_frame_21_7 : std_logic;
signal \c0.n20350\ : std_logic;
signal rx_data_3 : std_logic;
signal \c0.data_in_frame_23_3\ : std_logic;
signal \c0.n25484\ : std_logic;
signal \c0.n62\ : std_logic;
signal \c0.n21_adj_4481\ : std_logic;
signal \c0.n6_adj_4462\ : std_logic;
signal \c0.n30_adj_4482\ : std_logic;
signal \c0.n9_adj_4273\ : std_logic;
signal rx_data_7 : std_logic;
signal \c0.n23598\ : std_logic;
signal \c0.data_in_frame_8_4\ : std_logic;
signal data_in_frame_6_3 : std_logic;
signal \c0.n23267\ : std_logic;
signal \c0.n18_cascade_\ : std_logic;
signal \c0.n16_adj_4666\ : std_logic;
signal \c0.n28_adj_4667\ : std_logic;
signal \c0.n24_adj_4653_cascade_\ : std_logic;
signal \c0.n22369\ : std_logic;
signal \c0.n6_adj_4587\ : std_logic;
signal \c0.n22586\ : std_logic;
signal \c0.data_in_frame_19_6\ : std_logic;
signal \c0.data_in_frame_19_7\ : std_logic;
signal \c0.n23433\ : std_logic;
signal \c0.n15_adj_4625\ : std_logic;
signal \c0.n17_adj_4626\ : std_logic;
signal \c0.n16_adj_4627\ : std_logic;
signal \c0.n15_adj_4625_cascade_\ : std_logic;
signal \c0.n18\ : std_logic;
signal \c0.n22605\ : std_logic;
signal \c0.n13767\ : std_logic;
signal \c0.n19_adj_4595\ : std_logic;
signal \c0.n24_adj_4628\ : std_logic;
signal \c0.n14_adj_4629_cascade_\ : std_logic;
signal \c0.n23178\ : std_logic;
signal \c0.n22234\ : std_logic;
signal \c0.n17830\ : std_logic;
signal rx_data_0 : std_logic;
signal \c0.n22104\ : std_logic;
signal \c0.data_in_frame_23_0\ : std_logic;
signal \c0.n9_adj_4552\ : std_logic;
signal rx_data_5 : std_logic;
signal \c0.n22134\ : std_logic;
signal \c0.data_in_frame_28_5\ : std_logic;
signal rx_data_2 : std_logic;
signal n22110 : std_logic;
signal data_in_frame_22_2 : std_logic;
signal \CLK_c\ : std_logic;
signal \c0.data_in_frame_24_0\ : std_logic;
signal \c0.n29_adj_4362\ : std_logic;
signal \c0.n24_adj_4531\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \PIN_12_wire\ : std_logic;
signal \PIN_13_wire\ : std_logic;
signal \PIN_1_wire\ : std_logic;
signal \PIN_22_wire\ : std_logic;
signal \PIN_23_wire\ : std_logic;
signal \PIN_24_wire\ : std_logic;
signal \PIN_2_wire\ : std_logic;
signal \PIN_3_wire\ : std_logic;
signal \PIN_7_wire\ : std_logic;
signal \PIN_8_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    \PIN_12_wire\ <= PIN_12;
    \PIN_13_wire\ <= PIN_13;
    PIN_1 <= \PIN_1_wire\;
    PIN_22 <= \PIN_22_wire\;
    PIN_23 <= \PIN_23_wire\;
    PIN_24 <= \PIN_24_wire\;
    PIN_2 <= \PIN_2_wire\;
    PIN_3 <= \PIN_3_wire\;
    \PIN_7_wire\ <= PIN_7;
    \PIN_8_wire\ <= PIN_8;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81286\,
            DIN => \N__81285\,
            DOUT => \N__81284\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81286\,
            PADOUT => \N__81285\,
            PADIN => \N__81284\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__26751\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81277\,
            DIN => \N__81276\,
            DOUT => \N__81275\,
            PACKAGEPIN => \PIN_12_wire\
        );

    \PIN_12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81277\,
            PADOUT => \N__81276\,
            PADIN => \N__81275\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_12_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81268\,
            DIN => \N__81267\,
            DOUT => \N__81266\,
            PACKAGEPIN => \PIN_13_wire\
        );

    \PIN_13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81268\,
            PADOUT => \N__81267\,
            PADIN => \N__81266\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_13_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81259\,
            DIN => \N__81258\,
            DOUT => \N__81257\,
            PACKAGEPIN => \PIN_1_wire\
        );

    \PIN_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81259\,
            PADOUT => \N__81258\,
            PADIN => \N__81257\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81250\,
            DIN => \N__81249\,
            DOUT => \N__81248\,
            PACKAGEPIN => \PIN_22_wire\
        );

    \PIN_22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81250\,
            PADOUT => \N__81249\,
            PADIN => \N__81248\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81241\,
            DIN => \N__81240\,
            DOUT => \N__81239\,
            PACKAGEPIN => \PIN_23_wire\
        );

    \PIN_23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81241\,
            PADOUT => \N__81240\,
            PADIN => \N__81239\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81232\,
            DIN => \N__81231\,
            DOUT => \N__81230\,
            PACKAGEPIN => \PIN_24_wire\
        );

    \PIN_24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81232\,
            PADOUT => \N__81231\,
            PADIN => \N__81230\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81223\,
            DIN => \N__81222\,
            DOUT => \N__81221\,
            PACKAGEPIN => \PIN_2_wire\
        );

    \PIN_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81223\,
            PADOUT => \N__81222\,
            PADIN => \N__81221\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81214\,
            DIN => \N__81213\,
            DOUT => \N__81212\,
            PACKAGEPIN => \PIN_3_wire\
        );

    \PIN_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81214\,
            PADOUT => \N__81213\,
            PADIN => \N__81212\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81205\,
            DIN => \N__81204\,
            DOUT => \N__81203\,
            PACKAGEPIN => \PIN_7_wire\
        );

    \PIN_7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81205\,
            PADOUT => \N__81204\,
            PADIN => \N__81203\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_7_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81196\,
            DIN => \N__81195\,
            DOUT => \N__81194\,
            PACKAGEPIN => \PIN_8_wire\
        );

    \PIN_8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81196\,
            PADOUT => \N__81195\,
            PADIN => \N__81194\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_8_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81187\,
            DIN => \N__81186\,
            DOUT => \N__81185\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81187\,
            PADOUT => \N__81186\,
            PADIN => \N__81185\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall1_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__81178\,
            DIN => \N__81177\,
            DOUT => \N__81176\,
            PACKAGEPIN => PIN_4
        );

    \hall1_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81178\,
            PADOUT => \N__81177\,
            PADIN => \N__81176\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall2_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__81169\,
            DIN => \N__81168\,
            DOUT => \N__81167\,
            PACKAGEPIN => PIN_5
        );

    \hall2_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81169\,
            PADOUT => \N__81168\,
            PADIN => \N__81167\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall3_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__81160\,
            DIN => \N__81159\,
            DOUT => \N__81158\,
            PACKAGEPIN => PIN_6
        );

    \hall3_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81160\,
            PADOUT => \N__81159\,
            PADIN => \N__81158\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__81151\,
            DIN => \N__81150\,
            DOUT => \N__81149\,
            PACKAGEPIN => PIN_11
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81151\,
            PADOUT => \N__81150\,
            PADIN => \N__81149\,
            CLOCKENABLE => 'H',
            DIN0 => \LED_c\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__81142\,
            DIN => \N__81141\,
            DOUT => \N__81140\,
            PACKAGEPIN => PIN_10
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81142\,
            PADOUT => \N__81141\,
            PADIN => \N__81140\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__28599\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__26757\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__81133\,
            DIN => \N__81132\,
            DOUT => \N__81131\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__81133\,
            PADOUT => \N__81132\,
            PADIN => \N__81131\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__20379\ : CascadeMux
    port map (
            O => \N__81114\,
            I => \N__81111\
        );

    \I__20378\ : InMux
    port map (
            O => \N__81111\,
            I => \N__81108\
        );

    \I__20377\ : LocalMux
    port map (
            O => \N__81108\,
            I => \N__81105\
        );

    \I__20376\ : Span4Mux_h
    port map (
            O => \N__81105\,
            I => \N__81100\
        );

    \I__20375\ : InMux
    port map (
            O => \N__81104\,
            I => \N__81097\
        );

    \I__20374\ : InMux
    port map (
            O => \N__81103\,
            I => \N__81094\
        );

    \I__20373\ : Span4Mux_v
    port map (
            O => \N__81100\,
            I => \N__81091\
        );

    \I__20372\ : LocalMux
    port map (
            O => \N__81097\,
            I => \N__81086\
        );

    \I__20371\ : LocalMux
    port map (
            O => \N__81094\,
            I => \N__81086\
        );

    \I__20370\ : Odrv4
    port map (
            O => \N__81091\,
            I => \c0.n19_adj_4595\
        );

    \I__20369\ : Odrv12
    port map (
            O => \N__81086\,
            I => \c0.n19_adj_4595\
        );

    \I__20368\ : InMux
    port map (
            O => \N__81081\,
            I => \N__81078\
        );

    \I__20367\ : LocalMux
    port map (
            O => \N__81078\,
            I => \c0.n24_adj_4628\
        );

    \I__20366\ : CascadeMux
    port map (
            O => \N__81075\,
            I => \c0.n14_adj_4629_cascade_\
        );

    \I__20365\ : InMux
    port map (
            O => \N__81072\,
            I => \N__81068\
        );

    \I__20364\ : InMux
    port map (
            O => \N__81071\,
            I => \N__81065\
        );

    \I__20363\ : LocalMux
    port map (
            O => \N__81068\,
            I => \N__81062\
        );

    \I__20362\ : LocalMux
    port map (
            O => \N__81065\,
            I => \N__81059\
        );

    \I__20361\ : Span4Mux_v
    port map (
            O => \N__81062\,
            I => \N__81054\
        );

    \I__20360\ : Span4Mux_h
    port map (
            O => \N__81059\,
            I => \N__81051\
        );

    \I__20359\ : InMux
    port map (
            O => \N__81058\,
            I => \N__81048\
        );

    \I__20358\ : InMux
    port map (
            O => \N__81057\,
            I => \N__81045\
        );

    \I__20357\ : Span4Mux_h
    port map (
            O => \N__81054\,
            I => \N__81042\
        );

    \I__20356\ : Span4Mux_h
    port map (
            O => \N__81051\,
            I => \N__81039\
        );

    \I__20355\ : LocalMux
    port map (
            O => \N__81048\,
            I => \N__81036\
        );

    \I__20354\ : LocalMux
    port map (
            O => \N__81045\,
            I => \N__81033\
        );

    \I__20353\ : Span4Mux_v
    port map (
            O => \N__81042\,
            I => \N__81028\
        );

    \I__20352\ : Span4Mux_v
    port map (
            O => \N__81039\,
            I => \N__81025\
        );

    \I__20351\ : Span4Mux_v
    port map (
            O => \N__81036\,
            I => \N__81020\
        );

    \I__20350\ : Span4Mux_h
    port map (
            O => \N__81033\,
            I => \N__81020\
        );

    \I__20349\ : InMux
    port map (
            O => \N__81032\,
            I => \N__81015\
        );

    \I__20348\ : InMux
    port map (
            O => \N__81031\,
            I => \N__81015\
        );

    \I__20347\ : Odrv4
    port map (
            O => \N__81028\,
            I => \c0.n23178\
        );

    \I__20346\ : Odrv4
    port map (
            O => \N__81025\,
            I => \c0.n23178\
        );

    \I__20345\ : Odrv4
    port map (
            O => \N__81020\,
            I => \c0.n23178\
        );

    \I__20344\ : LocalMux
    port map (
            O => \N__81015\,
            I => \c0.n23178\
        );

    \I__20343\ : InMux
    port map (
            O => \N__81006\,
            I => \N__81003\
        );

    \I__20342\ : LocalMux
    port map (
            O => \N__81003\,
            I => \N__80999\
        );

    \I__20341\ : InMux
    port map (
            O => \N__81002\,
            I => \N__80996\
        );

    \I__20340\ : Span4Mux_v
    port map (
            O => \N__80999\,
            I => \N__80991\
        );

    \I__20339\ : LocalMux
    port map (
            O => \N__80996\,
            I => \N__80991\
        );

    \I__20338\ : Odrv4
    port map (
            O => \N__80991\,
            I => \c0.n22234\
        );

    \I__20337\ : InMux
    port map (
            O => \N__80988\,
            I => \N__80983\
        );

    \I__20336\ : InMux
    port map (
            O => \N__80987\,
            I => \N__80979\
        );

    \I__20335\ : CascadeMux
    port map (
            O => \N__80986\,
            I => \N__80976\
        );

    \I__20334\ : LocalMux
    port map (
            O => \N__80983\,
            I => \N__80970\
        );

    \I__20333\ : CascadeMux
    port map (
            O => \N__80982\,
            I => \N__80967\
        );

    \I__20332\ : LocalMux
    port map (
            O => \N__80979\,
            I => \N__80963\
        );

    \I__20331\ : InMux
    port map (
            O => \N__80976\,
            I => \N__80960\
        );

    \I__20330\ : InMux
    port map (
            O => \N__80975\,
            I => \N__80957\
        );

    \I__20329\ : InMux
    port map (
            O => \N__80974\,
            I => \N__80952\
        );

    \I__20328\ : InMux
    port map (
            O => \N__80973\,
            I => \N__80952\
        );

    \I__20327\ : Span4Mux_v
    port map (
            O => \N__80970\,
            I => \N__80948\
        );

    \I__20326\ : InMux
    port map (
            O => \N__80967\,
            I => \N__80945\
        );

    \I__20325\ : InMux
    port map (
            O => \N__80966\,
            I => \N__80937\
        );

    \I__20324\ : Span4Mux_v
    port map (
            O => \N__80963\,
            I => \N__80928\
        );

    \I__20323\ : LocalMux
    port map (
            O => \N__80960\,
            I => \N__80928\
        );

    \I__20322\ : LocalMux
    port map (
            O => \N__80957\,
            I => \N__80928\
        );

    \I__20321\ : LocalMux
    port map (
            O => \N__80952\,
            I => \N__80928\
        );

    \I__20320\ : CascadeMux
    port map (
            O => \N__80951\,
            I => \N__80925\
        );

    \I__20319\ : Span4Mux_h
    port map (
            O => \N__80948\,
            I => \N__80913\
        );

    \I__20318\ : LocalMux
    port map (
            O => \N__80945\,
            I => \N__80913\
        );

    \I__20317\ : InMux
    port map (
            O => \N__80944\,
            I => \N__80908\
        );

    \I__20316\ : InMux
    port map (
            O => \N__80943\,
            I => \N__80908\
        );

    \I__20315\ : InMux
    port map (
            O => \N__80942\,
            I => \N__80905\
        );

    \I__20314\ : InMux
    port map (
            O => \N__80941\,
            I => \N__80900\
        );

    \I__20313\ : InMux
    port map (
            O => \N__80940\,
            I => \N__80900\
        );

    \I__20312\ : LocalMux
    port map (
            O => \N__80937\,
            I => \N__80894\
        );

    \I__20311\ : Span4Mux_v
    port map (
            O => \N__80928\,
            I => \N__80894\
        );

    \I__20310\ : InMux
    port map (
            O => \N__80925\,
            I => \N__80889\
        );

    \I__20309\ : InMux
    port map (
            O => \N__80924\,
            I => \N__80889\
        );

    \I__20308\ : InMux
    port map (
            O => \N__80923\,
            I => \N__80885\
        );

    \I__20307\ : InMux
    port map (
            O => \N__80922\,
            I => \N__80882\
        );

    \I__20306\ : InMux
    port map (
            O => \N__80921\,
            I => \N__80875\
        );

    \I__20305\ : InMux
    port map (
            O => \N__80920\,
            I => \N__80875\
        );

    \I__20304\ : InMux
    port map (
            O => \N__80919\,
            I => \N__80875\
        );

    \I__20303\ : InMux
    port map (
            O => \N__80918\,
            I => \N__80872\
        );

    \I__20302\ : Span4Mux_v
    port map (
            O => \N__80913\,
            I => \N__80868\
        );

    \I__20301\ : LocalMux
    port map (
            O => \N__80908\,
            I => \N__80864\
        );

    \I__20300\ : LocalMux
    port map (
            O => \N__80905\,
            I => \N__80859\
        );

    \I__20299\ : LocalMux
    port map (
            O => \N__80900\,
            I => \N__80859\
        );

    \I__20298\ : InMux
    port map (
            O => \N__80899\,
            I => \N__80856\
        );

    \I__20297\ : Span4Mux_h
    port map (
            O => \N__80894\,
            I => \N__80853\
        );

    \I__20296\ : LocalMux
    port map (
            O => \N__80889\,
            I => \N__80850\
        );

    \I__20295\ : InMux
    port map (
            O => \N__80888\,
            I => \N__80847\
        );

    \I__20294\ : LocalMux
    port map (
            O => \N__80885\,
            I => \N__80844\
        );

    \I__20293\ : LocalMux
    port map (
            O => \N__80882\,
            I => \N__80840\
        );

    \I__20292\ : LocalMux
    port map (
            O => \N__80875\,
            I => \N__80837\
        );

    \I__20291\ : LocalMux
    port map (
            O => \N__80872\,
            I => \N__80834\
        );

    \I__20290\ : InMux
    port map (
            O => \N__80871\,
            I => \N__80831\
        );

    \I__20289\ : Span4Mux_v
    port map (
            O => \N__80868\,
            I => \N__80828\
        );

    \I__20288\ : InMux
    port map (
            O => \N__80867\,
            I => \N__80825\
        );

    \I__20287\ : Span4Mux_h
    port map (
            O => \N__80864\,
            I => \N__80820\
        );

    \I__20286\ : Span4Mux_v
    port map (
            O => \N__80859\,
            I => \N__80820\
        );

    \I__20285\ : LocalMux
    port map (
            O => \N__80856\,
            I => \N__80813\
        );

    \I__20284\ : Span4Mux_h
    port map (
            O => \N__80853\,
            I => \N__80813\
        );

    \I__20283\ : Span4Mux_v
    port map (
            O => \N__80850\,
            I => \N__80813\
        );

    \I__20282\ : LocalMux
    port map (
            O => \N__80847\,
            I => \N__80810\
        );

    \I__20281\ : Span4Mux_v
    port map (
            O => \N__80844\,
            I => \N__80807\
        );

    \I__20280\ : InMux
    port map (
            O => \N__80843\,
            I => \N__80804\
        );

    \I__20279\ : Span4Mux_h
    port map (
            O => \N__80840\,
            I => \N__80799\
        );

    \I__20278\ : Span4Mux_v
    port map (
            O => \N__80837\,
            I => \N__80799\
        );

    \I__20277\ : Sp12to4
    port map (
            O => \N__80834\,
            I => \N__80796\
        );

    \I__20276\ : LocalMux
    port map (
            O => \N__80831\,
            I => \N__80793\
        );

    \I__20275\ : Span4Mux_h
    port map (
            O => \N__80828\,
            I => \N__80790\
        );

    \I__20274\ : LocalMux
    port map (
            O => \N__80825\,
            I => \N__80787\
        );

    \I__20273\ : Span4Mux_h
    port map (
            O => \N__80820\,
            I => \N__80784\
        );

    \I__20272\ : Span4Mux_v
    port map (
            O => \N__80813\,
            I => \N__80781\
        );

    \I__20271\ : Span4Mux_v
    port map (
            O => \N__80810\,
            I => \N__80776\
        );

    \I__20270\ : Span4Mux_h
    port map (
            O => \N__80807\,
            I => \N__80776\
        );

    \I__20269\ : LocalMux
    port map (
            O => \N__80804\,
            I => \N__80769\
        );

    \I__20268\ : Sp12to4
    port map (
            O => \N__80799\,
            I => \N__80769\
        );

    \I__20267\ : Span12Mux_v
    port map (
            O => \N__80796\,
            I => \N__80769\
        );

    \I__20266\ : Span4Mux_h
    port map (
            O => \N__80793\,
            I => \N__80764\
        );

    \I__20265\ : Span4Mux_h
    port map (
            O => \N__80790\,
            I => \N__80764\
        );

    \I__20264\ : Span4Mux_v
    port map (
            O => \N__80787\,
            I => \N__80757\
        );

    \I__20263\ : Span4Mux_h
    port map (
            O => \N__80784\,
            I => \N__80757\
        );

    \I__20262\ : Span4Mux_v
    port map (
            O => \N__80781\,
            I => \N__80757\
        );

    \I__20261\ : Odrv4
    port map (
            O => \N__80776\,
            I => \c0.n17830\
        );

    \I__20260\ : Odrv12
    port map (
            O => \N__80769\,
            I => \c0.n17830\
        );

    \I__20259\ : Odrv4
    port map (
            O => \N__80764\,
            I => \c0.n17830\
        );

    \I__20258\ : Odrv4
    port map (
            O => \N__80757\,
            I => \c0.n17830\
        );

    \I__20257\ : InMux
    port map (
            O => \N__80748\,
            I => \N__80743\
        );

    \I__20256\ : CascadeMux
    port map (
            O => \N__80747\,
            I => \N__80730\
        );

    \I__20255\ : InMux
    port map (
            O => \N__80746\,
            I => \N__80726\
        );

    \I__20254\ : LocalMux
    port map (
            O => \N__80743\,
            I => \N__80723\
        );

    \I__20253\ : InMux
    port map (
            O => \N__80742\,
            I => \N__80720\
        );

    \I__20252\ : InMux
    port map (
            O => \N__80741\,
            I => \N__80715\
        );

    \I__20251\ : InMux
    port map (
            O => \N__80740\,
            I => \N__80712\
        );

    \I__20250\ : CascadeMux
    port map (
            O => \N__80739\,
            I => \N__80708\
        );

    \I__20249\ : InMux
    port map (
            O => \N__80738\,
            I => \N__80704\
        );

    \I__20248\ : InMux
    port map (
            O => \N__80737\,
            I => \N__80700\
        );

    \I__20247\ : CascadeMux
    port map (
            O => \N__80736\,
            I => \N__80697\
        );

    \I__20246\ : CascadeMux
    port map (
            O => \N__80735\,
            I => \N__80693\
        );

    \I__20245\ : InMux
    port map (
            O => \N__80734\,
            I => \N__80688\
        );

    \I__20244\ : InMux
    port map (
            O => \N__80733\,
            I => \N__80688\
        );

    \I__20243\ : InMux
    port map (
            O => \N__80730\,
            I => \N__80685\
        );

    \I__20242\ : InMux
    port map (
            O => \N__80729\,
            I => \N__80682\
        );

    \I__20241\ : LocalMux
    port map (
            O => \N__80726\,
            I => \N__80679\
        );

    \I__20240\ : Span4Mux_h
    port map (
            O => \N__80723\,
            I => \N__80674\
        );

    \I__20239\ : LocalMux
    port map (
            O => \N__80720\,
            I => \N__80674\
        );

    \I__20238\ : InMux
    port map (
            O => \N__80719\,
            I => \N__80668\
        );

    \I__20237\ : InMux
    port map (
            O => \N__80718\,
            I => \N__80665\
        );

    \I__20236\ : LocalMux
    port map (
            O => \N__80715\,
            I => \N__80662\
        );

    \I__20235\ : LocalMux
    port map (
            O => \N__80712\,
            I => \N__80659\
        );

    \I__20234\ : InMux
    port map (
            O => \N__80711\,
            I => \N__80656\
        );

    \I__20233\ : InMux
    port map (
            O => \N__80708\,
            I => \N__80650\
        );

    \I__20232\ : InMux
    port map (
            O => \N__80707\,
            I => \N__80650\
        );

    \I__20231\ : LocalMux
    port map (
            O => \N__80704\,
            I => \N__80647\
        );

    \I__20230\ : InMux
    port map (
            O => \N__80703\,
            I => \N__80644\
        );

    \I__20229\ : LocalMux
    port map (
            O => \N__80700\,
            I => \N__80641\
        );

    \I__20228\ : InMux
    port map (
            O => \N__80697\,
            I => \N__80638\
        );

    \I__20227\ : InMux
    port map (
            O => \N__80696\,
            I => \N__80635\
        );

    \I__20226\ : InMux
    port map (
            O => \N__80693\,
            I => \N__80632\
        );

    \I__20225\ : LocalMux
    port map (
            O => \N__80688\,
            I => \N__80627\
        );

    \I__20224\ : LocalMux
    port map (
            O => \N__80685\,
            I => \N__80627\
        );

    \I__20223\ : LocalMux
    port map (
            O => \N__80682\,
            I => \N__80624\
        );

    \I__20222\ : Span4Mux_v
    port map (
            O => \N__80679\,
            I => \N__80619\
        );

    \I__20221\ : Span4Mux_v
    port map (
            O => \N__80674\,
            I => \N__80619\
        );

    \I__20220\ : CascadeMux
    port map (
            O => \N__80673\,
            I => \N__80612\
        );

    \I__20219\ : InMux
    port map (
            O => \N__80672\,
            I => \N__80609\
        );

    \I__20218\ : CascadeMux
    port map (
            O => \N__80671\,
            I => \N__80606\
        );

    \I__20217\ : LocalMux
    port map (
            O => \N__80668\,
            I => \N__80602\
        );

    \I__20216\ : LocalMux
    port map (
            O => \N__80665\,
            I => \N__80595\
        );

    \I__20215\ : Span4Mux_h
    port map (
            O => \N__80662\,
            I => \N__80595\
        );

    \I__20214\ : Span4Mux_v
    port map (
            O => \N__80659\,
            I => \N__80595\
        );

    \I__20213\ : LocalMux
    port map (
            O => \N__80656\,
            I => \N__80592\
        );

    \I__20212\ : InMux
    port map (
            O => \N__80655\,
            I => \N__80589\
        );

    \I__20211\ : LocalMux
    port map (
            O => \N__80650\,
            I => \N__80586\
        );

    \I__20210\ : Span4Mux_h
    port map (
            O => \N__80647\,
            I => \N__80581\
        );

    \I__20209\ : LocalMux
    port map (
            O => \N__80644\,
            I => \N__80581\
        );

    \I__20208\ : Span4Mux_v
    port map (
            O => \N__80641\,
            I => \N__80576\
        );

    \I__20207\ : LocalMux
    port map (
            O => \N__80638\,
            I => \N__80576\
        );

    \I__20206\ : LocalMux
    port map (
            O => \N__80635\,
            I => \N__80568\
        );

    \I__20205\ : LocalMux
    port map (
            O => \N__80632\,
            I => \N__80568\
        );

    \I__20204\ : Span4Mux_v
    port map (
            O => \N__80627\,
            I => \N__80568\
        );

    \I__20203\ : Span4Mux_v
    port map (
            O => \N__80624\,
            I => \N__80565\
        );

    \I__20202\ : Span4Mux_h
    port map (
            O => \N__80619\,
            I => \N__80562\
        );

    \I__20201\ : InMux
    port map (
            O => \N__80618\,
            I => \N__80557\
        );

    \I__20200\ : InMux
    port map (
            O => \N__80617\,
            I => \N__80557\
        );

    \I__20199\ : InMux
    port map (
            O => \N__80616\,
            I => \N__80554\
        );

    \I__20198\ : InMux
    port map (
            O => \N__80615\,
            I => \N__80549\
        );

    \I__20197\ : InMux
    port map (
            O => \N__80612\,
            I => \N__80549\
        );

    \I__20196\ : LocalMux
    port map (
            O => \N__80609\,
            I => \N__80546\
        );

    \I__20195\ : InMux
    port map (
            O => \N__80606\,
            I => \N__80543\
        );

    \I__20194\ : InMux
    port map (
            O => \N__80605\,
            I => \N__80540\
        );

    \I__20193\ : Span4Mux_v
    port map (
            O => \N__80602\,
            I => \N__80535\
        );

    \I__20192\ : Span4Mux_v
    port map (
            O => \N__80595\,
            I => \N__80535\
        );

    \I__20191\ : Span4Mux_v
    port map (
            O => \N__80592\,
            I => \N__80532\
        );

    \I__20190\ : LocalMux
    port map (
            O => \N__80589\,
            I => \N__80527\
        );

    \I__20189\ : Span4Mux_v
    port map (
            O => \N__80586\,
            I => \N__80527\
        );

    \I__20188\ : Span4Mux_v
    port map (
            O => \N__80581\,
            I => \N__80524\
        );

    \I__20187\ : Span4Mux_h
    port map (
            O => \N__80576\,
            I => \N__80521\
        );

    \I__20186\ : InMux
    port map (
            O => \N__80575\,
            I => \N__80518\
        );

    \I__20185\ : Span4Mux_v
    port map (
            O => \N__80568\,
            I => \N__80515\
        );

    \I__20184\ : Span4Mux_v
    port map (
            O => \N__80565\,
            I => \N__80510\
        );

    \I__20183\ : Span4Mux_h
    port map (
            O => \N__80562\,
            I => \N__80510\
        );

    \I__20182\ : LocalMux
    port map (
            O => \N__80557\,
            I => \N__80505\
        );

    \I__20181\ : LocalMux
    port map (
            O => \N__80554\,
            I => \N__80502\
        );

    \I__20180\ : LocalMux
    port map (
            O => \N__80549\,
            I => \N__80497\
        );

    \I__20179\ : Span4Mux_v
    port map (
            O => \N__80546\,
            I => \N__80497\
        );

    \I__20178\ : LocalMux
    port map (
            O => \N__80543\,
            I => \N__80492\
        );

    \I__20177\ : LocalMux
    port map (
            O => \N__80540\,
            I => \N__80492\
        );

    \I__20176\ : Span4Mux_h
    port map (
            O => \N__80535\,
            I => \N__80487\
        );

    \I__20175\ : Span4Mux_v
    port map (
            O => \N__80532\,
            I => \N__80487\
        );

    \I__20174\ : Span4Mux_v
    port map (
            O => \N__80527\,
            I => \N__80484\
        );

    \I__20173\ : Sp12to4
    port map (
            O => \N__80524\,
            I => \N__80481\
        );

    \I__20172\ : Sp12to4
    port map (
            O => \N__80521\,
            I => \N__80478\
        );

    \I__20171\ : LocalMux
    port map (
            O => \N__80518\,
            I => \N__80471\
        );

    \I__20170\ : Sp12to4
    port map (
            O => \N__80515\,
            I => \N__80471\
        );

    \I__20169\ : Sp12to4
    port map (
            O => \N__80510\,
            I => \N__80471\
        );

    \I__20168\ : InMux
    port map (
            O => \N__80509\,
            I => \N__80466\
        );

    \I__20167\ : InMux
    port map (
            O => \N__80508\,
            I => \N__80466\
        );

    \I__20166\ : Span12Mux_h
    port map (
            O => \N__80505\,
            I => \N__80463\
        );

    \I__20165\ : Span4Mux_h
    port map (
            O => \N__80502\,
            I => \N__80458\
        );

    \I__20164\ : Span4Mux_h
    port map (
            O => \N__80497\,
            I => \N__80458\
        );

    \I__20163\ : Span4Mux_v
    port map (
            O => \N__80492\,
            I => \N__80453\
        );

    \I__20162\ : Span4Mux_v
    port map (
            O => \N__80487\,
            I => \N__80453\
        );

    \I__20161\ : Sp12to4
    port map (
            O => \N__80484\,
            I => \N__80444\
        );

    \I__20160\ : Span12Mux_h
    port map (
            O => \N__80481\,
            I => \N__80444\
        );

    \I__20159\ : Span12Mux_v
    port map (
            O => \N__80478\,
            I => \N__80444\
        );

    \I__20158\ : Span12Mux_h
    port map (
            O => \N__80471\,
            I => \N__80444\
        );

    \I__20157\ : LocalMux
    port map (
            O => \N__80466\,
            I => rx_data_0
        );

    \I__20156\ : Odrv12
    port map (
            O => \N__80463\,
            I => rx_data_0
        );

    \I__20155\ : Odrv4
    port map (
            O => \N__80458\,
            I => rx_data_0
        );

    \I__20154\ : Odrv4
    port map (
            O => \N__80453\,
            I => rx_data_0
        );

    \I__20153\ : Odrv12
    port map (
            O => \N__80444\,
            I => rx_data_0
        );

    \I__20152\ : InMux
    port map (
            O => \N__80433\,
            I => \N__80407\
        );

    \I__20151\ : InMux
    port map (
            O => \N__80432\,
            I => \N__80407\
        );

    \I__20150\ : InMux
    port map (
            O => \N__80431\,
            I => \N__80404\
        );

    \I__20149\ : InMux
    port map (
            O => \N__80430\,
            I => \N__80392\
        );

    \I__20148\ : InMux
    port map (
            O => \N__80429\,
            I => \N__80389\
        );

    \I__20147\ : InMux
    port map (
            O => \N__80428\,
            I => \N__80386\
        );

    \I__20146\ : InMux
    port map (
            O => \N__80427\,
            I => \N__80382\
        );

    \I__20145\ : InMux
    port map (
            O => \N__80426\,
            I => \N__80379\
        );

    \I__20144\ : InMux
    port map (
            O => \N__80425\,
            I => \N__80376\
        );

    \I__20143\ : InMux
    port map (
            O => \N__80424\,
            I => \N__80373\
        );

    \I__20142\ : InMux
    port map (
            O => \N__80423\,
            I => \N__80368\
        );

    \I__20141\ : InMux
    port map (
            O => \N__80422\,
            I => \N__80368\
        );

    \I__20140\ : InMux
    port map (
            O => \N__80421\,
            I => \N__80365\
        );

    \I__20139\ : InMux
    port map (
            O => \N__80420\,
            I => \N__80360\
        );

    \I__20138\ : InMux
    port map (
            O => \N__80419\,
            I => \N__80360\
        );

    \I__20137\ : InMux
    port map (
            O => \N__80418\,
            I => \N__80355\
        );

    \I__20136\ : InMux
    port map (
            O => \N__80417\,
            I => \N__80355\
        );

    \I__20135\ : InMux
    port map (
            O => \N__80416\,
            I => \N__80344\
        );

    \I__20134\ : InMux
    port map (
            O => \N__80415\,
            I => \N__80344\
        );

    \I__20133\ : InMux
    port map (
            O => \N__80414\,
            I => \N__80344\
        );

    \I__20132\ : InMux
    port map (
            O => \N__80413\,
            I => \N__80344\
        );

    \I__20131\ : InMux
    port map (
            O => \N__80412\,
            I => \N__80344\
        );

    \I__20130\ : LocalMux
    port map (
            O => \N__80407\,
            I => \N__80341\
        );

    \I__20129\ : LocalMux
    port map (
            O => \N__80404\,
            I => \N__80338\
        );

    \I__20128\ : InMux
    port map (
            O => \N__80403\,
            I => \N__80329\
        );

    \I__20127\ : InMux
    port map (
            O => \N__80402\,
            I => \N__80329\
        );

    \I__20126\ : InMux
    port map (
            O => \N__80401\,
            I => \N__80329\
        );

    \I__20125\ : InMux
    port map (
            O => \N__80400\,
            I => \N__80329\
        );

    \I__20124\ : InMux
    port map (
            O => \N__80399\,
            I => \N__80325\
        );

    \I__20123\ : InMux
    port map (
            O => \N__80398\,
            I => \N__80315\
        );

    \I__20122\ : InMux
    port map (
            O => \N__80397\,
            I => \N__80312\
        );

    \I__20121\ : InMux
    port map (
            O => \N__80396\,
            I => \N__80307\
        );

    \I__20120\ : InMux
    port map (
            O => \N__80395\,
            I => \N__80307\
        );

    \I__20119\ : LocalMux
    port map (
            O => \N__80392\,
            I => \N__80304\
        );

    \I__20118\ : LocalMux
    port map (
            O => \N__80389\,
            I => \N__80299\
        );

    \I__20117\ : LocalMux
    port map (
            O => \N__80386\,
            I => \N__80299\
        );

    \I__20116\ : InMux
    port map (
            O => \N__80385\,
            I => \N__80296\
        );

    \I__20115\ : LocalMux
    port map (
            O => \N__80382\,
            I => \N__80293\
        );

    \I__20114\ : LocalMux
    port map (
            O => \N__80379\,
            I => \N__80288\
        );

    \I__20113\ : LocalMux
    port map (
            O => \N__80376\,
            I => \N__80288\
        );

    \I__20112\ : LocalMux
    port map (
            O => \N__80373\,
            I => \N__80283\
        );

    \I__20111\ : LocalMux
    port map (
            O => \N__80368\,
            I => \N__80283\
        );

    \I__20110\ : LocalMux
    port map (
            O => \N__80365\,
            I => \N__80276\
        );

    \I__20109\ : LocalMux
    port map (
            O => \N__80360\,
            I => \N__80276\
        );

    \I__20108\ : LocalMux
    port map (
            O => \N__80355\,
            I => \N__80276\
        );

    \I__20107\ : LocalMux
    port map (
            O => \N__80344\,
            I => \N__80267\
        );

    \I__20106\ : Span4Mux_v
    port map (
            O => \N__80341\,
            I => \N__80267\
        );

    \I__20105\ : Span4Mux_v
    port map (
            O => \N__80338\,
            I => \N__80267\
        );

    \I__20104\ : LocalMux
    port map (
            O => \N__80329\,
            I => \N__80267\
        );

    \I__20103\ : InMux
    port map (
            O => \N__80328\,
            I => \N__80256\
        );

    \I__20102\ : LocalMux
    port map (
            O => \N__80325\,
            I => \N__80253\
        );

    \I__20101\ : InMux
    port map (
            O => \N__80324\,
            I => \N__80250\
        );

    \I__20100\ : InMux
    port map (
            O => \N__80323\,
            I => \N__80241\
        );

    \I__20099\ : InMux
    port map (
            O => \N__80322\,
            I => \N__80241\
        );

    \I__20098\ : InMux
    port map (
            O => \N__80321\,
            I => \N__80241\
        );

    \I__20097\ : InMux
    port map (
            O => \N__80320\,
            I => \N__80241\
        );

    \I__20096\ : InMux
    port map (
            O => \N__80319\,
            I => \N__80236\
        );

    \I__20095\ : InMux
    port map (
            O => \N__80318\,
            I => \N__80236\
        );

    \I__20094\ : LocalMux
    port map (
            O => \N__80315\,
            I => \N__80233\
        );

    \I__20093\ : LocalMux
    port map (
            O => \N__80312\,
            I => \N__80230\
        );

    \I__20092\ : LocalMux
    port map (
            O => \N__80307\,
            I => \N__80227\
        );

    \I__20091\ : Span4Mux_v
    port map (
            O => \N__80304\,
            I => \N__80224\
        );

    \I__20090\ : Span4Mux_v
    port map (
            O => \N__80299\,
            I => \N__80221\
        );

    \I__20089\ : LocalMux
    port map (
            O => \N__80296\,
            I => \N__80218\
        );

    \I__20088\ : Span4Mux_h
    port map (
            O => \N__80293\,
            I => \N__80213\
        );

    \I__20087\ : Span4Mux_v
    port map (
            O => \N__80288\,
            I => \N__80213\
        );

    \I__20086\ : Span4Mux_v
    port map (
            O => \N__80283\,
            I => \N__80206\
        );

    \I__20085\ : Span4Mux_v
    port map (
            O => \N__80276\,
            I => \N__80206\
        );

    \I__20084\ : Span4Mux_h
    port map (
            O => \N__80267\,
            I => \N__80206\
        );

    \I__20083\ : InMux
    port map (
            O => \N__80266\,
            I => \N__80203\
        );

    \I__20082\ : InMux
    port map (
            O => \N__80265\,
            I => \N__80200\
        );

    \I__20081\ : InMux
    port map (
            O => \N__80264\,
            I => \N__80197\
        );

    \I__20080\ : InMux
    port map (
            O => \N__80263\,
            I => \N__80186\
        );

    \I__20079\ : InMux
    port map (
            O => \N__80262\,
            I => \N__80186\
        );

    \I__20078\ : InMux
    port map (
            O => \N__80261\,
            I => \N__80186\
        );

    \I__20077\ : InMux
    port map (
            O => \N__80260\,
            I => \N__80186\
        );

    \I__20076\ : InMux
    port map (
            O => \N__80259\,
            I => \N__80186\
        );

    \I__20075\ : LocalMux
    port map (
            O => \N__80256\,
            I => \N__80183\
        );

    \I__20074\ : Span4Mux_h
    port map (
            O => \N__80253\,
            I => \N__80180\
        );

    \I__20073\ : LocalMux
    port map (
            O => \N__80250\,
            I => \N__80171\
        );

    \I__20072\ : LocalMux
    port map (
            O => \N__80241\,
            I => \N__80171\
        );

    \I__20071\ : LocalMux
    port map (
            O => \N__80236\,
            I => \N__80171\
        );

    \I__20070\ : Span12Mux_v
    port map (
            O => \N__80233\,
            I => \N__80171\
        );

    \I__20069\ : Span4Mux_v
    port map (
            O => \N__80230\,
            I => \N__80162\
        );

    \I__20068\ : Span4Mux_v
    port map (
            O => \N__80227\,
            I => \N__80162\
        );

    \I__20067\ : Span4Mux_h
    port map (
            O => \N__80224\,
            I => \N__80162\
        );

    \I__20066\ : Span4Mux_h
    port map (
            O => \N__80221\,
            I => \N__80162\
        );

    \I__20065\ : Span4Mux_h
    port map (
            O => \N__80218\,
            I => \N__80155\
        );

    \I__20064\ : Span4Mux_v
    port map (
            O => \N__80213\,
            I => \N__80155\
        );

    \I__20063\ : Span4Mux_h
    port map (
            O => \N__80206\,
            I => \N__80155\
        );

    \I__20062\ : LocalMux
    port map (
            O => \N__80203\,
            I => \c0.n22104\
        );

    \I__20061\ : LocalMux
    port map (
            O => \N__80200\,
            I => \c0.n22104\
        );

    \I__20060\ : LocalMux
    port map (
            O => \N__80197\,
            I => \c0.n22104\
        );

    \I__20059\ : LocalMux
    port map (
            O => \N__80186\,
            I => \c0.n22104\
        );

    \I__20058\ : Odrv4
    port map (
            O => \N__80183\,
            I => \c0.n22104\
        );

    \I__20057\ : Odrv4
    port map (
            O => \N__80180\,
            I => \c0.n22104\
        );

    \I__20056\ : Odrv12
    port map (
            O => \N__80171\,
            I => \c0.n22104\
        );

    \I__20055\ : Odrv4
    port map (
            O => \N__80162\,
            I => \c0.n22104\
        );

    \I__20054\ : Odrv4
    port map (
            O => \N__80155\,
            I => \c0.n22104\
        );

    \I__20053\ : InMux
    port map (
            O => \N__80136\,
            I => \N__80132\
        );

    \I__20052\ : InMux
    port map (
            O => \N__80135\,
            I => \N__80128\
        );

    \I__20051\ : LocalMux
    port map (
            O => \N__80132\,
            I => \N__80125\
        );

    \I__20050\ : CascadeMux
    port map (
            O => \N__80131\,
            I => \N__80122\
        );

    \I__20049\ : LocalMux
    port map (
            O => \N__80128\,
            I => \N__80119\
        );

    \I__20048\ : Span4Mux_h
    port map (
            O => \N__80125\,
            I => \N__80116\
        );

    \I__20047\ : InMux
    port map (
            O => \N__80122\,
            I => \N__80113\
        );

    \I__20046\ : Span4Mux_h
    port map (
            O => \N__80119\,
            I => \N__80110\
        );

    \I__20045\ : Span4Mux_h
    port map (
            O => \N__80116\,
            I => \N__80107\
        );

    \I__20044\ : LocalMux
    port map (
            O => \N__80113\,
            I => \c0.data_in_frame_23_0\
        );

    \I__20043\ : Odrv4
    port map (
            O => \N__80110\,
            I => \c0.data_in_frame_23_0\
        );

    \I__20042\ : Odrv4
    port map (
            O => \N__80107\,
            I => \c0.data_in_frame_23_0\
        );

    \I__20041\ : CascadeMux
    port map (
            O => \N__80100\,
            I => \N__80090\
        );

    \I__20040\ : CascadeMux
    port map (
            O => \N__80099\,
            I => \N__80087\
        );

    \I__20039\ : CascadeMux
    port map (
            O => \N__80098\,
            I => \N__80084\
        );

    \I__20038\ : CascadeMux
    port map (
            O => \N__80097\,
            I => \N__80081\
        );

    \I__20037\ : InMux
    port map (
            O => \N__80096\,
            I => \N__80076\
        );

    \I__20036\ : InMux
    port map (
            O => \N__80095\,
            I => \N__80073\
        );

    \I__20035\ : InMux
    port map (
            O => \N__80094\,
            I => \N__80070\
        );

    \I__20034\ : InMux
    port map (
            O => \N__80093\,
            I => \N__80067\
        );

    \I__20033\ : InMux
    port map (
            O => \N__80090\,
            I => \N__80064\
        );

    \I__20032\ : InMux
    port map (
            O => \N__80087\,
            I => \N__80061\
        );

    \I__20031\ : InMux
    port map (
            O => \N__80084\,
            I => \N__80055\
        );

    \I__20030\ : InMux
    port map (
            O => \N__80081\,
            I => \N__80055\
        );

    \I__20029\ : CascadeMux
    port map (
            O => \N__80080\,
            I => \N__80052\
        );

    \I__20028\ : InMux
    port map (
            O => \N__80079\,
            I => \N__80048\
        );

    \I__20027\ : LocalMux
    port map (
            O => \N__80076\,
            I => \N__80045\
        );

    \I__20026\ : LocalMux
    port map (
            O => \N__80073\,
            I => \N__80041\
        );

    \I__20025\ : LocalMux
    port map (
            O => \N__80070\,
            I => \N__80036\
        );

    \I__20024\ : LocalMux
    port map (
            O => \N__80067\,
            I => \N__80036\
        );

    \I__20023\ : LocalMux
    port map (
            O => \N__80064\,
            I => \N__80033\
        );

    \I__20022\ : LocalMux
    port map (
            O => \N__80061\,
            I => \N__80026\
        );

    \I__20021\ : InMux
    port map (
            O => \N__80060\,
            I => \N__80023\
        );

    \I__20020\ : LocalMux
    port map (
            O => \N__80055\,
            I => \N__80020\
        );

    \I__20019\ : InMux
    port map (
            O => \N__80052\,
            I => \N__80017\
        );

    \I__20018\ : InMux
    port map (
            O => \N__80051\,
            I => \N__80013\
        );

    \I__20017\ : LocalMux
    port map (
            O => \N__80048\,
            I => \N__80010\
        );

    \I__20016\ : Span4Mux_h
    port map (
            O => \N__80045\,
            I => \N__80004\
        );

    \I__20015\ : InMux
    port map (
            O => \N__80044\,
            I => \N__80001\
        );

    \I__20014\ : Span4Mux_h
    port map (
            O => \N__80041\,
            I => \N__79998\
        );

    \I__20013\ : Span4Mux_v
    port map (
            O => \N__80036\,
            I => \N__79995\
        );

    \I__20012\ : Span4Mux_h
    port map (
            O => \N__80033\,
            I => \N__79992\
        );

    \I__20011\ : CascadeMux
    port map (
            O => \N__80032\,
            I => \N__79989\
        );

    \I__20010\ : InMux
    port map (
            O => \N__80031\,
            I => \N__79980\
        );

    \I__20009\ : InMux
    port map (
            O => \N__80030\,
            I => \N__79975\
        );

    \I__20008\ : InMux
    port map (
            O => \N__80029\,
            I => \N__79975\
        );

    \I__20007\ : Span4Mux_h
    port map (
            O => \N__80026\,
            I => \N__79972\
        );

    \I__20006\ : LocalMux
    port map (
            O => \N__80023\,
            I => \N__79967\
        );

    \I__20005\ : Span4Mux_v
    port map (
            O => \N__80020\,
            I => \N__79967\
        );

    \I__20004\ : LocalMux
    port map (
            O => \N__80017\,
            I => \N__79964\
        );

    \I__20003\ : InMux
    port map (
            O => \N__80016\,
            I => \N__79961\
        );

    \I__20002\ : LocalMux
    port map (
            O => \N__80013\,
            I => \N__79958\
        );

    \I__20001\ : Span4Mux_h
    port map (
            O => \N__80010\,
            I => \N__79955\
        );

    \I__20000\ : CascadeMux
    port map (
            O => \N__80009\,
            I => \N__79949\
        );

    \I__19999\ : InMux
    port map (
            O => \N__80008\,
            I => \N__79944\
        );

    \I__19998\ : InMux
    port map (
            O => \N__80007\,
            I => \N__79941\
        );

    \I__19997\ : Span4Mux_h
    port map (
            O => \N__80004\,
            I => \N__79938\
        );

    \I__19996\ : LocalMux
    port map (
            O => \N__80001\,
            I => \N__79929\
        );

    \I__19995\ : Span4Mux_h
    port map (
            O => \N__79998\,
            I => \N__79929\
        );

    \I__19994\ : Span4Mux_h
    port map (
            O => \N__79995\,
            I => \N__79929\
        );

    \I__19993\ : Span4Mux_v
    port map (
            O => \N__79992\,
            I => \N__79929\
        );

    \I__19992\ : InMux
    port map (
            O => \N__79989\,
            I => \N__79922\
        );

    \I__19991\ : InMux
    port map (
            O => \N__79988\,
            I => \N__79922\
        );

    \I__19990\ : InMux
    port map (
            O => \N__79987\,
            I => \N__79922\
        );

    \I__19989\ : InMux
    port map (
            O => \N__79986\,
            I => \N__79919\
        );

    \I__19988\ : InMux
    port map (
            O => \N__79985\,
            I => \N__79914\
        );

    \I__19987\ : InMux
    port map (
            O => \N__79984\,
            I => \N__79914\
        );

    \I__19986\ : InMux
    port map (
            O => \N__79983\,
            I => \N__79911\
        );

    \I__19985\ : LocalMux
    port map (
            O => \N__79980\,
            I => \N__79908\
        );

    \I__19984\ : LocalMux
    port map (
            O => \N__79975\,
            I => \N__79901\
        );

    \I__19983\ : Span4Mux_h
    port map (
            O => \N__79972\,
            I => \N__79901\
        );

    \I__19982\ : Span4Mux_h
    port map (
            O => \N__79967\,
            I => \N__79901\
        );

    \I__19981\ : Span4Mux_v
    port map (
            O => \N__79964\,
            I => \N__79892\
        );

    \I__19980\ : LocalMux
    port map (
            O => \N__79961\,
            I => \N__79892\
        );

    \I__19979\ : Span4Mux_h
    port map (
            O => \N__79958\,
            I => \N__79892\
        );

    \I__19978\ : Span4Mux_v
    port map (
            O => \N__79955\,
            I => \N__79892\
        );

    \I__19977\ : CascadeMux
    port map (
            O => \N__79954\,
            I => \N__79889\
        );

    \I__19976\ : InMux
    port map (
            O => \N__79953\,
            I => \N__79886\
        );

    \I__19975\ : InMux
    port map (
            O => \N__79952\,
            I => \N__79883\
        );

    \I__19974\ : InMux
    port map (
            O => \N__79949\,
            I => \N__79878\
        );

    \I__19973\ : InMux
    port map (
            O => \N__79948\,
            I => \N__79878\
        );

    \I__19972\ : InMux
    port map (
            O => \N__79947\,
            I => \N__79875\
        );

    \I__19971\ : LocalMux
    port map (
            O => \N__79944\,
            I => \N__79868\
        );

    \I__19970\ : LocalMux
    port map (
            O => \N__79941\,
            I => \N__79868\
        );

    \I__19969\ : Span4Mux_h
    port map (
            O => \N__79938\,
            I => \N__79868\
        );

    \I__19968\ : Span4Mux_v
    port map (
            O => \N__79929\,
            I => \N__79865\
        );

    \I__19967\ : LocalMux
    port map (
            O => \N__79922\,
            I => \N__79860\
        );

    \I__19966\ : LocalMux
    port map (
            O => \N__79919\,
            I => \N__79860\
        );

    \I__19965\ : LocalMux
    port map (
            O => \N__79914\,
            I => \N__79857\
        );

    \I__19964\ : LocalMux
    port map (
            O => \N__79911\,
            I => \N__79848\
        );

    \I__19963\ : Span12Mux_s10_v
    port map (
            O => \N__79908\,
            I => \N__79848\
        );

    \I__19962\ : Sp12to4
    port map (
            O => \N__79901\,
            I => \N__79848\
        );

    \I__19961\ : Sp12to4
    port map (
            O => \N__79892\,
            I => \N__79848\
        );

    \I__19960\ : InMux
    port map (
            O => \N__79889\,
            I => \N__79845\
        );

    \I__19959\ : LocalMux
    port map (
            O => \N__79886\,
            I => \N__79842\
        );

    \I__19958\ : LocalMux
    port map (
            O => \N__79883\,
            I => \N__79833\
        );

    \I__19957\ : LocalMux
    port map (
            O => \N__79878\,
            I => \N__79833\
        );

    \I__19956\ : LocalMux
    port map (
            O => \N__79875\,
            I => \N__79833\
        );

    \I__19955\ : Span4Mux_v
    port map (
            O => \N__79868\,
            I => \N__79833\
        );

    \I__19954\ : Span4Mux_v
    port map (
            O => \N__79865\,
            I => \N__79830\
        );

    \I__19953\ : Span4Mux_v
    port map (
            O => \N__79860\,
            I => \N__79827\
        );

    \I__19952\ : Span12Mux_v
    port map (
            O => \N__79857\,
            I => \N__79824\
        );

    \I__19951\ : Span12Mux_v
    port map (
            O => \N__79848\,
            I => \N__79821\
        );

    \I__19950\ : LocalMux
    port map (
            O => \N__79845\,
            I => \N__79814\
        );

    \I__19949\ : Span4Mux_h
    port map (
            O => \N__79842\,
            I => \N__79814\
        );

    \I__19948\ : Span4Mux_v
    port map (
            O => \N__79833\,
            I => \N__79814\
        );

    \I__19947\ : Span4Mux_v
    port map (
            O => \N__79830\,
            I => \N__79811\
        );

    \I__19946\ : Odrv4
    port map (
            O => \N__79827\,
            I => \c0.n9_adj_4552\
        );

    \I__19945\ : Odrv12
    port map (
            O => \N__79824\,
            I => \c0.n9_adj_4552\
        );

    \I__19944\ : Odrv12
    port map (
            O => \N__79821\,
            I => \c0.n9_adj_4552\
        );

    \I__19943\ : Odrv4
    port map (
            O => \N__79814\,
            I => \c0.n9_adj_4552\
        );

    \I__19942\ : Odrv4
    port map (
            O => \N__79811\,
            I => \c0.n9_adj_4552\
        );

    \I__19941\ : CascadeMux
    port map (
            O => \N__79800\,
            I => \N__79797\
        );

    \I__19940\ : InMux
    port map (
            O => \N__79797\,
            I => \N__79793\
        );

    \I__19939\ : CascadeMux
    port map (
            O => \N__79796\,
            I => \N__79788\
        );

    \I__19938\ : LocalMux
    port map (
            O => \N__79793\,
            I => \N__79781\
        );

    \I__19937\ : InMux
    port map (
            O => \N__79792\,
            I => \N__79778\
        );

    \I__19936\ : InMux
    port map (
            O => \N__79791\,
            I => \N__79769\
        );

    \I__19935\ : InMux
    port map (
            O => \N__79788\,
            I => \N__79769\
        );

    \I__19934\ : InMux
    port map (
            O => \N__79787\,
            I => \N__79769\
        );

    \I__19933\ : InMux
    port map (
            O => \N__79786\,
            I => \N__79766\
        );

    \I__19932\ : InMux
    port map (
            O => \N__79785\,
            I => \N__79763\
        );

    \I__19931\ : InMux
    port map (
            O => \N__79784\,
            I => \N__79760\
        );

    \I__19930\ : Span4Mux_h
    port map (
            O => \N__79781\,
            I => \N__79751\
        );

    \I__19929\ : LocalMux
    port map (
            O => \N__79778\,
            I => \N__79751\
        );

    \I__19928\ : InMux
    port map (
            O => \N__79777\,
            I => \N__79746\
        );

    \I__19927\ : InMux
    port map (
            O => \N__79776\,
            I => \N__79746\
        );

    \I__19926\ : LocalMux
    port map (
            O => \N__79769\,
            I => \N__79743\
        );

    \I__19925\ : LocalMux
    port map (
            O => \N__79766\,
            I => \N__79740\
        );

    \I__19924\ : LocalMux
    port map (
            O => \N__79763\,
            I => \N__79737\
        );

    \I__19923\ : LocalMux
    port map (
            O => \N__79760\,
            I => \N__79734\
        );

    \I__19922\ : InMux
    port map (
            O => \N__79759\,
            I => \N__79729\
        );

    \I__19921\ : InMux
    port map (
            O => \N__79758\,
            I => \N__79729\
        );

    \I__19920\ : InMux
    port map (
            O => \N__79757\,
            I => \N__79724\
        );

    \I__19919\ : CascadeMux
    port map (
            O => \N__79756\,
            I => \N__79721\
        );

    \I__19918\ : Span4Mux_v
    port map (
            O => \N__79751\,
            I => \N__79718\
        );

    \I__19917\ : LocalMux
    port map (
            O => \N__79746\,
            I => \N__79709\
        );

    \I__19916\ : Span4Mux_v
    port map (
            O => \N__79743\,
            I => \N__79709\
        );

    \I__19915\ : Span4Mux_h
    port map (
            O => \N__79740\,
            I => \N__79709\
        );

    \I__19914\ : Span4Mux_v
    port map (
            O => \N__79737\,
            I => \N__79709\
        );

    \I__19913\ : Span4Mux_h
    port map (
            O => \N__79734\,
            I => \N__79704\
        );

    \I__19912\ : LocalMux
    port map (
            O => \N__79729\,
            I => \N__79704\
        );

    \I__19911\ : CascadeMux
    port map (
            O => \N__79728\,
            I => \N__79699\
        );

    \I__19910\ : InMux
    port map (
            O => \N__79727\,
            I => \N__79695\
        );

    \I__19909\ : LocalMux
    port map (
            O => \N__79724\,
            I => \N__79692\
        );

    \I__19908\ : InMux
    port map (
            O => \N__79721\,
            I => \N__79689\
        );

    \I__19907\ : Span4Mux_h
    port map (
            O => \N__79718\,
            I => \N__79686\
        );

    \I__19906\ : Span4Mux_h
    port map (
            O => \N__79709\,
            I => \N__79681\
        );

    \I__19905\ : Span4Mux_v
    port map (
            O => \N__79704\,
            I => \N__79681\
        );

    \I__19904\ : InMux
    port map (
            O => \N__79703\,
            I => \N__79678\
        );

    \I__19903\ : InMux
    port map (
            O => \N__79702\,
            I => \N__79674\
        );

    \I__19902\ : InMux
    port map (
            O => \N__79699\,
            I => \N__79671\
        );

    \I__19901\ : InMux
    port map (
            O => \N__79698\,
            I => \N__79668\
        );

    \I__19900\ : LocalMux
    port map (
            O => \N__79695\,
            I => \N__79665\
        );

    \I__19899\ : Span4Mux_h
    port map (
            O => \N__79692\,
            I => \N__79662\
        );

    \I__19898\ : LocalMux
    port map (
            O => \N__79689\,
            I => \N__79653\
        );

    \I__19897\ : Span4Mux_h
    port map (
            O => \N__79686\,
            I => \N__79653\
        );

    \I__19896\ : Span4Mux_h
    port map (
            O => \N__79681\,
            I => \N__79653\
        );

    \I__19895\ : LocalMux
    port map (
            O => \N__79678\,
            I => \N__79653\
        );

    \I__19894\ : CascadeMux
    port map (
            O => \N__79677\,
            I => \N__79650\
        );

    \I__19893\ : LocalMux
    port map (
            O => \N__79674\,
            I => \N__79641\
        );

    \I__19892\ : LocalMux
    port map (
            O => \N__79671\,
            I => \N__79641\
        );

    \I__19891\ : LocalMux
    port map (
            O => \N__79668\,
            I => \N__79632\
        );

    \I__19890\ : Span4Mux_h
    port map (
            O => \N__79665\,
            I => \N__79632\
        );

    \I__19889\ : Span4Mux_v
    port map (
            O => \N__79662\,
            I => \N__79632\
        );

    \I__19888\ : Span4Mux_v
    port map (
            O => \N__79653\,
            I => \N__79632\
        );

    \I__19887\ : InMux
    port map (
            O => \N__79650\,
            I => \N__79629\
        );

    \I__19886\ : CascadeMux
    port map (
            O => \N__79649\,
            I => \N__79623\
        );

    \I__19885\ : InMux
    port map (
            O => \N__79648\,
            I => \N__79619\
        );

    \I__19884\ : InMux
    port map (
            O => \N__79647\,
            I => \N__79616\
        );

    \I__19883\ : InMux
    port map (
            O => \N__79646\,
            I => \N__79613\
        );

    \I__19882\ : Span4Mux_v
    port map (
            O => \N__79641\,
            I => \N__79608\
        );

    \I__19881\ : Span4Mux_v
    port map (
            O => \N__79632\,
            I => \N__79608\
        );

    \I__19880\ : LocalMux
    port map (
            O => \N__79629\,
            I => \N__79605\
        );

    \I__19879\ : InMux
    port map (
            O => \N__79628\,
            I => \N__79602\
        );

    \I__19878\ : InMux
    port map (
            O => \N__79627\,
            I => \N__79599\
        );

    \I__19877\ : InMux
    port map (
            O => \N__79626\,
            I => \N__79596\
        );

    \I__19876\ : InMux
    port map (
            O => \N__79623\,
            I => \N__79593\
        );

    \I__19875\ : InMux
    port map (
            O => \N__79622\,
            I => \N__79590\
        );

    \I__19874\ : LocalMux
    port map (
            O => \N__79619\,
            I => \N__79582\
        );

    \I__19873\ : LocalMux
    port map (
            O => \N__79616\,
            I => \N__79582\
        );

    \I__19872\ : LocalMux
    port map (
            O => \N__79613\,
            I => \N__79579\
        );

    \I__19871\ : Span4Mux_h
    port map (
            O => \N__79608\,
            I => \N__79576\
        );

    \I__19870\ : Span4Mux_h
    port map (
            O => \N__79605\,
            I => \N__79571\
        );

    \I__19869\ : LocalMux
    port map (
            O => \N__79602\,
            I => \N__79571\
        );

    \I__19868\ : LocalMux
    port map (
            O => \N__79599\,
            I => \N__79568\
        );

    \I__19867\ : LocalMux
    port map (
            O => \N__79596\,
            I => \N__79565\
        );

    \I__19866\ : LocalMux
    port map (
            O => \N__79593\,
            I => \N__79560\
        );

    \I__19865\ : LocalMux
    port map (
            O => \N__79590\,
            I => \N__79560\
        );

    \I__19864\ : InMux
    port map (
            O => \N__79589\,
            I => \N__79557\
        );

    \I__19863\ : InMux
    port map (
            O => \N__79588\,
            I => \N__79554\
        );

    \I__19862\ : InMux
    port map (
            O => \N__79587\,
            I => \N__79551\
        );

    \I__19861\ : Span12Mux_h
    port map (
            O => \N__79582\,
            I => \N__79548\
        );

    \I__19860\ : Span4Mux_h
    port map (
            O => \N__79579\,
            I => \N__79543\
        );

    \I__19859\ : Span4Mux_v
    port map (
            O => \N__79576\,
            I => \N__79543\
        );

    \I__19858\ : Sp12to4
    port map (
            O => \N__79571\,
            I => \N__79537\
        );

    \I__19857\ : Span12Mux_v
    port map (
            O => \N__79568\,
            I => \N__79537\
        );

    \I__19856\ : Span12Mux_h
    port map (
            O => \N__79565\,
            I => \N__79532\
        );

    \I__19855\ : Sp12to4
    port map (
            O => \N__79560\,
            I => \N__79532\
        );

    \I__19854\ : LocalMux
    port map (
            O => \N__79557\,
            I => \N__79527\
        );

    \I__19853\ : LocalMux
    port map (
            O => \N__79554\,
            I => \N__79527\
        );

    \I__19852\ : LocalMux
    port map (
            O => \N__79551\,
            I => \N__79522\
        );

    \I__19851\ : Span12Mux_v
    port map (
            O => \N__79548\,
            I => \N__79522\
        );

    \I__19850\ : Span4Mux_v
    port map (
            O => \N__79543\,
            I => \N__79519\
        );

    \I__19849\ : InMux
    port map (
            O => \N__79542\,
            I => \N__79516\
        );

    \I__19848\ : Span12Mux_v
    port map (
            O => \N__79537\,
            I => \N__79513\
        );

    \I__19847\ : Span12Mux_v
    port map (
            O => \N__79532\,
            I => \N__79510\
        );

    \I__19846\ : Span12Mux_h
    port map (
            O => \N__79527\,
            I => \N__79505\
        );

    \I__19845\ : Span12Mux_h
    port map (
            O => \N__79522\,
            I => \N__79505\
        );

    \I__19844\ : Span4Mux_v
    port map (
            O => \N__79519\,
            I => \N__79502\
        );

    \I__19843\ : LocalMux
    port map (
            O => \N__79516\,
            I => rx_data_5
        );

    \I__19842\ : Odrv12
    port map (
            O => \N__79513\,
            I => rx_data_5
        );

    \I__19841\ : Odrv12
    port map (
            O => \N__79510\,
            I => rx_data_5
        );

    \I__19840\ : Odrv12
    port map (
            O => \N__79505\,
            I => rx_data_5
        );

    \I__19839\ : Odrv4
    port map (
            O => \N__79502\,
            I => rx_data_5
        );

    \I__19838\ : InMux
    port map (
            O => \N__79491\,
            I => \N__79485\
        );

    \I__19837\ : InMux
    port map (
            O => \N__79490\,
            I => \N__79478\
        );

    \I__19836\ : InMux
    port map (
            O => \N__79489\,
            I => \N__79473\
        );

    \I__19835\ : InMux
    port map (
            O => \N__79488\,
            I => \N__79468\
        );

    \I__19834\ : LocalMux
    port map (
            O => \N__79485\,
            I => \N__79465\
        );

    \I__19833\ : InMux
    port map (
            O => \N__79484\,
            I => \N__79458\
        );

    \I__19832\ : InMux
    port map (
            O => \N__79483\,
            I => \N__79458\
        );

    \I__19831\ : InMux
    port map (
            O => \N__79482\,
            I => \N__79453\
        );

    \I__19830\ : InMux
    port map (
            O => \N__79481\,
            I => \N__79450\
        );

    \I__19829\ : LocalMux
    port map (
            O => \N__79478\,
            I => \N__79447\
        );

    \I__19828\ : CascadeMux
    port map (
            O => \N__79477\,
            I => \N__79444\
        );

    \I__19827\ : InMux
    port map (
            O => \N__79476\,
            I => \N__79436\
        );

    \I__19826\ : LocalMux
    port map (
            O => \N__79473\,
            I => \N__79433\
        );

    \I__19825\ : InMux
    port map (
            O => \N__79472\,
            I => \N__79428\
        );

    \I__19824\ : InMux
    port map (
            O => \N__79471\,
            I => \N__79428\
        );

    \I__19823\ : LocalMux
    port map (
            O => \N__79468\,
            I => \N__79425\
        );

    \I__19822\ : Span4Mux_h
    port map (
            O => \N__79465\,
            I => \N__79422\
        );

    \I__19821\ : InMux
    port map (
            O => \N__79464\,
            I => \N__79415\
        );

    \I__19820\ : InMux
    port map (
            O => \N__79463\,
            I => \N__79415\
        );

    \I__19819\ : LocalMux
    port map (
            O => \N__79458\,
            I => \N__79412\
        );

    \I__19818\ : InMux
    port map (
            O => \N__79457\,
            I => \N__79407\
        );

    \I__19817\ : InMux
    port map (
            O => \N__79456\,
            I => \N__79407\
        );

    \I__19816\ : LocalMux
    port map (
            O => \N__79453\,
            I => \N__79404\
        );

    \I__19815\ : LocalMux
    port map (
            O => \N__79450\,
            I => \N__79399\
        );

    \I__19814\ : Span4Mux_v
    port map (
            O => \N__79447\,
            I => \N__79399\
        );

    \I__19813\ : InMux
    port map (
            O => \N__79444\,
            I => \N__79393\
        );

    \I__19812\ : InMux
    port map (
            O => \N__79443\,
            I => \N__79388\
        );

    \I__19811\ : InMux
    port map (
            O => \N__79442\,
            I => \N__79388\
        );

    \I__19810\ : InMux
    port map (
            O => \N__79441\,
            I => \N__79385\
        );

    \I__19809\ : InMux
    port map (
            O => \N__79440\,
            I => \N__79380\
        );

    \I__19808\ : InMux
    port map (
            O => \N__79439\,
            I => \N__79380\
        );

    \I__19807\ : LocalMux
    port map (
            O => \N__79436\,
            I => \N__79373\
        );

    \I__19806\ : Span4Mux_v
    port map (
            O => \N__79433\,
            I => \N__79373\
        );

    \I__19805\ : LocalMux
    port map (
            O => \N__79428\,
            I => \N__79373\
        );

    \I__19804\ : Span4Mux_v
    port map (
            O => \N__79425\,
            I => \N__79370\
        );

    \I__19803\ : Span4Mux_v
    port map (
            O => \N__79422\,
            I => \N__79367\
        );

    \I__19802\ : InMux
    port map (
            O => \N__79421\,
            I => \N__79351\
        );

    \I__19801\ : InMux
    port map (
            O => \N__79420\,
            I => \N__79348\
        );

    \I__19800\ : LocalMux
    port map (
            O => \N__79415\,
            I => \N__79345\
        );

    \I__19799\ : Span12Mux_s7_v
    port map (
            O => \N__79412\,
            I => \N__79342\
        );

    \I__19798\ : LocalMux
    port map (
            O => \N__79407\,
            I => \N__79337\
        );

    \I__19797\ : Span4Mux_v
    port map (
            O => \N__79404\,
            I => \N__79337\
        );

    \I__19796\ : Span4Mux_h
    port map (
            O => \N__79399\,
            I => \N__79334\
        );

    \I__19795\ : InMux
    port map (
            O => \N__79398\,
            I => \N__79327\
        );

    \I__19794\ : InMux
    port map (
            O => \N__79397\,
            I => \N__79327\
        );

    \I__19793\ : InMux
    port map (
            O => \N__79396\,
            I => \N__79327\
        );

    \I__19792\ : LocalMux
    port map (
            O => \N__79393\,
            I => \N__79324\
        );

    \I__19791\ : LocalMux
    port map (
            O => \N__79388\,
            I => \N__79321\
        );

    \I__19790\ : LocalMux
    port map (
            O => \N__79385\,
            I => \N__79316\
        );

    \I__19789\ : LocalMux
    port map (
            O => \N__79380\,
            I => \N__79316\
        );

    \I__19788\ : Span4Mux_v
    port map (
            O => \N__79373\,
            I => \N__79311\
        );

    \I__19787\ : Span4Mux_h
    port map (
            O => \N__79370\,
            I => \N__79311\
        );

    \I__19786\ : Span4Mux_v
    port map (
            O => \N__79367\,
            I => \N__79308\
        );

    \I__19785\ : InMux
    port map (
            O => \N__79366\,
            I => \N__79305\
        );

    \I__19784\ : InMux
    port map (
            O => \N__79365\,
            I => \N__79300\
        );

    \I__19783\ : InMux
    port map (
            O => \N__79364\,
            I => \N__79300\
        );

    \I__19782\ : InMux
    port map (
            O => \N__79363\,
            I => \N__79295\
        );

    \I__19781\ : InMux
    port map (
            O => \N__79362\,
            I => \N__79295\
        );

    \I__19780\ : InMux
    port map (
            O => \N__79361\,
            I => \N__79288\
        );

    \I__19779\ : InMux
    port map (
            O => \N__79360\,
            I => \N__79288\
        );

    \I__19778\ : InMux
    port map (
            O => \N__79359\,
            I => \N__79288\
        );

    \I__19777\ : InMux
    port map (
            O => \N__79358\,
            I => \N__79277\
        );

    \I__19776\ : InMux
    port map (
            O => \N__79357\,
            I => \N__79277\
        );

    \I__19775\ : InMux
    port map (
            O => \N__79356\,
            I => \N__79277\
        );

    \I__19774\ : InMux
    port map (
            O => \N__79355\,
            I => \N__79277\
        );

    \I__19773\ : InMux
    port map (
            O => \N__79354\,
            I => \N__79277\
        );

    \I__19772\ : LocalMux
    port map (
            O => \N__79351\,
            I => \N__79274\
        );

    \I__19771\ : LocalMux
    port map (
            O => \N__79348\,
            I => \N__79269\
        );

    \I__19770\ : Span4Mux_v
    port map (
            O => \N__79345\,
            I => \N__79269\
        );

    \I__19769\ : Span12Mux_v
    port map (
            O => \N__79342\,
            I => \N__79266\
        );

    \I__19768\ : Span4Mux_h
    port map (
            O => \N__79337\,
            I => \N__79261\
        );

    \I__19767\ : Span4Mux_h
    port map (
            O => \N__79334\,
            I => \N__79261\
        );

    \I__19766\ : LocalMux
    port map (
            O => \N__79327\,
            I => \N__79248\
        );

    \I__19765\ : Span4Mux_v
    port map (
            O => \N__79324\,
            I => \N__79248\
        );

    \I__19764\ : Span4Mux_h
    port map (
            O => \N__79321\,
            I => \N__79248\
        );

    \I__19763\ : Span4Mux_v
    port map (
            O => \N__79316\,
            I => \N__79248\
        );

    \I__19762\ : Span4Mux_h
    port map (
            O => \N__79311\,
            I => \N__79248\
        );

    \I__19761\ : Span4Mux_h
    port map (
            O => \N__79308\,
            I => \N__79248\
        );

    \I__19760\ : LocalMux
    port map (
            O => \N__79305\,
            I => \c0.n22134\
        );

    \I__19759\ : LocalMux
    port map (
            O => \N__79300\,
            I => \c0.n22134\
        );

    \I__19758\ : LocalMux
    port map (
            O => \N__79295\,
            I => \c0.n22134\
        );

    \I__19757\ : LocalMux
    port map (
            O => \N__79288\,
            I => \c0.n22134\
        );

    \I__19756\ : LocalMux
    port map (
            O => \N__79277\,
            I => \c0.n22134\
        );

    \I__19755\ : Odrv4
    port map (
            O => \N__79274\,
            I => \c0.n22134\
        );

    \I__19754\ : Odrv4
    port map (
            O => \N__79269\,
            I => \c0.n22134\
        );

    \I__19753\ : Odrv12
    port map (
            O => \N__79266\,
            I => \c0.n22134\
        );

    \I__19752\ : Odrv4
    port map (
            O => \N__79261\,
            I => \c0.n22134\
        );

    \I__19751\ : Odrv4
    port map (
            O => \N__79248\,
            I => \c0.n22134\
        );

    \I__19750\ : CascadeMux
    port map (
            O => \N__79227\,
            I => \N__79223\
        );

    \I__19749\ : InMux
    port map (
            O => \N__79226\,
            I => \N__79220\
        );

    \I__19748\ : InMux
    port map (
            O => \N__79223\,
            I => \N__79217\
        );

    \I__19747\ : LocalMux
    port map (
            O => \N__79220\,
            I => \N__79214\
        );

    \I__19746\ : LocalMux
    port map (
            O => \N__79217\,
            I => \c0.data_in_frame_28_5\
        );

    \I__19745\ : Odrv4
    port map (
            O => \N__79214\,
            I => \c0.data_in_frame_28_5\
        );

    \I__19744\ : InMux
    port map (
            O => \N__79209\,
            I => \N__79206\
        );

    \I__19743\ : LocalMux
    port map (
            O => \N__79206\,
            I => \N__79200\
        );

    \I__19742\ : InMux
    port map (
            O => \N__79205\,
            I => \N__79197\
        );

    \I__19741\ : CascadeMux
    port map (
            O => \N__79204\,
            I => \N__79194\
        );

    \I__19740\ : InMux
    port map (
            O => \N__79203\,
            I => \N__79186\
        );

    \I__19739\ : Span4Mux_h
    port map (
            O => \N__79200\,
            I => \N__79177\
        );

    \I__19738\ : LocalMux
    port map (
            O => \N__79197\,
            I => \N__79177\
        );

    \I__19737\ : InMux
    port map (
            O => \N__79194\,
            I => \N__79174\
        );

    \I__19736\ : CascadeMux
    port map (
            O => \N__79193\,
            I => \N__79169\
        );

    \I__19735\ : InMux
    port map (
            O => \N__79192\,
            I => \N__79164\
        );

    \I__19734\ : CascadeMux
    port map (
            O => \N__79191\,
            I => \N__79161\
        );

    \I__19733\ : InMux
    port map (
            O => \N__79190\,
            I => \N__79158\
        );

    \I__19732\ : InMux
    port map (
            O => \N__79189\,
            I => \N__79155\
        );

    \I__19731\ : LocalMux
    port map (
            O => \N__79186\,
            I => \N__79152\
        );

    \I__19730\ : InMux
    port map (
            O => \N__79185\,
            I => \N__79149\
        );

    \I__19729\ : CascadeMux
    port map (
            O => \N__79184\,
            I => \N__79145\
        );

    \I__19728\ : CascadeMux
    port map (
            O => \N__79183\,
            I => \N__79142\
        );

    \I__19727\ : CascadeMux
    port map (
            O => \N__79182\,
            I => \N__79137\
        );

    \I__19726\ : Span4Mux_v
    port map (
            O => \N__79177\,
            I => \N__79132\
        );

    \I__19725\ : LocalMux
    port map (
            O => \N__79174\,
            I => \N__79132\
        );

    \I__19724\ : InMux
    port map (
            O => \N__79173\,
            I => \N__79129\
        );

    \I__19723\ : InMux
    port map (
            O => \N__79172\,
            I => \N__79126\
        );

    \I__19722\ : InMux
    port map (
            O => \N__79169\,
            I => \N__79120\
        );

    \I__19721\ : InMux
    port map (
            O => \N__79168\,
            I => \N__79120\
        );

    \I__19720\ : InMux
    port map (
            O => \N__79167\,
            I => \N__79117\
        );

    \I__19719\ : LocalMux
    port map (
            O => \N__79164\,
            I => \N__79114\
        );

    \I__19718\ : InMux
    port map (
            O => \N__79161\,
            I => \N__79111\
        );

    \I__19717\ : LocalMux
    port map (
            O => \N__79158\,
            I => \N__79101\
        );

    \I__19716\ : LocalMux
    port map (
            O => \N__79155\,
            I => \N__79101\
        );

    \I__19715\ : Span4Mux_h
    port map (
            O => \N__79152\,
            I => \N__79096\
        );

    \I__19714\ : LocalMux
    port map (
            O => \N__79149\,
            I => \N__79096\
        );

    \I__19713\ : InMux
    port map (
            O => \N__79148\,
            I => \N__79093\
        );

    \I__19712\ : InMux
    port map (
            O => \N__79145\,
            I => \N__79088\
        );

    \I__19711\ : InMux
    port map (
            O => \N__79142\,
            I => \N__79088\
        );

    \I__19710\ : CascadeMux
    port map (
            O => \N__79141\,
            I => \N__79085\
        );

    \I__19709\ : InMux
    port map (
            O => \N__79140\,
            I => \N__79078\
        );

    \I__19708\ : InMux
    port map (
            O => \N__79137\,
            I => \N__79078\
        );

    \I__19707\ : Span4Mux_h
    port map (
            O => \N__79132\,
            I => \N__79075\
        );

    \I__19706\ : LocalMux
    port map (
            O => \N__79129\,
            I => \N__79072\
        );

    \I__19705\ : LocalMux
    port map (
            O => \N__79126\,
            I => \N__79069\
        );

    \I__19704\ : InMux
    port map (
            O => \N__79125\,
            I => \N__79066\
        );

    \I__19703\ : LocalMux
    port map (
            O => \N__79120\,
            I => \N__79063\
        );

    \I__19702\ : LocalMux
    port map (
            O => \N__79117\,
            I => \N__79060\
        );

    \I__19701\ : Span4Mux_v
    port map (
            O => \N__79114\,
            I => \N__79055\
        );

    \I__19700\ : LocalMux
    port map (
            O => \N__79111\,
            I => \N__79055\
        );

    \I__19699\ : InMux
    port map (
            O => \N__79110\,
            I => \N__79052\
        );

    \I__19698\ : InMux
    port map (
            O => \N__79109\,
            I => \N__79046\
        );

    \I__19697\ : InMux
    port map (
            O => \N__79108\,
            I => \N__79046\
        );

    \I__19696\ : InMux
    port map (
            O => \N__79107\,
            I => \N__79043\
        );

    \I__19695\ : InMux
    port map (
            O => \N__79106\,
            I => \N__79040\
        );

    \I__19694\ : Span4Mux_v
    port map (
            O => \N__79101\,
            I => \N__79037\
        );

    \I__19693\ : Span4Mux_h
    port map (
            O => \N__79096\,
            I => \N__79034\
        );

    \I__19692\ : LocalMux
    port map (
            O => \N__79093\,
            I => \N__79029\
        );

    \I__19691\ : LocalMux
    port map (
            O => \N__79088\,
            I => \N__79029\
        );

    \I__19690\ : InMux
    port map (
            O => \N__79085\,
            I => \N__79022\
        );

    \I__19689\ : InMux
    port map (
            O => \N__79084\,
            I => \N__79022\
        );

    \I__19688\ : InMux
    port map (
            O => \N__79083\,
            I => \N__79022\
        );

    \I__19687\ : LocalMux
    port map (
            O => \N__79078\,
            I => \N__79019\
        );

    \I__19686\ : Span4Mux_v
    port map (
            O => \N__79075\,
            I => \N__79016\
        );

    \I__19685\ : Span4Mux_h
    port map (
            O => \N__79072\,
            I => \N__79009\
        );

    \I__19684\ : Span4Mux_v
    port map (
            O => \N__79069\,
            I => \N__79009\
        );

    \I__19683\ : LocalMux
    port map (
            O => \N__79066\,
            I => \N__79009\
        );

    \I__19682\ : Span4Mux_v
    port map (
            O => \N__79063\,
            I => \N__79006\
        );

    \I__19681\ : Span4Mux_v
    port map (
            O => \N__79060\,
            I => \N__79001\
        );

    \I__19680\ : Span4Mux_h
    port map (
            O => \N__79055\,
            I => \N__79001\
        );

    \I__19679\ : LocalMux
    port map (
            O => \N__79052\,
            I => \N__78998\
        );

    \I__19678\ : CascadeMux
    port map (
            O => \N__79051\,
            I => \N__78995\
        );

    \I__19677\ : LocalMux
    port map (
            O => \N__79046\,
            I => \N__78985\
        );

    \I__19676\ : LocalMux
    port map (
            O => \N__79043\,
            I => \N__78985\
        );

    \I__19675\ : LocalMux
    port map (
            O => \N__79040\,
            I => \N__78985\
        );

    \I__19674\ : Sp12to4
    port map (
            O => \N__79037\,
            I => \N__78985\
        );

    \I__19673\ : Span4Mux_v
    port map (
            O => \N__79034\,
            I => \N__78980\
        );

    \I__19672\ : Span4Mux_v
    port map (
            O => \N__79029\,
            I => \N__78980\
        );

    \I__19671\ : LocalMux
    port map (
            O => \N__79022\,
            I => \N__78975\
        );

    \I__19670\ : Span4Mux_h
    port map (
            O => \N__79019\,
            I => \N__78970\
        );

    \I__19669\ : Span4Mux_v
    port map (
            O => \N__79016\,
            I => \N__78970\
        );

    \I__19668\ : Span4Mux_v
    port map (
            O => \N__79009\,
            I => \N__78963\
        );

    \I__19667\ : Span4Mux_v
    port map (
            O => \N__79006\,
            I => \N__78963\
        );

    \I__19666\ : Span4Mux_v
    port map (
            O => \N__79001\,
            I => \N__78963\
        );

    \I__19665\ : Span4Mux_h
    port map (
            O => \N__78998\,
            I => \N__78960\
        );

    \I__19664\ : InMux
    port map (
            O => \N__78995\,
            I => \N__78955\
        );

    \I__19663\ : InMux
    port map (
            O => \N__78994\,
            I => \N__78955\
        );

    \I__19662\ : Span12Mux_h
    port map (
            O => \N__78985\,
            I => \N__78952\
        );

    \I__19661\ : Sp12to4
    port map (
            O => \N__78980\,
            I => \N__78949\
        );

    \I__19660\ : InMux
    port map (
            O => \N__78979\,
            I => \N__78946\
        );

    \I__19659\ : InMux
    port map (
            O => \N__78978\,
            I => \N__78943\
        );

    \I__19658\ : Span4Mux_h
    port map (
            O => \N__78975\,
            I => \N__78938\
        );

    \I__19657\ : Span4Mux_h
    port map (
            O => \N__78970\,
            I => \N__78938\
        );

    \I__19656\ : Span4Mux_h
    port map (
            O => \N__78963\,
            I => \N__78933\
        );

    \I__19655\ : Span4Mux_v
    port map (
            O => \N__78960\,
            I => \N__78933\
        );

    \I__19654\ : LocalMux
    port map (
            O => \N__78955\,
            I => \N__78926\
        );

    \I__19653\ : Span12Mux_v
    port map (
            O => \N__78952\,
            I => \N__78926\
        );

    \I__19652\ : Span12Mux_v
    port map (
            O => \N__78949\,
            I => \N__78926\
        );

    \I__19651\ : LocalMux
    port map (
            O => \N__78946\,
            I => rx_data_2
        );

    \I__19650\ : LocalMux
    port map (
            O => \N__78943\,
            I => rx_data_2
        );

    \I__19649\ : Odrv4
    port map (
            O => \N__78938\,
            I => rx_data_2
        );

    \I__19648\ : Odrv4
    port map (
            O => \N__78933\,
            I => rx_data_2
        );

    \I__19647\ : Odrv12
    port map (
            O => \N__78926\,
            I => rx_data_2
        );

    \I__19646\ : InMux
    port map (
            O => \N__78915\,
            I => \N__78912\
        );

    \I__19645\ : LocalMux
    port map (
            O => \N__78912\,
            I => \N__78908\
        );

    \I__19644\ : InMux
    port map (
            O => \N__78911\,
            I => \N__78905\
        );

    \I__19643\ : Span4Mux_v
    port map (
            O => \N__78908\,
            I => \N__78901\
        );

    \I__19642\ : LocalMux
    port map (
            O => \N__78905\,
            I => \N__78898\
        );

    \I__19641\ : InMux
    port map (
            O => \N__78904\,
            I => \N__78892\
        );

    \I__19640\ : Span4Mux_h
    port map (
            O => \N__78901\,
            I => \N__78887\
        );

    \I__19639\ : Span4Mux_v
    port map (
            O => \N__78898\,
            I => \N__78884\
        );

    \I__19638\ : InMux
    port map (
            O => \N__78897\,
            I => \N__78881\
        );

    \I__19637\ : InMux
    port map (
            O => \N__78896\,
            I => \N__78876\
        );

    \I__19636\ : InMux
    port map (
            O => \N__78895\,
            I => \N__78876\
        );

    \I__19635\ : LocalMux
    port map (
            O => \N__78892\,
            I => \N__78873\
        );

    \I__19634\ : InMux
    port map (
            O => \N__78891\,
            I => \N__78870\
        );

    \I__19633\ : InMux
    port map (
            O => \N__78890\,
            I => \N__78867\
        );

    \I__19632\ : Odrv4
    port map (
            O => \N__78887\,
            I => n22110
        );

    \I__19631\ : Odrv4
    port map (
            O => \N__78884\,
            I => n22110
        );

    \I__19630\ : LocalMux
    port map (
            O => \N__78881\,
            I => n22110
        );

    \I__19629\ : LocalMux
    port map (
            O => \N__78876\,
            I => n22110
        );

    \I__19628\ : Odrv12
    port map (
            O => \N__78873\,
            I => n22110
        );

    \I__19627\ : LocalMux
    port map (
            O => \N__78870\,
            I => n22110
        );

    \I__19626\ : LocalMux
    port map (
            O => \N__78867\,
            I => n22110
        );

    \I__19625\ : InMux
    port map (
            O => \N__78852\,
            I => \N__78849\
        );

    \I__19624\ : LocalMux
    port map (
            O => \N__78849\,
            I => \N__78846\
        );

    \I__19623\ : Span4Mux_h
    port map (
            O => \N__78846\,
            I => \N__78843\
        );

    \I__19622\ : Span4Mux_v
    port map (
            O => \N__78843\,
            I => \N__78838\
        );

    \I__19621\ : InMux
    port map (
            O => \N__78842\,
            I => \N__78833\
        );

    \I__19620\ : InMux
    port map (
            O => \N__78841\,
            I => \N__78833\
        );

    \I__19619\ : Span4Mux_v
    port map (
            O => \N__78838\,
            I => \N__78830\
        );

    \I__19618\ : LocalMux
    port map (
            O => \N__78833\,
            I => data_in_frame_22_2
        );

    \I__19617\ : Odrv4
    port map (
            O => \N__78830\,
            I => data_in_frame_22_2
        );

    \I__19616\ : ClkMux
    port map (
            O => \N__78825\,
            I => \N__78033\
        );

    \I__19615\ : ClkMux
    port map (
            O => \N__78824\,
            I => \N__78033\
        );

    \I__19614\ : ClkMux
    port map (
            O => \N__78823\,
            I => \N__78033\
        );

    \I__19613\ : ClkMux
    port map (
            O => \N__78822\,
            I => \N__78033\
        );

    \I__19612\ : ClkMux
    port map (
            O => \N__78821\,
            I => \N__78033\
        );

    \I__19611\ : ClkMux
    port map (
            O => \N__78820\,
            I => \N__78033\
        );

    \I__19610\ : ClkMux
    port map (
            O => \N__78819\,
            I => \N__78033\
        );

    \I__19609\ : ClkMux
    port map (
            O => \N__78818\,
            I => \N__78033\
        );

    \I__19608\ : ClkMux
    port map (
            O => \N__78817\,
            I => \N__78033\
        );

    \I__19607\ : ClkMux
    port map (
            O => \N__78816\,
            I => \N__78033\
        );

    \I__19606\ : ClkMux
    port map (
            O => \N__78815\,
            I => \N__78033\
        );

    \I__19605\ : ClkMux
    port map (
            O => \N__78814\,
            I => \N__78033\
        );

    \I__19604\ : ClkMux
    port map (
            O => \N__78813\,
            I => \N__78033\
        );

    \I__19603\ : ClkMux
    port map (
            O => \N__78812\,
            I => \N__78033\
        );

    \I__19602\ : ClkMux
    port map (
            O => \N__78811\,
            I => \N__78033\
        );

    \I__19601\ : ClkMux
    port map (
            O => \N__78810\,
            I => \N__78033\
        );

    \I__19600\ : ClkMux
    port map (
            O => \N__78809\,
            I => \N__78033\
        );

    \I__19599\ : ClkMux
    port map (
            O => \N__78808\,
            I => \N__78033\
        );

    \I__19598\ : ClkMux
    port map (
            O => \N__78807\,
            I => \N__78033\
        );

    \I__19597\ : ClkMux
    port map (
            O => \N__78806\,
            I => \N__78033\
        );

    \I__19596\ : ClkMux
    port map (
            O => \N__78805\,
            I => \N__78033\
        );

    \I__19595\ : ClkMux
    port map (
            O => \N__78804\,
            I => \N__78033\
        );

    \I__19594\ : ClkMux
    port map (
            O => \N__78803\,
            I => \N__78033\
        );

    \I__19593\ : ClkMux
    port map (
            O => \N__78802\,
            I => \N__78033\
        );

    \I__19592\ : ClkMux
    port map (
            O => \N__78801\,
            I => \N__78033\
        );

    \I__19591\ : ClkMux
    port map (
            O => \N__78800\,
            I => \N__78033\
        );

    \I__19590\ : ClkMux
    port map (
            O => \N__78799\,
            I => \N__78033\
        );

    \I__19589\ : ClkMux
    port map (
            O => \N__78798\,
            I => \N__78033\
        );

    \I__19588\ : ClkMux
    port map (
            O => \N__78797\,
            I => \N__78033\
        );

    \I__19587\ : ClkMux
    port map (
            O => \N__78796\,
            I => \N__78033\
        );

    \I__19586\ : ClkMux
    port map (
            O => \N__78795\,
            I => \N__78033\
        );

    \I__19585\ : ClkMux
    port map (
            O => \N__78794\,
            I => \N__78033\
        );

    \I__19584\ : ClkMux
    port map (
            O => \N__78793\,
            I => \N__78033\
        );

    \I__19583\ : ClkMux
    port map (
            O => \N__78792\,
            I => \N__78033\
        );

    \I__19582\ : ClkMux
    port map (
            O => \N__78791\,
            I => \N__78033\
        );

    \I__19581\ : ClkMux
    port map (
            O => \N__78790\,
            I => \N__78033\
        );

    \I__19580\ : ClkMux
    port map (
            O => \N__78789\,
            I => \N__78033\
        );

    \I__19579\ : ClkMux
    port map (
            O => \N__78788\,
            I => \N__78033\
        );

    \I__19578\ : ClkMux
    port map (
            O => \N__78787\,
            I => \N__78033\
        );

    \I__19577\ : ClkMux
    port map (
            O => \N__78786\,
            I => \N__78033\
        );

    \I__19576\ : ClkMux
    port map (
            O => \N__78785\,
            I => \N__78033\
        );

    \I__19575\ : ClkMux
    port map (
            O => \N__78784\,
            I => \N__78033\
        );

    \I__19574\ : ClkMux
    port map (
            O => \N__78783\,
            I => \N__78033\
        );

    \I__19573\ : ClkMux
    port map (
            O => \N__78782\,
            I => \N__78033\
        );

    \I__19572\ : ClkMux
    port map (
            O => \N__78781\,
            I => \N__78033\
        );

    \I__19571\ : ClkMux
    port map (
            O => \N__78780\,
            I => \N__78033\
        );

    \I__19570\ : ClkMux
    port map (
            O => \N__78779\,
            I => \N__78033\
        );

    \I__19569\ : ClkMux
    port map (
            O => \N__78778\,
            I => \N__78033\
        );

    \I__19568\ : ClkMux
    port map (
            O => \N__78777\,
            I => \N__78033\
        );

    \I__19567\ : ClkMux
    port map (
            O => \N__78776\,
            I => \N__78033\
        );

    \I__19566\ : ClkMux
    port map (
            O => \N__78775\,
            I => \N__78033\
        );

    \I__19565\ : ClkMux
    port map (
            O => \N__78774\,
            I => \N__78033\
        );

    \I__19564\ : ClkMux
    port map (
            O => \N__78773\,
            I => \N__78033\
        );

    \I__19563\ : ClkMux
    port map (
            O => \N__78772\,
            I => \N__78033\
        );

    \I__19562\ : ClkMux
    port map (
            O => \N__78771\,
            I => \N__78033\
        );

    \I__19561\ : ClkMux
    port map (
            O => \N__78770\,
            I => \N__78033\
        );

    \I__19560\ : ClkMux
    port map (
            O => \N__78769\,
            I => \N__78033\
        );

    \I__19559\ : ClkMux
    port map (
            O => \N__78768\,
            I => \N__78033\
        );

    \I__19558\ : ClkMux
    port map (
            O => \N__78767\,
            I => \N__78033\
        );

    \I__19557\ : ClkMux
    port map (
            O => \N__78766\,
            I => \N__78033\
        );

    \I__19556\ : ClkMux
    port map (
            O => \N__78765\,
            I => \N__78033\
        );

    \I__19555\ : ClkMux
    port map (
            O => \N__78764\,
            I => \N__78033\
        );

    \I__19554\ : ClkMux
    port map (
            O => \N__78763\,
            I => \N__78033\
        );

    \I__19553\ : ClkMux
    port map (
            O => \N__78762\,
            I => \N__78033\
        );

    \I__19552\ : ClkMux
    port map (
            O => \N__78761\,
            I => \N__78033\
        );

    \I__19551\ : ClkMux
    port map (
            O => \N__78760\,
            I => \N__78033\
        );

    \I__19550\ : ClkMux
    port map (
            O => \N__78759\,
            I => \N__78033\
        );

    \I__19549\ : ClkMux
    port map (
            O => \N__78758\,
            I => \N__78033\
        );

    \I__19548\ : ClkMux
    port map (
            O => \N__78757\,
            I => \N__78033\
        );

    \I__19547\ : ClkMux
    port map (
            O => \N__78756\,
            I => \N__78033\
        );

    \I__19546\ : ClkMux
    port map (
            O => \N__78755\,
            I => \N__78033\
        );

    \I__19545\ : ClkMux
    port map (
            O => \N__78754\,
            I => \N__78033\
        );

    \I__19544\ : ClkMux
    port map (
            O => \N__78753\,
            I => \N__78033\
        );

    \I__19543\ : ClkMux
    port map (
            O => \N__78752\,
            I => \N__78033\
        );

    \I__19542\ : ClkMux
    port map (
            O => \N__78751\,
            I => \N__78033\
        );

    \I__19541\ : ClkMux
    port map (
            O => \N__78750\,
            I => \N__78033\
        );

    \I__19540\ : ClkMux
    port map (
            O => \N__78749\,
            I => \N__78033\
        );

    \I__19539\ : ClkMux
    port map (
            O => \N__78748\,
            I => \N__78033\
        );

    \I__19538\ : ClkMux
    port map (
            O => \N__78747\,
            I => \N__78033\
        );

    \I__19537\ : ClkMux
    port map (
            O => \N__78746\,
            I => \N__78033\
        );

    \I__19536\ : ClkMux
    port map (
            O => \N__78745\,
            I => \N__78033\
        );

    \I__19535\ : ClkMux
    port map (
            O => \N__78744\,
            I => \N__78033\
        );

    \I__19534\ : ClkMux
    port map (
            O => \N__78743\,
            I => \N__78033\
        );

    \I__19533\ : ClkMux
    port map (
            O => \N__78742\,
            I => \N__78033\
        );

    \I__19532\ : ClkMux
    port map (
            O => \N__78741\,
            I => \N__78033\
        );

    \I__19531\ : ClkMux
    port map (
            O => \N__78740\,
            I => \N__78033\
        );

    \I__19530\ : ClkMux
    port map (
            O => \N__78739\,
            I => \N__78033\
        );

    \I__19529\ : ClkMux
    port map (
            O => \N__78738\,
            I => \N__78033\
        );

    \I__19528\ : ClkMux
    port map (
            O => \N__78737\,
            I => \N__78033\
        );

    \I__19527\ : ClkMux
    port map (
            O => \N__78736\,
            I => \N__78033\
        );

    \I__19526\ : ClkMux
    port map (
            O => \N__78735\,
            I => \N__78033\
        );

    \I__19525\ : ClkMux
    port map (
            O => \N__78734\,
            I => \N__78033\
        );

    \I__19524\ : ClkMux
    port map (
            O => \N__78733\,
            I => \N__78033\
        );

    \I__19523\ : ClkMux
    port map (
            O => \N__78732\,
            I => \N__78033\
        );

    \I__19522\ : ClkMux
    port map (
            O => \N__78731\,
            I => \N__78033\
        );

    \I__19521\ : ClkMux
    port map (
            O => \N__78730\,
            I => \N__78033\
        );

    \I__19520\ : ClkMux
    port map (
            O => \N__78729\,
            I => \N__78033\
        );

    \I__19519\ : ClkMux
    port map (
            O => \N__78728\,
            I => \N__78033\
        );

    \I__19518\ : ClkMux
    port map (
            O => \N__78727\,
            I => \N__78033\
        );

    \I__19517\ : ClkMux
    port map (
            O => \N__78726\,
            I => \N__78033\
        );

    \I__19516\ : ClkMux
    port map (
            O => \N__78725\,
            I => \N__78033\
        );

    \I__19515\ : ClkMux
    port map (
            O => \N__78724\,
            I => \N__78033\
        );

    \I__19514\ : ClkMux
    port map (
            O => \N__78723\,
            I => \N__78033\
        );

    \I__19513\ : ClkMux
    port map (
            O => \N__78722\,
            I => \N__78033\
        );

    \I__19512\ : ClkMux
    port map (
            O => \N__78721\,
            I => \N__78033\
        );

    \I__19511\ : ClkMux
    port map (
            O => \N__78720\,
            I => \N__78033\
        );

    \I__19510\ : ClkMux
    port map (
            O => \N__78719\,
            I => \N__78033\
        );

    \I__19509\ : ClkMux
    port map (
            O => \N__78718\,
            I => \N__78033\
        );

    \I__19508\ : ClkMux
    port map (
            O => \N__78717\,
            I => \N__78033\
        );

    \I__19507\ : ClkMux
    port map (
            O => \N__78716\,
            I => \N__78033\
        );

    \I__19506\ : ClkMux
    port map (
            O => \N__78715\,
            I => \N__78033\
        );

    \I__19505\ : ClkMux
    port map (
            O => \N__78714\,
            I => \N__78033\
        );

    \I__19504\ : ClkMux
    port map (
            O => \N__78713\,
            I => \N__78033\
        );

    \I__19503\ : ClkMux
    port map (
            O => \N__78712\,
            I => \N__78033\
        );

    \I__19502\ : ClkMux
    port map (
            O => \N__78711\,
            I => \N__78033\
        );

    \I__19501\ : ClkMux
    port map (
            O => \N__78710\,
            I => \N__78033\
        );

    \I__19500\ : ClkMux
    port map (
            O => \N__78709\,
            I => \N__78033\
        );

    \I__19499\ : ClkMux
    port map (
            O => \N__78708\,
            I => \N__78033\
        );

    \I__19498\ : ClkMux
    port map (
            O => \N__78707\,
            I => \N__78033\
        );

    \I__19497\ : ClkMux
    port map (
            O => \N__78706\,
            I => \N__78033\
        );

    \I__19496\ : ClkMux
    port map (
            O => \N__78705\,
            I => \N__78033\
        );

    \I__19495\ : ClkMux
    port map (
            O => \N__78704\,
            I => \N__78033\
        );

    \I__19494\ : ClkMux
    port map (
            O => \N__78703\,
            I => \N__78033\
        );

    \I__19493\ : ClkMux
    port map (
            O => \N__78702\,
            I => \N__78033\
        );

    \I__19492\ : ClkMux
    port map (
            O => \N__78701\,
            I => \N__78033\
        );

    \I__19491\ : ClkMux
    port map (
            O => \N__78700\,
            I => \N__78033\
        );

    \I__19490\ : ClkMux
    port map (
            O => \N__78699\,
            I => \N__78033\
        );

    \I__19489\ : ClkMux
    port map (
            O => \N__78698\,
            I => \N__78033\
        );

    \I__19488\ : ClkMux
    port map (
            O => \N__78697\,
            I => \N__78033\
        );

    \I__19487\ : ClkMux
    port map (
            O => \N__78696\,
            I => \N__78033\
        );

    \I__19486\ : ClkMux
    port map (
            O => \N__78695\,
            I => \N__78033\
        );

    \I__19485\ : ClkMux
    port map (
            O => \N__78694\,
            I => \N__78033\
        );

    \I__19484\ : ClkMux
    port map (
            O => \N__78693\,
            I => \N__78033\
        );

    \I__19483\ : ClkMux
    port map (
            O => \N__78692\,
            I => \N__78033\
        );

    \I__19482\ : ClkMux
    port map (
            O => \N__78691\,
            I => \N__78033\
        );

    \I__19481\ : ClkMux
    port map (
            O => \N__78690\,
            I => \N__78033\
        );

    \I__19480\ : ClkMux
    port map (
            O => \N__78689\,
            I => \N__78033\
        );

    \I__19479\ : ClkMux
    port map (
            O => \N__78688\,
            I => \N__78033\
        );

    \I__19478\ : ClkMux
    port map (
            O => \N__78687\,
            I => \N__78033\
        );

    \I__19477\ : ClkMux
    port map (
            O => \N__78686\,
            I => \N__78033\
        );

    \I__19476\ : ClkMux
    port map (
            O => \N__78685\,
            I => \N__78033\
        );

    \I__19475\ : ClkMux
    port map (
            O => \N__78684\,
            I => \N__78033\
        );

    \I__19474\ : ClkMux
    port map (
            O => \N__78683\,
            I => \N__78033\
        );

    \I__19473\ : ClkMux
    port map (
            O => \N__78682\,
            I => \N__78033\
        );

    \I__19472\ : ClkMux
    port map (
            O => \N__78681\,
            I => \N__78033\
        );

    \I__19471\ : ClkMux
    port map (
            O => \N__78680\,
            I => \N__78033\
        );

    \I__19470\ : ClkMux
    port map (
            O => \N__78679\,
            I => \N__78033\
        );

    \I__19469\ : ClkMux
    port map (
            O => \N__78678\,
            I => \N__78033\
        );

    \I__19468\ : ClkMux
    port map (
            O => \N__78677\,
            I => \N__78033\
        );

    \I__19467\ : ClkMux
    port map (
            O => \N__78676\,
            I => \N__78033\
        );

    \I__19466\ : ClkMux
    port map (
            O => \N__78675\,
            I => \N__78033\
        );

    \I__19465\ : ClkMux
    port map (
            O => \N__78674\,
            I => \N__78033\
        );

    \I__19464\ : ClkMux
    port map (
            O => \N__78673\,
            I => \N__78033\
        );

    \I__19463\ : ClkMux
    port map (
            O => \N__78672\,
            I => \N__78033\
        );

    \I__19462\ : ClkMux
    port map (
            O => \N__78671\,
            I => \N__78033\
        );

    \I__19461\ : ClkMux
    port map (
            O => \N__78670\,
            I => \N__78033\
        );

    \I__19460\ : ClkMux
    port map (
            O => \N__78669\,
            I => \N__78033\
        );

    \I__19459\ : ClkMux
    port map (
            O => \N__78668\,
            I => \N__78033\
        );

    \I__19458\ : ClkMux
    port map (
            O => \N__78667\,
            I => \N__78033\
        );

    \I__19457\ : ClkMux
    port map (
            O => \N__78666\,
            I => \N__78033\
        );

    \I__19456\ : ClkMux
    port map (
            O => \N__78665\,
            I => \N__78033\
        );

    \I__19455\ : ClkMux
    port map (
            O => \N__78664\,
            I => \N__78033\
        );

    \I__19454\ : ClkMux
    port map (
            O => \N__78663\,
            I => \N__78033\
        );

    \I__19453\ : ClkMux
    port map (
            O => \N__78662\,
            I => \N__78033\
        );

    \I__19452\ : ClkMux
    port map (
            O => \N__78661\,
            I => \N__78033\
        );

    \I__19451\ : ClkMux
    port map (
            O => \N__78660\,
            I => \N__78033\
        );

    \I__19450\ : ClkMux
    port map (
            O => \N__78659\,
            I => \N__78033\
        );

    \I__19449\ : ClkMux
    port map (
            O => \N__78658\,
            I => \N__78033\
        );

    \I__19448\ : ClkMux
    port map (
            O => \N__78657\,
            I => \N__78033\
        );

    \I__19447\ : ClkMux
    port map (
            O => \N__78656\,
            I => \N__78033\
        );

    \I__19446\ : ClkMux
    port map (
            O => \N__78655\,
            I => \N__78033\
        );

    \I__19445\ : ClkMux
    port map (
            O => \N__78654\,
            I => \N__78033\
        );

    \I__19444\ : ClkMux
    port map (
            O => \N__78653\,
            I => \N__78033\
        );

    \I__19443\ : ClkMux
    port map (
            O => \N__78652\,
            I => \N__78033\
        );

    \I__19442\ : ClkMux
    port map (
            O => \N__78651\,
            I => \N__78033\
        );

    \I__19441\ : ClkMux
    port map (
            O => \N__78650\,
            I => \N__78033\
        );

    \I__19440\ : ClkMux
    port map (
            O => \N__78649\,
            I => \N__78033\
        );

    \I__19439\ : ClkMux
    port map (
            O => \N__78648\,
            I => \N__78033\
        );

    \I__19438\ : ClkMux
    port map (
            O => \N__78647\,
            I => \N__78033\
        );

    \I__19437\ : ClkMux
    port map (
            O => \N__78646\,
            I => \N__78033\
        );

    \I__19436\ : ClkMux
    port map (
            O => \N__78645\,
            I => \N__78033\
        );

    \I__19435\ : ClkMux
    port map (
            O => \N__78644\,
            I => \N__78033\
        );

    \I__19434\ : ClkMux
    port map (
            O => \N__78643\,
            I => \N__78033\
        );

    \I__19433\ : ClkMux
    port map (
            O => \N__78642\,
            I => \N__78033\
        );

    \I__19432\ : ClkMux
    port map (
            O => \N__78641\,
            I => \N__78033\
        );

    \I__19431\ : ClkMux
    port map (
            O => \N__78640\,
            I => \N__78033\
        );

    \I__19430\ : ClkMux
    port map (
            O => \N__78639\,
            I => \N__78033\
        );

    \I__19429\ : ClkMux
    port map (
            O => \N__78638\,
            I => \N__78033\
        );

    \I__19428\ : ClkMux
    port map (
            O => \N__78637\,
            I => \N__78033\
        );

    \I__19427\ : ClkMux
    port map (
            O => \N__78636\,
            I => \N__78033\
        );

    \I__19426\ : ClkMux
    port map (
            O => \N__78635\,
            I => \N__78033\
        );

    \I__19425\ : ClkMux
    port map (
            O => \N__78634\,
            I => \N__78033\
        );

    \I__19424\ : ClkMux
    port map (
            O => \N__78633\,
            I => \N__78033\
        );

    \I__19423\ : ClkMux
    port map (
            O => \N__78632\,
            I => \N__78033\
        );

    \I__19422\ : ClkMux
    port map (
            O => \N__78631\,
            I => \N__78033\
        );

    \I__19421\ : ClkMux
    port map (
            O => \N__78630\,
            I => \N__78033\
        );

    \I__19420\ : ClkMux
    port map (
            O => \N__78629\,
            I => \N__78033\
        );

    \I__19419\ : ClkMux
    port map (
            O => \N__78628\,
            I => \N__78033\
        );

    \I__19418\ : ClkMux
    port map (
            O => \N__78627\,
            I => \N__78033\
        );

    \I__19417\ : ClkMux
    port map (
            O => \N__78626\,
            I => \N__78033\
        );

    \I__19416\ : ClkMux
    port map (
            O => \N__78625\,
            I => \N__78033\
        );

    \I__19415\ : ClkMux
    port map (
            O => \N__78624\,
            I => \N__78033\
        );

    \I__19414\ : ClkMux
    port map (
            O => \N__78623\,
            I => \N__78033\
        );

    \I__19413\ : ClkMux
    port map (
            O => \N__78622\,
            I => \N__78033\
        );

    \I__19412\ : ClkMux
    port map (
            O => \N__78621\,
            I => \N__78033\
        );

    \I__19411\ : ClkMux
    port map (
            O => \N__78620\,
            I => \N__78033\
        );

    \I__19410\ : ClkMux
    port map (
            O => \N__78619\,
            I => \N__78033\
        );

    \I__19409\ : ClkMux
    port map (
            O => \N__78618\,
            I => \N__78033\
        );

    \I__19408\ : ClkMux
    port map (
            O => \N__78617\,
            I => \N__78033\
        );

    \I__19407\ : ClkMux
    port map (
            O => \N__78616\,
            I => \N__78033\
        );

    \I__19406\ : ClkMux
    port map (
            O => \N__78615\,
            I => \N__78033\
        );

    \I__19405\ : ClkMux
    port map (
            O => \N__78614\,
            I => \N__78033\
        );

    \I__19404\ : ClkMux
    port map (
            O => \N__78613\,
            I => \N__78033\
        );

    \I__19403\ : ClkMux
    port map (
            O => \N__78612\,
            I => \N__78033\
        );

    \I__19402\ : ClkMux
    port map (
            O => \N__78611\,
            I => \N__78033\
        );

    \I__19401\ : ClkMux
    port map (
            O => \N__78610\,
            I => \N__78033\
        );

    \I__19400\ : ClkMux
    port map (
            O => \N__78609\,
            I => \N__78033\
        );

    \I__19399\ : ClkMux
    port map (
            O => \N__78608\,
            I => \N__78033\
        );

    \I__19398\ : ClkMux
    port map (
            O => \N__78607\,
            I => \N__78033\
        );

    \I__19397\ : ClkMux
    port map (
            O => \N__78606\,
            I => \N__78033\
        );

    \I__19396\ : ClkMux
    port map (
            O => \N__78605\,
            I => \N__78033\
        );

    \I__19395\ : ClkMux
    port map (
            O => \N__78604\,
            I => \N__78033\
        );

    \I__19394\ : ClkMux
    port map (
            O => \N__78603\,
            I => \N__78033\
        );

    \I__19393\ : ClkMux
    port map (
            O => \N__78602\,
            I => \N__78033\
        );

    \I__19392\ : ClkMux
    port map (
            O => \N__78601\,
            I => \N__78033\
        );

    \I__19391\ : ClkMux
    port map (
            O => \N__78600\,
            I => \N__78033\
        );

    \I__19390\ : ClkMux
    port map (
            O => \N__78599\,
            I => \N__78033\
        );

    \I__19389\ : ClkMux
    port map (
            O => \N__78598\,
            I => \N__78033\
        );

    \I__19388\ : ClkMux
    port map (
            O => \N__78597\,
            I => \N__78033\
        );

    \I__19387\ : ClkMux
    port map (
            O => \N__78596\,
            I => \N__78033\
        );

    \I__19386\ : ClkMux
    port map (
            O => \N__78595\,
            I => \N__78033\
        );

    \I__19385\ : ClkMux
    port map (
            O => \N__78594\,
            I => \N__78033\
        );

    \I__19384\ : ClkMux
    port map (
            O => \N__78593\,
            I => \N__78033\
        );

    \I__19383\ : ClkMux
    port map (
            O => \N__78592\,
            I => \N__78033\
        );

    \I__19382\ : ClkMux
    port map (
            O => \N__78591\,
            I => \N__78033\
        );

    \I__19381\ : ClkMux
    port map (
            O => \N__78590\,
            I => \N__78033\
        );

    \I__19380\ : ClkMux
    port map (
            O => \N__78589\,
            I => \N__78033\
        );

    \I__19379\ : ClkMux
    port map (
            O => \N__78588\,
            I => \N__78033\
        );

    \I__19378\ : ClkMux
    port map (
            O => \N__78587\,
            I => \N__78033\
        );

    \I__19377\ : ClkMux
    port map (
            O => \N__78586\,
            I => \N__78033\
        );

    \I__19376\ : ClkMux
    port map (
            O => \N__78585\,
            I => \N__78033\
        );

    \I__19375\ : ClkMux
    port map (
            O => \N__78584\,
            I => \N__78033\
        );

    \I__19374\ : ClkMux
    port map (
            O => \N__78583\,
            I => \N__78033\
        );

    \I__19373\ : ClkMux
    port map (
            O => \N__78582\,
            I => \N__78033\
        );

    \I__19372\ : ClkMux
    port map (
            O => \N__78581\,
            I => \N__78033\
        );

    \I__19371\ : ClkMux
    port map (
            O => \N__78580\,
            I => \N__78033\
        );

    \I__19370\ : ClkMux
    port map (
            O => \N__78579\,
            I => \N__78033\
        );

    \I__19369\ : ClkMux
    port map (
            O => \N__78578\,
            I => \N__78033\
        );

    \I__19368\ : ClkMux
    port map (
            O => \N__78577\,
            I => \N__78033\
        );

    \I__19367\ : ClkMux
    port map (
            O => \N__78576\,
            I => \N__78033\
        );

    \I__19366\ : ClkMux
    port map (
            O => \N__78575\,
            I => \N__78033\
        );

    \I__19365\ : ClkMux
    port map (
            O => \N__78574\,
            I => \N__78033\
        );

    \I__19364\ : ClkMux
    port map (
            O => \N__78573\,
            I => \N__78033\
        );

    \I__19363\ : ClkMux
    port map (
            O => \N__78572\,
            I => \N__78033\
        );

    \I__19362\ : ClkMux
    port map (
            O => \N__78571\,
            I => \N__78033\
        );

    \I__19361\ : ClkMux
    port map (
            O => \N__78570\,
            I => \N__78033\
        );

    \I__19360\ : ClkMux
    port map (
            O => \N__78569\,
            I => \N__78033\
        );

    \I__19359\ : ClkMux
    port map (
            O => \N__78568\,
            I => \N__78033\
        );

    \I__19358\ : ClkMux
    port map (
            O => \N__78567\,
            I => \N__78033\
        );

    \I__19357\ : ClkMux
    port map (
            O => \N__78566\,
            I => \N__78033\
        );

    \I__19356\ : ClkMux
    port map (
            O => \N__78565\,
            I => \N__78033\
        );

    \I__19355\ : ClkMux
    port map (
            O => \N__78564\,
            I => \N__78033\
        );

    \I__19354\ : ClkMux
    port map (
            O => \N__78563\,
            I => \N__78033\
        );

    \I__19353\ : ClkMux
    port map (
            O => \N__78562\,
            I => \N__78033\
        );

    \I__19352\ : GlobalMux
    port map (
            O => \N__78033\,
            I => \N__78030\
        );

    \I__19351\ : gio2CtrlBuf
    port map (
            O => \N__78030\,
            I => \CLK_c\
        );

    \I__19350\ : InMux
    port map (
            O => \N__78027\,
            I => \N__78021\
        );

    \I__19349\ : InMux
    port map (
            O => \N__78026\,
            I => \N__78014\
        );

    \I__19348\ : InMux
    port map (
            O => \N__78025\,
            I => \N__78009\
        );

    \I__19347\ : InMux
    port map (
            O => \N__78024\,
            I => \N__78009\
        );

    \I__19346\ : LocalMux
    port map (
            O => \N__78021\,
            I => \N__78006\
        );

    \I__19345\ : InMux
    port map (
            O => \N__78020\,
            I => \N__78003\
        );

    \I__19344\ : InMux
    port map (
            O => \N__78019\,
            I => \N__77998\
        );

    \I__19343\ : InMux
    port map (
            O => \N__78018\,
            I => \N__77998\
        );

    \I__19342\ : CascadeMux
    port map (
            O => \N__78017\,
            I => \N__77995\
        );

    \I__19341\ : LocalMux
    port map (
            O => \N__78014\,
            I => \N__77992\
        );

    \I__19340\ : LocalMux
    port map (
            O => \N__78009\,
            I => \N__77987\
        );

    \I__19339\ : Span4Mux_v
    port map (
            O => \N__78006\,
            I => \N__77987\
        );

    \I__19338\ : LocalMux
    port map (
            O => \N__78003\,
            I => \N__77982\
        );

    \I__19337\ : LocalMux
    port map (
            O => \N__77998\,
            I => \N__77982\
        );

    \I__19336\ : InMux
    port map (
            O => \N__77995\,
            I => \N__77979\
        );

    \I__19335\ : Span4Mux_v
    port map (
            O => \N__77992\,
            I => \N__77976\
        );

    \I__19334\ : Span4Mux_h
    port map (
            O => \N__77987\,
            I => \N__77971\
        );

    \I__19333\ : Span4Mux_v
    port map (
            O => \N__77982\,
            I => \N__77971\
        );

    \I__19332\ : LocalMux
    port map (
            O => \N__77979\,
            I => \N__77966\
        );

    \I__19331\ : Span4Mux_h
    port map (
            O => \N__77976\,
            I => \N__77966\
        );

    \I__19330\ : Span4Mux_h
    port map (
            O => \N__77971\,
            I => \N__77963\
        );

    \I__19329\ : Odrv4
    port map (
            O => \N__77966\,
            I => \c0.data_in_frame_24_0\
        );

    \I__19328\ : Odrv4
    port map (
            O => \N__77963\,
            I => \c0.data_in_frame_24_0\
        );

    \I__19327\ : InMux
    port map (
            O => \N__77958\,
            I => \N__77951\
        );

    \I__19326\ : InMux
    port map (
            O => \N__77957\,
            I => \N__77948\
        );

    \I__19325\ : InMux
    port map (
            O => \N__77956\,
            I => \N__77945\
        );

    \I__19324\ : InMux
    port map (
            O => \N__77955\,
            I => \N__77942\
        );

    \I__19323\ : InMux
    port map (
            O => \N__77954\,
            I => \N__77939\
        );

    \I__19322\ : LocalMux
    port map (
            O => \N__77951\,
            I => \N__77933\
        );

    \I__19321\ : LocalMux
    port map (
            O => \N__77948\,
            I => \N__77933\
        );

    \I__19320\ : LocalMux
    port map (
            O => \N__77945\,
            I => \N__77928\
        );

    \I__19319\ : LocalMux
    port map (
            O => \N__77942\,
            I => \N__77928\
        );

    \I__19318\ : LocalMux
    port map (
            O => \N__77939\,
            I => \N__77925\
        );

    \I__19317\ : InMux
    port map (
            O => \N__77938\,
            I => \N__77922\
        );

    \I__19316\ : Span4Mux_v
    port map (
            O => \N__77933\,
            I => \N__77919\
        );

    \I__19315\ : Span4Mux_h
    port map (
            O => \N__77928\,
            I => \N__77914\
        );

    \I__19314\ : Span4Mux_v
    port map (
            O => \N__77925\,
            I => \N__77914\
        );

    \I__19313\ : LocalMux
    port map (
            O => \N__77922\,
            I => \N__77911\
        );

    \I__19312\ : Span4Mux_v
    port map (
            O => \N__77919\,
            I => \N__77906\
        );

    \I__19311\ : Span4Mux_v
    port map (
            O => \N__77914\,
            I => \N__77906\
        );

    \I__19310\ : Span12Mux_h
    port map (
            O => \N__77911\,
            I => \N__77903\
        );

    \I__19309\ : Odrv4
    port map (
            O => \N__77906\,
            I => \c0.n29_adj_4362\
        );

    \I__19308\ : Odrv12
    port map (
            O => \N__77903\,
            I => \c0.n29_adj_4362\
        );

    \I__19307\ : InMux
    port map (
            O => \N__77898\,
            I => \N__77895\
        );

    \I__19306\ : LocalMux
    port map (
            O => \N__77895\,
            I => \N__77892\
        );

    \I__19305\ : Span4Mux_v
    port map (
            O => \N__77892\,
            I => \N__77889\
        );

    \I__19304\ : Span4Mux_h
    port map (
            O => \N__77889\,
            I => \N__77886\
        );

    \I__19303\ : Odrv4
    port map (
            O => \N__77886\,
            I => \c0.n24_adj_4531\
        );

    \I__19302\ : InMux
    port map (
            O => \N__77883\,
            I => \N__77880\
        );

    \I__19301\ : LocalMux
    port map (
            O => \N__77880\,
            I => \N__77876\
        );

    \I__19300\ : InMux
    port map (
            O => \N__77879\,
            I => \N__77873\
        );

    \I__19299\ : Span4Mux_h
    port map (
            O => \N__77876\,
            I => \N__77869\
        );

    \I__19298\ : LocalMux
    port map (
            O => \N__77873\,
            I => \N__77866\
        );

    \I__19297\ : InMux
    port map (
            O => \N__77872\,
            I => \N__77863\
        );

    \I__19296\ : Span4Mux_h
    port map (
            O => \N__77869\,
            I => \N__77858\
        );

    \I__19295\ : Span4Mux_v
    port map (
            O => \N__77866\,
            I => \N__77858\
        );

    \I__19294\ : LocalMux
    port map (
            O => \N__77863\,
            I => \N__77853\
        );

    \I__19293\ : Span4Mux_v
    port map (
            O => \N__77858\,
            I => \N__77850\
        );

    \I__19292\ : InMux
    port map (
            O => \N__77857\,
            I => \N__77847\
        );

    \I__19291\ : InMux
    port map (
            O => \N__77856\,
            I => \N__77841\
        );

    \I__19290\ : Span12Mux_v
    port map (
            O => \N__77853\,
            I => \N__77838\
        );

    \I__19289\ : Span4Mux_h
    port map (
            O => \N__77850\,
            I => \N__77833\
        );

    \I__19288\ : LocalMux
    port map (
            O => \N__77847\,
            I => \N__77833\
        );

    \I__19287\ : InMux
    port map (
            O => \N__77846\,
            I => \N__77826\
        );

    \I__19286\ : InMux
    port map (
            O => \N__77845\,
            I => \N__77826\
        );

    \I__19285\ : InMux
    port map (
            O => \N__77844\,
            I => \N__77826\
        );

    \I__19284\ : LocalMux
    port map (
            O => \N__77841\,
            I => data_in_frame_6_3
        );

    \I__19283\ : Odrv12
    port map (
            O => \N__77838\,
            I => data_in_frame_6_3
        );

    \I__19282\ : Odrv4
    port map (
            O => \N__77833\,
            I => data_in_frame_6_3
        );

    \I__19281\ : LocalMux
    port map (
            O => \N__77826\,
            I => data_in_frame_6_3
        );

    \I__19280\ : InMux
    port map (
            O => \N__77817\,
            I => \N__77813\
        );

    \I__19279\ : InMux
    port map (
            O => \N__77816\,
            I => \N__77807\
        );

    \I__19278\ : LocalMux
    port map (
            O => \N__77813\,
            I => \N__77804\
        );

    \I__19277\ : InMux
    port map (
            O => \N__77812\,
            I => \N__77799\
        );

    \I__19276\ : InMux
    port map (
            O => \N__77811\,
            I => \N__77799\
        );

    \I__19275\ : InMux
    port map (
            O => \N__77810\,
            I => \N__77796\
        );

    \I__19274\ : LocalMux
    port map (
            O => \N__77807\,
            I => \N__77793\
        );

    \I__19273\ : Span4Mux_v
    port map (
            O => \N__77804\,
            I => \N__77789\
        );

    \I__19272\ : LocalMux
    port map (
            O => \N__77799\,
            I => \N__77784\
        );

    \I__19271\ : LocalMux
    port map (
            O => \N__77796\,
            I => \N__77784\
        );

    \I__19270\ : Span4Mux_v
    port map (
            O => \N__77793\,
            I => \N__77781\
        );

    \I__19269\ : InMux
    port map (
            O => \N__77792\,
            I => \N__77778\
        );

    \I__19268\ : Span4Mux_h
    port map (
            O => \N__77789\,
            I => \N__77771\
        );

    \I__19267\ : Span4Mux_v
    port map (
            O => \N__77784\,
            I => \N__77771\
        );

    \I__19266\ : Span4Mux_v
    port map (
            O => \N__77781\,
            I => \N__77766\
        );

    \I__19265\ : LocalMux
    port map (
            O => \N__77778\,
            I => \N__77766\
        );

    \I__19264\ : InMux
    port map (
            O => \N__77777\,
            I => \N__77761\
        );

    \I__19263\ : InMux
    port map (
            O => \N__77776\,
            I => \N__77761\
        );

    \I__19262\ : Odrv4
    port map (
            O => \N__77771\,
            I => \c0.n23267\
        );

    \I__19261\ : Odrv4
    port map (
            O => \N__77766\,
            I => \c0.n23267\
        );

    \I__19260\ : LocalMux
    port map (
            O => \N__77761\,
            I => \c0.n23267\
        );

    \I__19259\ : CascadeMux
    port map (
            O => \N__77754\,
            I => \c0.n18_cascade_\
        );

    \I__19258\ : InMux
    port map (
            O => \N__77751\,
            I => \N__77748\
        );

    \I__19257\ : LocalMux
    port map (
            O => \N__77748\,
            I => \N__77745\
        );

    \I__19256\ : Span4Mux_h
    port map (
            O => \N__77745\,
            I => \N__77742\
        );

    \I__19255\ : Odrv4
    port map (
            O => \N__77742\,
            I => \c0.n16_adj_4666\
        );

    \I__19254\ : InMux
    port map (
            O => \N__77739\,
            I => \N__77736\
        );

    \I__19253\ : LocalMux
    port map (
            O => \N__77736\,
            I => \c0.n28_adj_4667\
        );

    \I__19252\ : CascadeMux
    port map (
            O => \N__77733\,
            I => \c0.n24_adj_4653_cascade_\
        );

    \I__19251\ : InMux
    port map (
            O => \N__77730\,
            I => \N__77727\
        );

    \I__19250\ : LocalMux
    port map (
            O => \N__77727\,
            I => \N__77723\
        );

    \I__19249\ : InMux
    port map (
            O => \N__77726\,
            I => \N__77720\
        );

    \I__19248\ : Span4Mux_v
    port map (
            O => \N__77723\,
            I => \N__77715\
        );

    \I__19247\ : LocalMux
    port map (
            O => \N__77720\,
            I => \N__77715\
        );

    \I__19246\ : Span4Mux_h
    port map (
            O => \N__77715\,
            I => \N__77712\
        );

    \I__19245\ : Odrv4
    port map (
            O => \N__77712\,
            I => \c0.n22369\
        );

    \I__19244\ : InMux
    port map (
            O => \N__77709\,
            I => \N__77706\
        );

    \I__19243\ : LocalMux
    port map (
            O => \N__77706\,
            I => \N__77702\
        );

    \I__19242\ : CascadeMux
    port map (
            O => \N__77705\,
            I => \N__77699\
        );

    \I__19241\ : Span4Mux_h
    port map (
            O => \N__77702\,
            I => \N__77696\
        );

    \I__19240\ : InMux
    port map (
            O => \N__77699\,
            I => \N__77693\
        );

    \I__19239\ : Odrv4
    port map (
            O => \N__77696\,
            I => \c0.n6_adj_4587\
        );

    \I__19238\ : LocalMux
    port map (
            O => \N__77693\,
            I => \c0.n6_adj_4587\
        );

    \I__19237\ : InMux
    port map (
            O => \N__77688\,
            I => \N__77684\
        );

    \I__19236\ : InMux
    port map (
            O => \N__77687\,
            I => \N__77681\
        );

    \I__19235\ : LocalMux
    port map (
            O => \N__77684\,
            I => \N__77678\
        );

    \I__19234\ : LocalMux
    port map (
            O => \N__77681\,
            I => \N__77675\
        );

    \I__19233\ : Span4Mux_h
    port map (
            O => \N__77678\,
            I => \N__77668\
        );

    \I__19232\ : Span4Mux_h
    port map (
            O => \N__77675\,
            I => \N__77668\
        );

    \I__19231\ : InMux
    port map (
            O => \N__77674\,
            I => \N__77663\
        );

    \I__19230\ : InMux
    port map (
            O => \N__77673\,
            I => \N__77663\
        );

    \I__19229\ : Span4Mux_h
    port map (
            O => \N__77668\,
            I => \N__77658\
        );

    \I__19228\ : LocalMux
    port map (
            O => \N__77663\,
            I => \N__77658\
        );

    \I__19227\ : Odrv4
    port map (
            O => \N__77658\,
            I => \c0.n22586\
        );

    \I__19226\ : CascadeMux
    port map (
            O => \N__77655\,
            I => \N__77651\
        );

    \I__19225\ : InMux
    port map (
            O => \N__77654\,
            I => \N__77646\
        );

    \I__19224\ : InMux
    port map (
            O => \N__77651\,
            I => \N__77643\
        );

    \I__19223\ : InMux
    port map (
            O => \N__77650\,
            I => \N__77640\
        );

    \I__19222\ : CascadeMux
    port map (
            O => \N__77649\,
            I => \N__77635\
        );

    \I__19221\ : LocalMux
    port map (
            O => \N__77646\,
            I => \N__77632\
        );

    \I__19220\ : LocalMux
    port map (
            O => \N__77643\,
            I => \N__77629\
        );

    \I__19219\ : LocalMux
    port map (
            O => \N__77640\,
            I => \N__77626\
        );

    \I__19218\ : InMux
    port map (
            O => \N__77639\,
            I => \N__77623\
        );

    \I__19217\ : InMux
    port map (
            O => \N__77638\,
            I => \N__77620\
        );

    \I__19216\ : InMux
    port map (
            O => \N__77635\,
            I => \N__77617\
        );

    \I__19215\ : Span4Mux_v
    port map (
            O => \N__77632\,
            I => \N__77614\
        );

    \I__19214\ : Span4Mux_v
    port map (
            O => \N__77629\,
            I => \N__77611\
        );

    \I__19213\ : Span4Mux_v
    port map (
            O => \N__77626\,
            I => \N__77608\
        );

    \I__19212\ : LocalMux
    port map (
            O => \N__77623\,
            I => \N__77605\
        );

    \I__19211\ : LocalMux
    port map (
            O => \N__77620\,
            I => \N__77602\
        );

    \I__19210\ : LocalMux
    port map (
            O => \N__77617\,
            I => \N__77593\
        );

    \I__19209\ : Span4Mux_h
    port map (
            O => \N__77614\,
            I => \N__77593\
        );

    \I__19208\ : Span4Mux_v
    port map (
            O => \N__77611\,
            I => \N__77593\
        );

    \I__19207\ : Span4Mux_v
    port map (
            O => \N__77608\,
            I => \N__77593\
        );

    \I__19206\ : Span4Mux_v
    port map (
            O => \N__77605\,
            I => \N__77590\
        );

    \I__19205\ : Odrv12
    port map (
            O => \N__77602\,
            I => \c0.data_in_frame_19_6\
        );

    \I__19204\ : Odrv4
    port map (
            O => \N__77593\,
            I => \c0.data_in_frame_19_6\
        );

    \I__19203\ : Odrv4
    port map (
            O => \N__77590\,
            I => \c0.data_in_frame_19_6\
        );

    \I__19202\ : InMux
    port map (
            O => \N__77583\,
            I => \N__77580\
        );

    \I__19201\ : LocalMux
    port map (
            O => \N__77580\,
            I => \N__77575\
        );

    \I__19200\ : InMux
    port map (
            O => \N__77579\,
            I => \N__77570\
        );

    \I__19199\ : InMux
    port map (
            O => \N__77578\,
            I => \N__77566\
        );

    \I__19198\ : Span4Mux_v
    port map (
            O => \N__77575\,
            I => \N__77563\
        );

    \I__19197\ : InMux
    port map (
            O => \N__77574\,
            I => \N__77560\
        );

    \I__19196\ : InMux
    port map (
            O => \N__77573\,
            I => \N__77557\
        );

    \I__19195\ : LocalMux
    port map (
            O => \N__77570\,
            I => \N__77554\
        );

    \I__19194\ : CascadeMux
    port map (
            O => \N__77569\,
            I => \N__77551\
        );

    \I__19193\ : LocalMux
    port map (
            O => \N__77566\,
            I => \N__77546\
        );

    \I__19192\ : Span4Mux_h
    port map (
            O => \N__77563\,
            I => \N__77546\
        );

    \I__19191\ : LocalMux
    port map (
            O => \N__77560\,
            I => \N__77543\
        );

    \I__19190\ : LocalMux
    port map (
            O => \N__77557\,
            I => \N__77538\
        );

    \I__19189\ : Span4Mux_h
    port map (
            O => \N__77554\,
            I => \N__77538\
        );

    \I__19188\ : InMux
    port map (
            O => \N__77551\,
            I => \N__77535\
        );

    \I__19187\ : Span4Mux_v
    port map (
            O => \N__77546\,
            I => \N__77532\
        );

    \I__19186\ : Span4Mux_h
    port map (
            O => \N__77543\,
            I => \N__77529\
        );

    \I__19185\ : Span4Mux_v
    port map (
            O => \N__77538\,
            I => \N__77526\
        );

    \I__19184\ : LocalMux
    port map (
            O => \N__77535\,
            I => \c0.data_in_frame_19_7\
        );

    \I__19183\ : Odrv4
    port map (
            O => \N__77532\,
            I => \c0.data_in_frame_19_7\
        );

    \I__19182\ : Odrv4
    port map (
            O => \N__77529\,
            I => \c0.data_in_frame_19_7\
        );

    \I__19181\ : Odrv4
    port map (
            O => \N__77526\,
            I => \c0.data_in_frame_19_7\
        );

    \I__19180\ : InMux
    port map (
            O => \N__77517\,
            I => \N__77514\
        );

    \I__19179\ : LocalMux
    port map (
            O => \N__77514\,
            I => \N__77511\
        );

    \I__19178\ : Odrv12
    port map (
            O => \N__77511\,
            I => \c0.n23433\
        );

    \I__19177\ : InMux
    port map (
            O => \N__77508\,
            I => \N__77505\
        );

    \I__19176\ : LocalMux
    port map (
            O => \N__77505\,
            I => \c0.n15_adj_4625\
        );

    \I__19175\ : InMux
    port map (
            O => \N__77502\,
            I => \N__77498\
        );

    \I__19174\ : InMux
    port map (
            O => \N__77501\,
            I => \N__77495\
        );

    \I__19173\ : LocalMux
    port map (
            O => \N__77498\,
            I => \c0.n17_adj_4626\
        );

    \I__19172\ : LocalMux
    port map (
            O => \N__77495\,
            I => \c0.n17_adj_4626\
        );

    \I__19171\ : InMux
    port map (
            O => \N__77490\,
            I => \N__77486\
        );

    \I__19170\ : InMux
    port map (
            O => \N__77489\,
            I => \N__77483\
        );

    \I__19169\ : LocalMux
    port map (
            O => \N__77486\,
            I => \N__77480\
        );

    \I__19168\ : LocalMux
    port map (
            O => \N__77483\,
            I => \N__77477\
        );

    \I__19167\ : Span4Mux_v
    port map (
            O => \N__77480\,
            I => \N__77474\
        );

    \I__19166\ : Span4Mux_h
    port map (
            O => \N__77477\,
            I => \N__77471\
        );

    \I__19165\ : Odrv4
    port map (
            O => \N__77474\,
            I => \c0.n16_adj_4627\
        );

    \I__19164\ : Odrv4
    port map (
            O => \N__77471\,
            I => \c0.n16_adj_4627\
        );

    \I__19163\ : CascadeMux
    port map (
            O => \N__77466\,
            I => \c0.n15_adj_4625_cascade_\
        );

    \I__19162\ : InMux
    port map (
            O => \N__77463\,
            I => \N__77460\
        );

    \I__19161\ : LocalMux
    port map (
            O => \N__77460\,
            I => \c0.n18\
        );

    \I__19160\ : InMux
    port map (
            O => \N__77457\,
            I => \N__77454\
        );

    \I__19159\ : LocalMux
    port map (
            O => \N__77454\,
            I => \N__77450\
        );

    \I__19158\ : InMux
    port map (
            O => \N__77453\,
            I => \N__77447\
        );

    \I__19157\ : Span4Mux_v
    port map (
            O => \N__77450\,
            I => \N__77441\
        );

    \I__19156\ : LocalMux
    port map (
            O => \N__77447\,
            I => \N__77441\
        );

    \I__19155\ : InMux
    port map (
            O => \N__77446\,
            I => \N__77437\
        );

    \I__19154\ : Span4Mux_v
    port map (
            O => \N__77441\,
            I => \N__77434\
        );

    \I__19153\ : InMux
    port map (
            O => \N__77440\,
            I => \N__77431\
        );

    \I__19152\ : LocalMux
    port map (
            O => \N__77437\,
            I => \N__77428\
        );

    \I__19151\ : Odrv4
    port map (
            O => \N__77434\,
            I => \c0.n22605\
        );

    \I__19150\ : LocalMux
    port map (
            O => \N__77431\,
            I => \c0.n22605\
        );

    \I__19149\ : Odrv12
    port map (
            O => \N__77428\,
            I => \c0.n22605\
        );

    \I__19148\ : InMux
    port map (
            O => \N__77421\,
            I => \N__77418\
        );

    \I__19147\ : LocalMux
    port map (
            O => \N__77418\,
            I => \N__77414\
        );

    \I__19146\ : InMux
    port map (
            O => \N__77417\,
            I => \N__77411\
        );

    \I__19145\ : Span4Mux_v
    port map (
            O => \N__77414\,
            I => \N__77406\
        );

    \I__19144\ : LocalMux
    port map (
            O => \N__77411\,
            I => \N__77406\
        );

    \I__19143\ : Span4Mux_h
    port map (
            O => \N__77406\,
            I => \N__77402\
        );

    \I__19142\ : InMux
    port map (
            O => \N__77405\,
            I => \N__77399\
        );

    \I__19141\ : Odrv4
    port map (
            O => \N__77402\,
            I => \c0.n13767\
        );

    \I__19140\ : LocalMux
    port map (
            O => \N__77399\,
            I => \c0.n13767\
        );

    \I__19139\ : CascadeMux
    port map (
            O => \N__77394\,
            I => \N__77388\
        );

    \I__19138\ : InMux
    port map (
            O => \N__77393\,
            I => \N__77383\
        );

    \I__19137\ : InMux
    port map (
            O => \N__77392\,
            I => \N__77383\
        );

    \I__19136\ : InMux
    port map (
            O => \N__77391\,
            I => \N__77380\
        );

    \I__19135\ : InMux
    port map (
            O => \N__77388\,
            I => \N__77377\
        );

    \I__19134\ : LocalMux
    port map (
            O => \N__77383\,
            I => \N__77373\
        );

    \I__19133\ : LocalMux
    port map (
            O => \N__77380\,
            I => \N__77368\
        );

    \I__19132\ : LocalMux
    port map (
            O => \N__77377\,
            I => \N__77368\
        );

    \I__19131\ : InMux
    port map (
            O => \N__77376\,
            I => \N__77365\
        );

    \I__19130\ : Span4Mux_h
    port map (
            O => \N__77373\,
            I => \N__77362\
        );

    \I__19129\ : Odrv4
    port map (
            O => \N__77368\,
            I => \c0.n13468\
        );

    \I__19128\ : LocalMux
    port map (
            O => \N__77365\,
            I => \c0.n13468\
        );

    \I__19127\ : Odrv4
    port map (
            O => \N__77362\,
            I => \c0.n13468\
        );

    \I__19126\ : CascadeMux
    port map (
            O => \N__77355\,
            I => \c0.n20239_cascade_\
        );

    \I__19125\ : InMux
    port map (
            O => \N__77352\,
            I => \N__77348\
        );

    \I__19124\ : InMux
    port map (
            O => \N__77351\,
            I => \N__77345\
        );

    \I__19123\ : LocalMux
    port map (
            O => \N__77348\,
            I => \N__77342\
        );

    \I__19122\ : LocalMux
    port map (
            O => \N__77345\,
            I => \N__77336\
        );

    \I__19121\ : Span4Mux_v
    port map (
            O => \N__77342\,
            I => \N__77336\
        );

    \I__19120\ : InMux
    port map (
            O => \N__77341\,
            I => \N__77333\
        );

    \I__19119\ : Span4Mux_h
    port map (
            O => \N__77336\,
            I => \N__77329\
        );

    \I__19118\ : LocalMux
    port map (
            O => \N__77333\,
            I => \N__77326\
        );

    \I__19117\ : CascadeMux
    port map (
            O => \N__77332\,
            I => \N__77323\
        );

    \I__19116\ : Sp12to4
    port map (
            O => \N__77329\,
            I => \N__77318\
        );

    \I__19115\ : Sp12to4
    port map (
            O => \N__77326\,
            I => \N__77318\
        );

    \I__19114\ : InMux
    port map (
            O => \N__77323\,
            I => \N__77315\
        );

    \I__19113\ : Span12Mux_s10_v
    port map (
            O => \N__77318\,
            I => \N__77312\
        );

    \I__19112\ : LocalMux
    port map (
            O => \N__77315\,
            I => \c0.data_in_frame_26_4\
        );

    \I__19111\ : Odrv12
    port map (
            O => \N__77312\,
            I => \c0.data_in_frame_26_4\
        );

    \I__19110\ : InMux
    port map (
            O => \N__77307\,
            I => \N__77304\
        );

    \I__19109\ : LocalMux
    port map (
            O => \N__77304\,
            I => \N__77301\
        );

    \I__19108\ : Odrv12
    port map (
            O => \N__77301\,
            I => \c0.n10_adj_4457\
        );

    \I__19107\ : InMux
    port map (
            O => \N__77298\,
            I => \N__77295\
        );

    \I__19106\ : LocalMux
    port map (
            O => \N__77295\,
            I => \c0.n6_adj_4668\
        );

    \I__19105\ : CascadeMux
    port map (
            O => \N__77292\,
            I => \N__77288\
        );

    \I__19104\ : InMux
    port map (
            O => \N__77291\,
            I => \N__77284\
        );

    \I__19103\ : InMux
    port map (
            O => \N__77288\,
            I => \N__77281\
        );

    \I__19102\ : InMux
    port map (
            O => \N__77287\,
            I => \N__77277\
        );

    \I__19101\ : LocalMux
    port map (
            O => \N__77284\,
            I => \N__77274\
        );

    \I__19100\ : LocalMux
    port map (
            O => \N__77281\,
            I => \N__77270\
        );

    \I__19099\ : InMux
    port map (
            O => \N__77280\,
            I => \N__77267\
        );

    \I__19098\ : LocalMux
    port map (
            O => \N__77277\,
            I => \N__77261\
        );

    \I__19097\ : Span4Mux_h
    port map (
            O => \N__77274\,
            I => \N__77261\
        );

    \I__19096\ : InMux
    port map (
            O => \N__77273\,
            I => \N__77258\
        );

    \I__19095\ : Span4Mux_v
    port map (
            O => \N__77270\,
            I => \N__77255\
        );

    \I__19094\ : LocalMux
    port map (
            O => \N__77267\,
            I => \N__77252\
        );

    \I__19093\ : InMux
    port map (
            O => \N__77266\,
            I => \N__77249\
        );

    \I__19092\ : Span4Mux_h
    port map (
            O => \N__77261\,
            I => \N__77246\
        );

    \I__19091\ : LocalMux
    port map (
            O => \N__77258\,
            I => \N__77243\
        );

    \I__19090\ : Span4Mux_h
    port map (
            O => \N__77255\,
            I => \N__77238\
        );

    \I__19089\ : Span4Mux_h
    port map (
            O => \N__77252\,
            I => \N__77238\
        );

    \I__19088\ : LocalMux
    port map (
            O => \N__77249\,
            I => \c0.data_in_frame_23_2\
        );

    \I__19087\ : Odrv4
    port map (
            O => \N__77246\,
            I => \c0.data_in_frame_23_2\
        );

    \I__19086\ : Odrv12
    port map (
            O => \N__77243\,
            I => \c0.data_in_frame_23_2\
        );

    \I__19085\ : Odrv4
    port map (
            O => \N__77238\,
            I => \c0.data_in_frame_23_2\
        );

    \I__19084\ : InMux
    port map (
            O => \N__77229\,
            I => \N__77226\
        );

    \I__19083\ : LocalMux
    port map (
            O => \N__77226\,
            I => \N__77223\
        );

    \I__19082\ : Span4Mux_h
    port map (
            O => \N__77223\,
            I => \N__77220\
        );

    \I__19081\ : Odrv4
    port map (
            O => \N__77220\,
            I => \c0.n13314\
        );

    \I__19080\ : InMux
    port map (
            O => \N__77217\,
            I => \N__77213\
        );

    \I__19079\ : InMux
    port map (
            O => \N__77216\,
            I => \N__77210\
        );

    \I__19078\ : LocalMux
    port map (
            O => \N__77213\,
            I => \N__77204\
        );

    \I__19077\ : LocalMux
    port map (
            O => \N__77210\,
            I => \N__77204\
        );

    \I__19076\ : CascadeMux
    port map (
            O => \N__77209\,
            I => \N__77201\
        );

    \I__19075\ : Span4Mux_v
    port map (
            O => \N__77204\,
            I => \N__77198\
        );

    \I__19074\ : InMux
    port map (
            O => \N__77201\,
            I => \N__77195\
        );

    \I__19073\ : Odrv4
    port map (
            O => \N__77198\,
            I => \c0.n6227\
        );

    \I__19072\ : LocalMux
    port map (
            O => \N__77195\,
            I => \c0.n6227\
        );

    \I__19071\ : InMux
    port map (
            O => \N__77190\,
            I => \N__77184\
        );

    \I__19070\ : CascadeMux
    port map (
            O => \N__77189\,
            I => \N__77181\
        );

    \I__19069\ : InMux
    port map (
            O => \N__77188\,
            I => \N__77177\
        );

    \I__19068\ : InMux
    port map (
            O => \N__77187\,
            I => \N__77174\
        );

    \I__19067\ : LocalMux
    port map (
            O => \N__77184\,
            I => \N__77171\
        );

    \I__19066\ : InMux
    port map (
            O => \N__77181\,
            I => \N__77168\
        );

    \I__19065\ : InMux
    port map (
            O => \N__77180\,
            I => \N__77165\
        );

    \I__19064\ : LocalMux
    port map (
            O => \N__77177\,
            I => \N__77162\
        );

    \I__19063\ : LocalMux
    port map (
            O => \N__77174\,
            I => data_in_frame_21_7
        );

    \I__19062\ : Odrv4
    port map (
            O => \N__77171\,
            I => data_in_frame_21_7
        );

    \I__19061\ : LocalMux
    port map (
            O => \N__77168\,
            I => data_in_frame_21_7
        );

    \I__19060\ : LocalMux
    port map (
            O => \N__77165\,
            I => data_in_frame_21_7
        );

    \I__19059\ : Odrv4
    port map (
            O => \N__77162\,
            I => data_in_frame_21_7
        );

    \I__19058\ : InMux
    port map (
            O => \N__77151\,
            I => \N__77147\
        );

    \I__19057\ : InMux
    port map (
            O => \N__77150\,
            I => \N__77144\
        );

    \I__19056\ : LocalMux
    port map (
            O => \N__77147\,
            I => \N__77141\
        );

    \I__19055\ : LocalMux
    port map (
            O => \N__77144\,
            I => \N__77138\
        );

    \I__19054\ : Odrv4
    port map (
            O => \N__77141\,
            I => \c0.n20350\
        );

    \I__19053\ : Odrv4
    port map (
            O => \N__77138\,
            I => \c0.n20350\
        );

    \I__19052\ : CascadeMux
    port map (
            O => \N__77133\,
            I => \N__77125\
        );

    \I__19051\ : CascadeMux
    port map (
            O => \N__77132\,
            I => \N__77118\
        );

    \I__19050\ : InMux
    port map (
            O => \N__77131\,
            I => \N__77115\
        );

    \I__19049\ : InMux
    port map (
            O => \N__77130\,
            I => \N__77112\
        );

    \I__19048\ : InMux
    port map (
            O => \N__77129\,
            I => \N__77107\
        );

    \I__19047\ : InMux
    port map (
            O => \N__77128\,
            I => \N__77103\
        );

    \I__19046\ : InMux
    port map (
            O => \N__77125\,
            I => \N__77093\
        );

    \I__19045\ : InMux
    port map (
            O => \N__77124\,
            I => \N__77093\
        );

    \I__19044\ : InMux
    port map (
            O => \N__77123\,
            I => \N__77087\
        );

    \I__19043\ : InMux
    port map (
            O => \N__77122\,
            I => \N__77084\
        );

    \I__19042\ : CascadeMux
    port map (
            O => \N__77121\,
            I => \N__77081\
        );

    \I__19041\ : InMux
    port map (
            O => \N__77118\,
            I => \N__77078\
        );

    \I__19040\ : LocalMux
    port map (
            O => \N__77115\,
            I => \N__77075\
        );

    \I__19039\ : LocalMux
    port map (
            O => \N__77112\,
            I => \N__77072\
        );

    \I__19038\ : InMux
    port map (
            O => \N__77111\,
            I => \N__77069\
        );

    \I__19037\ : InMux
    port map (
            O => \N__77110\,
            I => \N__77066\
        );

    \I__19036\ : LocalMux
    port map (
            O => \N__77107\,
            I => \N__77062\
        );

    \I__19035\ : InMux
    port map (
            O => \N__77106\,
            I => \N__77059\
        );

    \I__19034\ : LocalMux
    port map (
            O => \N__77103\,
            I => \N__77055\
        );

    \I__19033\ : InMux
    port map (
            O => \N__77102\,
            I => \N__77052\
        );

    \I__19032\ : InMux
    port map (
            O => \N__77101\,
            I => \N__77049\
        );

    \I__19031\ : InMux
    port map (
            O => \N__77100\,
            I => \N__77046\
        );

    \I__19030\ : CascadeMux
    port map (
            O => \N__77099\,
            I => \N__77041\
        );

    \I__19029\ : CascadeMux
    port map (
            O => \N__77098\,
            I => \N__77038\
        );

    \I__19028\ : LocalMux
    port map (
            O => \N__77093\,
            I => \N__77035\
        );

    \I__19027\ : InMux
    port map (
            O => \N__77092\,
            I => \N__77028\
        );

    \I__19026\ : InMux
    port map (
            O => \N__77091\,
            I => \N__77028\
        );

    \I__19025\ : InMux
    port map (
            O => \N__77090\,
            I => \N__77028\
        );

    \I__19024\ : LocalMux
    port map (
            O => \N__77087\,
            I => \N__77023\
        );

    \I__19023\ : LocalMux
    port map (
            O => \N__77084\,
            I => \N__77023\
        );

    \I__19022\ : InMux
    port map (
            O => \N__77081\,
            I => \N__77020\
        );

    \I__19021\ : LocalMux
    port map (
            O => \N__77078\,
            I => \N__77017\
        );

    \I__19020\ : Span4Mux_h
    port map (
            O => \N__77075\,
            I => \N__77012\
        );

    \I__19019\ : Span4Mux_h
    port map (
            O => \N__77072\,
            I => \N__77012\
        );

    \I__19018\ : LocalMux
    port map (
            O => \N__77069\,
            I => \N__77009\
        );

    \I__19017\ : LocalMux
    port map (
            O => \N__77066\,
            I => \N__77006\
        );

    \I__19016\ : InMux
    port map (
            O => \N__77065\,
            I => \N__77003\
        );

    \I__19015\ : Span4Mux_v
    port map (
            O => \N__77062\,
            I => \N__76998\
        );

    \I__19014\ : LocalMux
    port map (
            O => \N__77059\,
            I => \N__76998\
        );

    \I__19013\ : InMux
    port map (
            O => \N__77058\,
            I => \N__76994\
        );

    \I__19012\ : Span4Mux_v
    port map (
            O => \N__77055\,
            I => \N__76985\
        );

    \I__19011\ : LocalMux
    port map (
            O => \N__77052\,
            I => \N__76985\
        );

    \I__19010\ : LocalMux
    port map (
            O => \N__77049\,
            I => \N__76985\
        );

    \I__19009\ : LocalMux
    port map (
            O => \N__77046\,
            I => \N__76985\
        );

    \I__19008\ : InMux
    port map (
            O => \N__77045\,
            I => \N__76982\
        );

    \I__19007\ : InMux
    port map (
            O => \N__77044\,
            I => \N__76979\
        );

    \I__19006\ : InMux
    port map (
            O => \N__77041\,
            I => \N__76974\
        );

    \I__19005\ : InMux
    port map (
            O => \N__77038\,
            I => \N__76974\
        );

    \I__19004\ : Span4Mux_v
    port map (
            O => \N__77035\,
            I => \N__76963\
        );

    \I__19003\ : LocalMux
    port map (
            O => \N__77028\,
            I => \N__76963\
        );

    \I__19002\ : Span4Mux_h
    port map (
            O => \N__77023\,
            I => \N__76963\
        );

    \I__19001\ : LocalMux
    port map (
            O => \N__77020\,
            I => \N__76963\
        );

    \I__19000\ : Span4Mux_v
    port map (
            O => \N__77017\,
            I => \N__76963\
        );

    \I__18999\ : Span4Mux_h
    port map (
            O => \N__77012\,
            I => \N__76958\
        );

    \I__18998\ : Span4Mux_v
    port map (
            O => \N__77009\,
            I => \N__76958\
        );

    \I__18997\ : Span4Mux_v
    port map (
            O => \N__77006\,
            I => \N__76955\
        );

    \I__18996\ : LocalMux
    port map (
            O => \N__77003\,
            I => \N__76949\
        );

    \I__18995\ : Span4Mux_h
    port map (
            O => \N__76998\,
            I => \N__76949\
        );

    \I__18994\ : InMux
    port map (
            O => \N__76997\,
            I => \N__76946\
        );

    \I__18993\ : LocalMux
    port map (
            O => \N__76994\,
            I => \N__76941\
        );

    \I__18992\ : Span4Mux_h
    port map (
            O => \N__76985\,
            I => \N__76936\
        );

    \I__18991\ : LocalMux
    port map (
            O => \N__76982\,
            I => \N__76936\
        );

    \I__18990\ : LocalMux
    port map (
            O => \N__76979\,
            I => \N__76933\
        );

    \I__18989\ : LocalMux
    port map (
            O => \N__76974\,
            I => \N__76926\
        );

    \I__18988\ : Span4Mux_h
    port map (
            O => \N__76963\,
            I => \N__76926\
        );

    \I__18987\ : Span4Mux_v
    port map (
            O => \N__76958\,
            I => \N__76926\
        );

    \I__18986\ : Span4Mux_v
    port map (
            O => \N__76955\,
            I => \N__76923\
        );

    \I__18985\ : InMux
    port map (
            O => \N__76954\,
            I => \N__76920\
        );

    \I__18984\ : Span4Mux_v
    port map (
            O => \N__76949\,
            I => \N__76917\
        );

    \I__18983\ : LocalMux
    port map (
            O => \N__76946\,
            I => \N__76913\
        );

    \I__18982\ : InMux
    port map (
            O => \N__76945\,
            I => \N__76909\
        );

    \I__18981\ : InMux
    port map (
            O => \N__76944\,
            I => \N__76906\
        );

    \I__18980\ : Span4Mux_v
    port map (
            O => \N__76941\,
            I => \N__76903\
        );

    \I__18979\ : Span4Mux_h
    port map (
            O => \N__76936\,
            I => \N__76900\
        );

    \I__18978\ : Span4Mux_h
    port map (
            O => \N__76933\,
            I => \N__76895\
        );

    \I__18977\ : Span4Mux_v
    port map (
            O => \N__76926\,
            I => \N__76895\
        );

    \I__18976\ : Span4Mux_v
    port map (
            O => \N__76923\,
            I => \N__76892\
        );

    \I__18975\ : LocalMux
    port map (
            O => \N__76920\,
            I => \N__76887\
        );

    \I__18974\ : Span4Mux_v
    port map (
            O => \N__76917\,
            I => \N__76887\
        );

    \I__18973\ : CascadeMux
    port map (
            O => \N__76916\,
            I => \N__76884\
        );

    \I__18972\ : Span4Mux_v
    port map (
            O => \N__76913\,
            I => \N__76880\
        );

    \I__18971\ : InMux
    port map (
            O => \N__76912\,
            I => \N__76877\
        );

    \I__18970\ : LocalMux
    port map (
            O => \N__76909\,
            I => \N__76874\
        );

    \I__18969\ : LocalMux
    port map (
            O => \N__76906\,
            I => \N__76865\
        );

    \I__18968\ : Span4Mux_h
    port map (
            O => \N__76903\,
            I => \N__76865\
        );

    \I__18967\ : Span4Mux_v
    port map (
            O => \N__76900\,
            I => \N__76865\
        );

    \I__18966\ : Span4Mux_v
    port map (
            O => \N__76895\,
            I => \N__76865\
        );

    \I__18965\ : Span4Mux_h
    port map (
            O => \N__76892\,
            I => \N__76860\
        );

    \I__18964\ : Span4Mux_v
    port map (
            O => \N__76887\,
            I => \N__76860\
        );

    \I__18963\ : InMux
    port map (
            O => \N__76884\,
            I => \N__76855\
        );

    \I__18962\ : InMux
    port map (
            O => \N__76883\,
            I => \N__76855\
        );

    \I__18961\ : Span4Mux_v
    port map (
            O => \N__76880\,
            I => \N__76852\
        );

    \I__18960\ : LocalMux
    port map (
            O => \N__76877\,
            I => \N__76845\
        );

    \I__18959\ : Span4Mux_v
    port map (
            O => \N__76874\,
            I => \N__76845\
        );

    \I__18958\ : Span4Mux_h
    port map (
            O => \N__76865\,
            I => \N__76845\
        );

    \I__18957\ : Span4Mux_h
    port map (
            O => \N__76860\,
            I => \N__76842\
        );

    \I__18956\ : LocalMux
    port map (
            O => \N__76855\,
            I => rx_data_3
        );

    \I__18955\ : Odrv4
    port map (
            O => \N__76852\,
            I => rx_data_3
        );

    \I__18954\ : Odrv4
    port map (
            O => \N__76845\,
            I => rx_data_3
        );

    \I__18953\ : Odrv4
    port map (
            O => \N__76842\,
            I => rx_data_3
        );

    \I__18952\ : InMux
    port map (
            O => \N__76833\,
            I => \N__76829\
        );

    \I__18951\ : InMux
    port map (
            O => \N__76832\,
            I => \N__76825\
        );

    \I__18950\ : LocalMux
    port map (
            O => \N__76829\,
            I => \N__76822\
        );

    \I__18949\ : InMux
    port map (
            O => \N__76828\,
            I => \N__76819\
        );

    \I__18948\ : LocalMux
    port map (
            O => \N__76825\,
            I => \N__76816\
        );

    \I__18947\ : Span4Mux_v
    port map (
            O => \N__76822\,
            I => \N__76810\
        );

    \I__18946\ : LocalMux
    port map (
            O => \N__76819\,
            I => \N__76810\
        );

    \I__18945\ : Span4Mux_h
    port map (
            O => \N__76816\,
            I => \N__76807\
        );

    \I__18944\ : CascadeMux
    port map (
            O => \N__76815\,
            I => \N__76804\
        );

    \I__18943\ : Span4Mux_h
    port map (
            O => \N__76810\,
            I => \N__76801\
        );

    \I__18942\ : Span4Mux_h
    port map (
            O => \N__76807\,
            I => \N__76798\
        );

    \I__18941\ : InMux
    port map (
            O => \N__76804\,
            I => \N__76794\
        );

    \I__18940\ : Span4Mux_h
    port map (
            O => \N__76801\,
            I => \N__76791\
        );

    \I__18939\ : Span4Mux_v
    port map (
            O => \N__76798\,
            I => \N__76788\
        );

    \I__18938\ : InMux
    port map (
            O => \N__76797\,
            I => \N__76785\
        );

    \I__18937\ : LocalMux
    port map (
            O => \N__76794\,
            I => \c0.data_in_frame_23_3\
        );

    \I__18936\ : Odrv4
    port map (
            O => \N__76791\,
            I => \c0.data_in_frame_23_3\
        );

    \I__18935\ : Odrv4
    port map (
            O => \N__76788\,
            I => \c0.data_in_frame_23_3\
        );

    \I__18934\ : LocalMux
    port map (
            O => \N__76785\,
            I => \c0.data_in_frame_23_3\
        );

    \I__18933\ : InMux
    port map (
            O => \N__76776\,
            I => \N__76773\
        );

    \I__18932\ : LocalMux
    port map (
            O => \N__76773\,
            I => \N__76770\
        );

    \I__18931\ : Odrv4
    port map (
            O => \N__76770\,
            I => \c0.n25484\
        );

    \I__18930\ : InMux
    port map (
            O => \N__76767\,
            I => \N__76764\
        );

    \I__18929\ : LocalMux
    port map (
            O => \N__76764\,
            I => \N__76761\
        );

    \I__18928\ : Odrv4
    port map (
            O => \N__76761\,
            I => \c0.n62\
        );

    \I__18927\ : CascadeMux
    port map (
            O => \N__76758\,
            I => \N__76755\
        );

    \I__18926\ : InMux
    port map (
            O => \N__76755\,
            I => \N__76752\
        );

    \I__18925\ : LocalMux
    port map (
            O => \N__76752\,
            I => \c0.n21_adj_4481\
        );

    \I__18924\ : InMux
    port map (
            O => \N__76749\,
            I => \N__76746\
        );

    \I__18923\ : LocalMux
    port map (
            O => \N__76746\,
            I => \N__76743\
        );

    \I__18922\ : Span4Mux_v
    port map (
            O => \N__76743\,
            I => \N__76738\
        );

    \I__18921\ : InMux
    port map (
            O => \N__76742\,
            I => \N__76735\
        );

    \I__18920\ : InMux
    port map (
            O => \N__76741\,
            I => \N__76732\
        );

    \I__18919\ : Span4Mux_h
    port map (
            O => \N__76738\,
            I => \N__76727\
        );

    \I__18918\ : LocalMux
    port map (
            O => \N__76735\,
            I => \N__76727\
        );

    \I__18917\ : LocalMux
    port map (
            O => \N__76732\,
            I => \N__76723\
        );

    \I__18916\ : Span4Mux_h
    port map (
            O => \N__76727\,
            I => \N__76720\
        );

    \I__18915\ : InMux
    port map (
            O => \N__76726\,
            I => \N__76717\
        );

    \I__18914\ : Odrv12
    port map (
            O => \N__76723\,
            I => \c0.n6_adj_4462\
        );

    \I__18913\ : Odrv4
    port map (
            O => \N__76720\,
            I => \c0.n6_adj_4462\
        );

    \I__18912\ : LocalMux
    port map (
            O => \N__76717\,
            I => \c0.n6_adj_4462\
        );

    \I__18911\ : InMux
    port map (
            O => \N__76710\,
            I => \N__76707\
        );

    \I__18910\ : LocalMux
    port map (
            O => \N__76707\,
            I => \N__76704\
        );

    \I__18909\ : Span4Mux_h
    port map (
            O => \N__76704\,
            I => \N__76701\
        );

    \I__18908\ : Span4Mux_h
    port map (
            O => \N__76701\,
            I => \N__76698\
        );

    \I__18907\ : Odrv4
    port map (
            O => \N__76698\,
            I => \c0.n30_adj_4482\
        );

    \I__18906\ : InMux
    port map (
            O => \N__76695\,
            I => \N__76688\
        );

    \I__18905\ : InMux
    port map (
            O => \N__76694\,
            I => \N__76688\
        );

    \I__18904\ : InMux
    port map (
            O => \N__76693\,
            I => \N__76684\
        );

    \I__18903\ : LocalMux
    port map (
            O => \N__76688\,
            I => \N__76679\
        );

    \I__18902\ : InMux
    port map (
            O => \N__76687\,
            I => \N__76676\
        );

    \I__18901\ : LocalMux
    port map (
            O => \N__76684\,
            I => \N__76671\
        );

    \I__18900\ : InMux
    port map (
            O => \N__76683\,
            I => \N__76668\
        );

    \I__18899\ : InMux
    port map (
            O => \N__76682\,
            I => \N__76665\
        );

    \I__18898\ : Span4Mux_v
    port map (
            O => \N__76679\,
            I => \N__76660\
        );

    \I__18897\ : LocalMux
    port map (
            O => \N__76676\,
            I => \N__76660\
        );

    \I__18896\ : InMux
    port map (
            O => \N__76675\,
            I => \N__76657\
        );

    \I__18895\ : InMux
    port map (
            O => \N__76674\,
            I => \N__76649\
        );

    \I__18894\ : Span4Mux_v
    port map (
            O => \N__76671\,
            I => \N__76644\
        );

    \I__18893\ : LocalMux
    port map (
            O => \N__76668\,
            I => \N__76644\
        );

    \I__18892\ : LocalMux
    port map (
            O => \N__76665\,
            I => \N__76641\
        );

    \I__18891\ : Span4Mux_v
    port map (
            O => \N__76660\,
            I => \N__76636\
        );

    \I__18890\ : LocalMux
    port map (
            O => \N__76657\,
            I => \N__76636\
        );

    \I__18889\ : InMux
    port map (
            O => \N__76656\,
            I => \N__76631\
        );

    \I__18888\ : InMux
    port map (
            O => \N__76655\,
            I => \N__76631\
        );

    \I__18887\ : InMux
    port map (
            O => \N__76654\,
            I => \N__76626\
        );

    \I__18886\ : InMux
    port map (
            O => \N__76653\,
            I => \N__76617\
        );

    \I__18885\ : InMux
    port map (
            O => \N__76652\,
            I => \N__76617\
        );

    \I__18884\ : LocalMux
    port map (
            O => \N__76649\,
            I => \N__76614\
        );

    \I__18883\ : Span4Mux_v
    port map (
            O => \N__76644\,
            I => \N__76607\
        );

    \I__18882\ : Span4Mux_v
    port map (
            O => \N__76641\,
            I => \N__76600\
        );

    \I__18881\ : Span4Mux_v
    port map (
            O => \N__76636\,
            I => \N__76600\
        );

    \I__18880\ : LocalMux
    port map (
            O => \N__76631\,
            I => \N__76600\
        );

    \I__18879\ : CascadeMux
    port map (
            O => \N__76630\,
            I => \N__76596\
        );

    \I__18878\ : InMux
    port map (
            O => \N__76629\,
            I => \N__76592\
        );

    \I__18877\ : LocalMux
    port map (
            O => \N__76626\,
            I => \N__76589\
        );

    \I__18876\ : InMux
    port map (
            O => \N__76625\,
            I => \N__76586\
        );

    \I__18875\ : InMux
    port map (
            O => \N__76624\,
            I => \N__76583\
        );

    \I__18874\ : InMux
    port map (
            O => \N__76623\,
            I => \N__76579\
        );

    \I__18873\ : InMux
    port map (
            O => \N__76622\,
            I => \N__76576\
        );

    \I__18872\ : LocalMux
    port map (
            O => \N__76617\,
            I => \N__76573\
        );

    \I__18871\ : Span4Mux_h
    port map (
            O => \N__76614\,
            I => \N__76570\
        );

    \I__18870\ : InMux
    port map (
            O => \N__76613\,
            I => \N__76567\
        );

    \I__18869\ : InMux
    port map (
            O => \N__76612\,
            I => \N__76564\
        );

    \I__18868\ : InMux
    port map (
            O => \N__76611\,
            I => \N__76559\
        );

    \I__18867\ : InMux
    port map (
            O => \N__76610\,
            I => \N__76559\
        );

    \I__18866\ : Span4Mux_h
    port map (
            O => \N__76607\,
            I => \N__76554\
        );

    \I__18865\ : Span4Mux_h
    port map (
            O => \N__76600\,
            I => \N__76554\
        );

    \I__18864\ : CascadeMux
    port map (
            O => \N__76599\,
            I => \N__76551\
        );

    \I__18863\ : InMux
    port map (
            O => \N__76596\,
            I => \N__76545\
        );

    \I__18862\ : InMux
    port map (
            O => \N__76595\,
            I => \N__76542\
        );

    \I__18861\ : LocalMux
    port map (
            O => \N__76592\,
            I => \N__76539\
        );

    \I__18860\ : Span4Mux_v
    port map (
            O => \N__76589\,
            I => \N__76536\
        );

    \I__18859\ : LocalMux
    port map (
            O => \N__76586\,
            I => \N__76531\
        );

    \I__18858\ : LocalMux
    port map (
            O => \N__76583\,
            I => \N__76531\
        );

    \I__18857\ : InMux
    port map (
            O => \N__76582\,
            I => \N__76526\
        );

    \I__18856\ : LocalMux
    port map (
            O => \N__76579\,
            I => \N__76520\
        );

    \I__18855\ : LocalMux
    port map (
            O => \N__76576\,
            I => \N__76520\
        );

    \I__18854\ : Span4Mux_v
    port map (
            O => \N__76573\,
            I => \N__76513\
        );

    \I__18853\ : Span4Mux_h
    port map (
            O => \N__76570\,
            I => \N__76513\
        );

    \I__18852\ : LocalMux
    port map (
            O => \N__76567\,
            I => \N__76513\
        );

    \I__18851\ : LocalMux
    port map (
            O => \N__76564\,
            I => \N__76510\
        );

    \I__18850\ : LocalMux
    port map (
            O => \N__76559\,
            I => \N__76505\
        );

    \I__18849\ : Span4Mux_v
    port map (
            O => \N__76554\,
            I => \N__76505\
        );

    \I__18848\ : InMux
    port map (
            O => \N__76551\,
            I => \N__76502\
        );

    \I__18847\ : InMux
    port map (
            O => \N__76550\,
            I => \N__76499\
        );

    \I__18846\ : InMux
    port map (
            O => \N__76549\,
            I => \N__76496\
        );

    \I__18845\ : InMux
    port map (
            O => \N__76548\,
            I => \N__76493\
        );

    \I__18844\ : LocalMux
    port map (
            O => \N__76545\,
            I => \N__76484\
        );

    \I__18843\ : LocalMux
    port map (
            O => \N__76542\,
            I => \N__76484\
        );

    \I__18842\ : Span4Mux_h
    port map (
            O => \N__76539\,
            I => \N__76484\
        );

    \I__18841\ : Span4Mux_v
    port map (
            O => \N__76536\,
            I => \N__76484\
        );

    \I__18840\ : Span4Mux_v
    port map (
            O => \N__76531\,
            I => \N__76481\
        );

    \I__18839\ : InMux
    port map (
            O => \N__76530\,
            I => \N__76478\
        );

    \I__18838\ : InMux
    port map (
            O => \N__76529\,
            I => \N__76475\
        );

    \I__18837\ : LocalMux
    port map (
            O => \N__76526\,
            I => \N__76472\
        );

    \I__18836\ : InMux
    port map (
            O => \N__76525\,
            I => \N__76469\
        );

    \I__18835\ : Span4Mux_v
    port map (
            O => \N__76520\,
            I => \N__76464\
        );

    \I__18834\ : Span4Mux_v
    port map (
            O => \N__76513\,
            I => \N__76464\
        );

    \I__18833\ : Span4Mux_h
    port map (
            O => \N__76510\,
            I => \N__76459\
        );

    \I__18832\ : Span4Mux_v
    port map (
            O => \N__76505\,
            I => \N__76459\
        );

    \I__18831\ : LocalMux
    port map (
            O => \N__76502\,
            I => \N__76456\
        );

    \I__18830\ : LocalMux
    port map (
            O => \N__76499\,
            I => \N__76449\
        );

    \I__18829\ : LocalMux
    port map (
            O => \N__76496\,
            I => \N__76449\
        );

    \I__18828\ : LocalMux
    port map (
            O => \N__76493\,
            I => \N__76449\
        );

    \I__18827\ : Span4Mux_h
    port map (
            O => \N__76484\,
            I => \N__76446\
        );

    \I__18826\ : Sp12to4
    port map (
            O => \N__76481\,
            I => \N__76443\
        );

    \I__18825\ : LocalMux
    port map (
            O => \N__76478\,
            I => \N__76434\
        );

    \I__18824\ : LocalMux
    port map (
            O => \N__76475\,
            I => \N__76434\
        );

    \I__18823\ : Span12Mux_v
    port map (
            O => \N__76472\,
            I => \N__76434\
        );

    \I__18822\ : LocalMux
    port map (
            O => \N__76469\,
            I => \N__76434\
        );

    \I__18821\ : Span4Mux_h
    port map (
            O => \N__76464\,
            I => \N__76429\
        );

    \I__18820\ : Span4Mux_v
    port map (
            O => \N__76459\,
            I => \N__76429\
        );

    \I__18819\ : Span4Mux_v
    port map (
            O => \N__76456\,
            I => \N__76426\
        );

    \I__18818\ : Span4Mux_v
    port map (
            O => \N__76449\,
            I => \N__76423\
        );

    \I__18817\ : Span4Mux_h
    port map (
            O => \N__76446\,
            I => \N__76420\
        );

    \I__18816\ : Span12Mux_h
    port map (
            O => \N__76443\,
            I => \N__76417\
        );

    \I__18815\ : Span12Mux_v
    port map (
            O => \N__76434\,
            I => \N__76414\
        );

    \I__18814\ : Span4Mux_v
    port map (
            O => \N__76429\,
            I => \N__76411\
        );

    \I__18813\ : Odrv4
    port map (
            O => \N__76426\,
            I => \c0.n9_adj_4273\
        );

    \I__18812\ : Odrv4
    port map (
            O => \N__76423\,
            I => \c0.n9_adj_4273\
        );

    \I__18811\ : Odrv4
    port map (
            O => \N__76420\,
            I => \c0.n9_adj_4273\
        );

    \I__18810\ : Odrv12
    port map (
            O => \N__76417\,
            I => \c0.n9_adj_4273\
        );

    \I__18809\ : Odrv12
    port map (
            O => \N__76414\,
            I => \c0.n9_adj_4273\
        );

    \I__18808\ : Odrv4
    port map (
            O => \N__76411\,
            I => \c0.n9_adj_4273\
        );

    \I__18807\ : CascadeMux
    port map (
            O => \N__76398\,
            I => \N__76395\
        );

    \I__18806\ : InMux
    port map (
            O => \N__76395\,
            I => \N__76390\
        );

    \I__18805\ : InMux
    port map (
            O => \N__76394\,
            I => \N__76386\
        );

    \I__18804\ : InMux
    port map (
            O => \N__76393\,
            I => \N__76379\
        );

    \I__18803\ : LocalMux
    port map (
            O => \N__76390\,
            I => \N__76375\
        );

    \I__18802\ : InMux
    port map (
            O => \N__76389\,
            I => \N__76372\
        );

    \I__18801\ : LocalMux
    port map (
            O => \N__76386\,
            I => \N__76369\
        );

    \I__18800\ : InMux
    port map (
            O => \N__76385\,
            I => \N__76366\
        );

    \I__18799\ : InMux
    port map (
            O => \N__76384\,
            I => \N__76362\
        );

    \I__18798\ : CascadeMux
    port map (
            O => \N__76383\,
            I => \N__76359\
        );

    \I__18797\ : CascadeMux
    port map (
            O => \N__76382\,
            I => \N__76356\
        );

    \I__18796\ : LocalMux
    port map (
            O => \N__76379\,
            I => \N__76351\
        );

    \I__18795\ : InMux
    port map (
            O => \N__76378\,
            I => \N__76348\
        );

    \I__18794\ : Span4Mux_h
    port map (
            O => \N__76375\,
            I => \N__76343\
        );

    \I__18793\ : LocalMux
    port map (
            O => \N__76372\,
            I => \N__76343\
        );

    \I__18792\ : Span4Mux_v
    port map (
            O => \N__76369\,
            I => \N__76338\
        );

    \I__18791\ : LocalMux
    port map (
            O => \N__76366\,
            I => \N__76338\
        );

    \I__18790\ : CascadeMux
    port map (
            O => \N__76365\,
            I => \N__76335\
        );

    \I__18789\ : LocalMux
    port map (
            O => \N__76362\,
            I => \N__76332\
        );

    \I__18788\ : InMux
    port map (
            O => \N__76359\,
            I => \N__76329\
        );

    \I__18787\ : InMux
    port map (
            O => \N__76356\,
            I => \N__76326\
        );

    \I__18786\ : InMux
    port map (
            O => \N__76355\,
            I => \N__76321\
        );

    \I__18785\ : InMux
    port map (
            O => \N__76354\,
            I => \N__76318\
        );

    \I__18784\ : Span4Mux_v
    port map (
            O => \N__76351\,
            I => \N__76310\
        );

    \I__18783\ : LocalMux
    port map (
            O => \N__76348\,
            I => \N__76310\
        );

    \I__18782\ : Span4Mux_v
    port map (
            O => \N__76343\,
            I => \N__76305\
        );

    \I__18781\ : Span4Mux_h
    port map (
            O => \N__76338\,
            I => \N__76305\
        );

    \I__18780\ : InMux
    port map (
            O => \N__76335\,
            I => \N__76302\
        );

    \I__18779\ : Span4Mux_h
    port map (
            O => \N__76332\,
            I => \N__76295\
        );

    \I__18778\ : LocalMux
    port map (
            O => \N__76329\,
            I => \N__76295\
        );

    \I__18777\ : LocalMux
    port map (
            O => \N__76326\,
            I => \N__76295\
        );

    \I__18776\ : CascadeMux
    port map (
            O => \N__76325\,
            I => \N__76290\
        );

    \I__18775\ : InMux
    port map (
            O => \N__76324\,
            I => \N__76286\
        );

    \I__18774\ : LocalMux
    port map (
            O => \N__76321\,
            I => \N__76282\
        );

    \I__18773\ : LocalMux
    port map (
            O => \N__76318\,
            I => \N__76279\
        );

    \I__18772\ : InMux
    port map (
            O => \N__76317\,
            I => \N__76276\
        );

    \I__18771\ : InMux
    port map (
            O => \N__76316\,
            I => \N__76271\
        );

    \I__18770\ : InMux
    port map (
            O => \N__76315\,
            I => \N__76268\
        );

    \I__18769\ : Span4Mux_v
    port map (
            O => \N__76310\,
            I => \N__76265\
        );

    \I__18768\ : Span4Mux_h
    port map (
            O => \N__76305\,
            I => \N__76260\
        );

    \I__18767\ : LocalMux
    port map (
            O => \N__76302\,
            I => \N__76260\
        );

    \I__18766\ : Span4Mux_v
    port map (
            O => \N__76295\,
            I => \N__76257\
        );

    \I__18765\ : CascadeMux
    port map (
            O => \N__76294\,
            I => \N__76254\
        );

    \I__18764\ : InMux
    port map (
            O => \N__76293\,
            I => \N__76251\
        );

    \I__18763\ : InMux
    port map (
            O => \N__76290\,
            I => \N__76248\
        );

    \I__18762\ : InMux
    port map (
            O => \N__76289\,
            I => \N__76245\
        );

    \I__18761\ : LocalMux
    port map (
            O => \N__76286\,
            I => \N__76242\
        );

    \I__18760\ : InMux
    port map (
            O => \N__76285\,
            I => \N__76239\
        );

    \I__18759\ : Span4Mux_v
    port map (
            O => \N__76282\,
            I => \N__76232\
        );

    \I__18758\ : Span4Mux_h
    port map (
            O => \N__76279\,
            I => \N__76232\
        );

    \I__18757\ : LocalMux
    port map (
            O => \N__76276\,
            I => \N__76232\
        );

    \I__18756\ : CascadeMux
    port map (
            O => \N__76275\,
            I => \N__76229\
        );

    \I__18755\ : InMux
    port map (
            O => \N__76274\,
            I => \N__76224\
        );

    \I__18754\ : LocalMux
    port map (
            O => \N__76271\,
            I => \N__76221\
        );

    \I__18753\ : LocalMux
    port map (
            O => \N__76268\,
            I => \N__76218\
        );

    \I__18752\ : Span4Mux_h
    port map (
            O => \N__76265\,
            I => \N__76215\
        );

    \I__18751\ : Span4Mux_v
    port map (
            O => \N__76260\,
            I => \N__76212\
        );

    \I__18750\ : Span4Mux_h
    port map (
            O => \N__76257\,
            I => \N__76209\
        );

    \I__18749\ : InMux
    port map (
            O => \N__76254\,
            I => \N__76206\
        );

    \I__18748\ : LocalMux
    port map (
            O => \N__76251\,
            I => \N__76199\
        );

    \I__18747\ : LocalMux
    port map (
            O => \N__76248\,
            I => \N__76199\
        );

    \I__18746\ : LocalMux
    port map (
            O => \N__76245\,
            I => \N__76199\
        );

    \I__18745\ : Span4Mux_v
    port map (
            O => \N__76242\,
            I => \N__76194\
        );

    \I__18744\ : LocalMux
    port map (
            O => \N__76239\,
            I => \N__76194\
        );

    \I__18743\ : Span4Mux_v
    port map (
            O => \N__76232\,
            I => \N__76191\
        );

    \I__18742\ : InMux
    port map (
            O => \N__76229\,
            I => \N__76188\
        );

    \I__18741\ : InMux
    port map (
            O => \N__76228\,
            I => \N__76183\
        );

    \I__18740\ : InMux
    port map (
            O => \N__76227\,
            I => \N__76183\
        );

    \I__18739\ : LocalMux
    port map (
            O => \N__76224\,
            I => \N__76180\
        );

    \I__18738\ : Span4Mux_v
    port map (
            O => \N__76221\,
            I => \N__76175\
        );

    \I__18737\ : Span4Mux_h
    port map (
            O => \N__76218\,
            I => \N__76175\
        );

    \I__18736\ : Sp12to4
    port map (
            O => \N__76215\,
            I => \N__76172\
        );

    \I__18735\ : Sp12to4
    port map (
            O => \N__76212\,
            I => \N__76167\
        );

    \I__18734\ : Sp12to4
    port map (
            O => \N__76209\,
            I => \N__76167\
        );

    \I__18733\ : LocalMux
    port map (
            O => \N__76206\,
            I => \N__76164\
        );

    \I__18732\ : Span4Mux_v
    port map (
            O => \N__76199\,
            I => \N__76161\
        );

    \I__18731\ : Span4Mux_h
    port map (
            O => \N__76194\,
            I => \N__76158\
        );

    \I__18730\ : Span4Mux_h
    port map (
            O => \N__76191\,
            I => \N__76155\
        );

    \I__18729\ : LocalMux
    port map (
            O => \N__76188\,
            I => \N__76135\
        );

    \I__18728\ : LocalMux
    port map (
            O => \N__76183\,
            I => \N__76135\
        );

    \I__18727\ : Span12Mux_h
    port map (
            O => \N__76180\,
            I => \N__76135\
        );

    \I__18726\ : Sp12to4
    port map (
            O => \N__76175\,
            I => \N__76135\
        );

    \I__18725\ : Span12Mux_h
    port map (
            O => \N__76172\,
            I => \N__76135\
        );

    \I__18724\ : Span12Mux_h
    port map (
            O => \N__76167\,
            I => \N__76135\
        );

    \I__18723\ : Span4Mux_v
    port map (
            O => \N__76164\,
            I => \N__76130\
        );

    \I__18722\ : Span4Mux_v
    port map (
            O => \N__76161\,
            I => \N__76130\
        );

    \I__18721\ : Span4Mux_v
    port map (
            O => \N__76158\,
            I => \N__76125\
        );

    \I__18720\ : Span4Mux_v
    port map (
            O => \N__76155\,
            I => \N__76125\
        );

    \I__18719\ : InMux
    port map (
            O => \N__76154\,
            I => \N__76122\
        );

    \I__18718\ : InMux
    port map (
            O => \N__76153\,
            I => \N__76117\
        );

    \I__18717\ : InMux
    port map (
            O => \N__76152\,
            I => \N__76117\
        );

    \I__18716\ : InMux
    port map (
            O => \N__76151\,
            I => \N__76112\
        );

    \I__18715\ : InMux
    port map (
            O => \N__76150\,
            I => \N__76112\
        );

    \I__18714\ : InMux
    port map (
            O => \N__76149\,
            I => \N__76107\
        );

    \I__18713\ : InMux
    port map (
            O => \N__76148\,
            I => \N__76107\
        );

    \I__18712\ : Span12Mux_v
    port map (
            O => \N__76135\,
            I => \N__76104\
        );

    \I__18711\ : Span4Mux_h
    port map (
            O => \N__76130\,
            I => \N__76099\
        );

    \I__18710\ : Span4Mux_v
    port map (
            O => \N__76125\,
            I => \N__76099\
        );

    \I__18709\ : LocalMux
    port map (
            O => \N__76122\,
            I => rx_data_7
        );

    \I__18708\ : LocalMux
    port map (
            O => \N__76117\,
            I => rx_data_7
        );

    \I__18707\ : LocalMux
    port map (
            O => \N__76112\,
            I => rx_data_7
        );

    \I__18706\ : LocalMux
    port map (
            O => \N__76107\,
            I => rx_data_7
        );

    \I__18705\ : Odrv12
    port map (
            O => \N__76104\,
            I => rx_data_7
        );

    \I__18704\ : Odrv4
    port map (
            O => \N__76099\,
            I => rx_data_7
        );

    \I__18703\ : InMux
    port map (
            O => \N__76086\,
            I => \N__76083\
        );

    \I__18702\ : LocalMux
    port map (
            O => \N__76083\,
            I => \N__76079\
        );

    \I__18701\ : InMux
    port map (
            O => \N__76082\,
            I => \N__76076\
        );

    \I__18700\ : Span4Mux_h
    port map (
            O => \N__76079\,
            I => \N__76071\
        );

    \I__18699\ : LocalMux
    port map (
            O => \N__76076\,
            I => \N__76071\
        );

    \I__18698\ : Span4Mux_h
    port map (
            O => \N__76071\,
            I => \N__76067\
        );

    \I__18697\ : CascadeMux
    port map (
            O => \N__76070\,
            I => \N__76064\
        );

    \I__18696\ : Sp12to4
    port map (
            O => \N__76067\,
            I => \N__76061\
        );

    \I__18695\ : InMux
    port map (
            O => \N__76064\,
            I => \N__76058\
        );

    \I__18694\ : Odrv12
    port map (
            O => \N__76061\,
            I => \c0.n23598\
        );

    \I__18693\ : LocalMux
    port map (
            O => \N__76058\,
            I => \c0.n23598\
        );

    \I__18692\ : InMux
    port map (
            O => \N__76053\,
            I => \N__76049\
        );

    \I__18691\ : InMux
    port map (
            O => \N__76052\,
            I => \N__76044\
        );

    \I__18690\ : LocalMux
    port map (
            O => \N__76049\,
            I => \N__76041\
        );

    \I__18689\ : CascadeMux
    port map (
            O => \N__76048\,
            I => \N__76038\
        );

    \I__18688\ : CascadeMux
    port map (
            O => \N__76047\,
            I => \N__76033\
        );

    \I__18687\ : LocalMux
    port map (
            O => \N__76044\,
            I => \N__76030\
        );

    \I__18686\ : Span4Mux_v
    port map (
            O => \N__76041\,
            I => \N__76027\
        );

    \I__18685\ : InMux
    port map (
            O => \N__76038\,
            I => \N__76022\
        );

    \I__18684\ : InMux
    port map (
            O => \N__76037\,
            I => \N__76022\
        );

    \I__18683\ : InMux
    port map (
            O => \N__76036\,
            I => \N__76019\
        );

    \I__18682\ : InMux
    port map (
            O => \N__76033\,
            I => \N__76016\
        );

    \I__18681\ : Span4Mux_h
    port map (
            O => \N__76030\,
            I => \N__76013\
        );

    \I__18680\ : Span4Mux_h
    port map (
            O => \N__76027\,
            I => \N__76008\
        );

    \I__18679\ : LocalMux
    port map (
            O => \N__76022\,
            I => \N__76008\
        );

    \I__18678\ : LocalMux
    port map (
            O => \N__76019\,
            I => \N__76005\
        );

    \I__18677\ : LocalMux
    port map (
            O => \N__76016\,
            I => \c0.data_in_frame_8_4\
        );

    \I__18676\ : Odrv4
    port map (
            O => \N__76013\,
            I => \c0.data_in_frame_8_4\
        );

    \I__18675\ : Odrv4
    port map (
            O => \N__76008\,
            I => \c0.data_in_frame_8_4\
        );

    \I__18674\ : Odrv12
    port map (
            O => \N__76005\,
            I => \c0.data_in_frame_8_4\
        );

    \I__18673\ : CascadeMux
    port map (
            O => \N__75996\,
            I => \N__75993\
        );

    \I__18672\ : InMux
    port map (
            O => \N__75993\,
            I => \N__75990\
        );

    \I__18671\ : LocalMux
    port map (
            O => \N__75990\,
            I => \N__75986\
        );

    \I__18670\ : CascadeMux
    port map (
            O => \N__75989\,
            I => \N__75983\
        );

    \I__18669\ : Span12Mux_s10_h
    port map (
            O => \N__75986\,
            I => \N__75980\
        );

    \I__18668\ : InMux
    port map (
            O => \N__75983\,
            I => \N__75977\
        );

    \I__18667\ : Span12Mux_v
    port map (
            O => \N__75980\,
            I => \N__75974\
        );

    \I__18666\ : LocalMux
    port map (
            O => \N__75977\,
            I => \c0.data_in_frame_26_6\
        );

    \I__18665\ : Odrv12
    port map (
            O => \N__75974\,
            I => \c0.data_in_frame_26_6\
        );

    \I__18664\ : InMux
    port map (
            O => \N__75969\,
            I => \N__75966\
        );

    \I__18663\ : LocalMux
    port map (
            O => \N__75966\,
            I => \N__75963\
        );

    \I__18662\ : Span12Mux_h
    port map (
            O => \N__75963\,
            I => \N__75959\
        );

    \I__18661\ : InMux
    port map (
            O => \N__75962\,
            I => \N__75956\
        );

    \I__18660\ : Odrv12
    port map (
            O => \N__75959\,
            I => \c0.n22769\
        );

    \I__18659\ : LocalMux
    port map (
            O => \N__75956\,
            I => \c0.n22769\
        );

    \I__18658\ : InMux
    port map (
            O => \N__75951\,
            I => \N__75948\
        );

    \I__18657\ : LocalMux
    port map (
            O => \N__75948\,
            I => \N__75943\
        );

    \I__18656\ : InMux
    port map (
            O => \N__75947\,
            I => \N__75940\
        );

    \I__18655\ : InMux
    port map (
            O => \N__75946\,
            I => \N__75935\
        );

    \I__18654\ : Span4Mux_h
    port map (
            O => \N__75943\,
            I => \N__75932\
        );

    \I__18653\ : LocalMux
    port map (
            O => \N__75940\,
            I => \N__75929\
        );

    \I__18652\ : InMux
    port map (
            O => \N__75939\,
            I => \N__75926\
        );

    \I__18651\ : CascadeMux
    port map (
            O => \N__75938\,
            I => \N__75923\
        );

    \I__18650\ : LocalMux
    port map (
            O => \N__75935\,
            I => \N__75920\
        );

    \I__18649\ : Span4Mux_v
    port map (
            O => \N__75932\,
            I => \N__75913\
        );

    \I__18648\ : Span4Mux_h
    port map (
            O => \N__75929\,
            I => \N__75913\
        );

    \I__18647\ : LocalMux
    port map (
            O => \N__75926\,
            I => \N__75913\
        );

    \I__18646\ : InMux
    port map (
            O => \N__75923\,
            I => \N__75910\
        );

    \I__18645\ : Span4Mux_h
    port map (
            O => \N__75920\,
            I => \N__75906\
        );

    \I__18644\ : Span4Mux_v
    port map (
            O => \N__75913\,
            I => \N__75903\
        );

    \I__18643\ : LocalMux
    port map (
            O => \N__75910\,
            I => \N__75900\
        );

    \I__18642\ : InMux
    port map (
            O => \N__75909\,
            I => \N__75897\
        );

    \I__18641\ : Span4Mux_h
    port map (
            O => \N__75906\,
            I => \N__75894\
        );

    \I__18640\ : Span4Mux_h
    port map (
            O => \N__75903\,
            I => \N__75891\
        );

    \I__18639\ : Span12Mux_v
    port map (
            O => \N__75900\,
            I => \N__75888\
        );

    \I__18638\ : LocalMux
    port map (
            O => \N__75897\,
            I => \N__75883\
        );

    \I__18637\ : Span4Mux_v
    port map (
            O => \N__75894\,
            I => \N__75883\
        );

    \I__18636\ : Span4Mux_h
    port map (
            O => \N__75891\,
            I => \N__75880\
        );

    \I__18635\ : Odrv12
    port map (
            O => \N__75888\,
            I => data_in_frame_21_5
        );

    \I__18634\ : Odrv4
    port map (
            O => \N__75883\,
            I => data_in_frame_21_5
        );

    \I__18633\ : Odrv4
    port map (
            O => \N__75880\,
            I => data_in_frame_21_5
        );

    \I__18632\ : InMux
    port map (
            O => \N__75873\,
            I => \N__75870\
        );

    \I__18631\ : LocalMux
    port map (
            O => \N__75870\,
            I => \N__75867\
        );

    \I__18630\ : Span4Mux_v
    port map (
            O => \N__75867\,
            I => \N__75864\
        );

    \I__18629\ : Span4Mux_h
    port map (
            O => \N__75864\,
            I => \N__75861\
        );

    \I__18628\ : Odrv4
    port map (
            O => \N__75861\,
            I => \c0.n22698\
        );

    \I__18627\ : CascadeMux
    port map (
            O => \N__75858\,
            I => \N__75854\
        );

    \I__18626\ : CascadeMux
    port map (
            O => \N__75857\,
            I => \N__75851\
        );

    \I__18625\ : InMux
    port map (
            O => \N__75854\,
            I => \N__75848\
        );

    \I__18624\ : InMux
    port map (
            O => \N__75851\,
            I => \N__75844\
        );

    \I__18623\ : LocalMux
    port map (
            O => \N__75848\,
            I => \N__75841\
        );

    \I__18622\ : InMux
    port map (
            O => \N__75847\,
            I => \N__75838\
        );

    \I__18621\ : LocalMux
    port map (
            O => \N__75844\,
            I => \N__75831\
        );

    \I__18620\ : Span4Mux_v
    port map (
            O => \N__75841\,
            I => \N__75831\
        );

    \I__18619\ : LocalMux
    port map (
            O => \N__75838\,
            I => \N__75831\
        );

    \I__18618\ : Span4Mux_h
    port map (
            O => \N__75831\,
            I => \N__75827\
        );

    \I__18617\ : CascadeMux
    port map (
            O => \N__75830\,
            I => \N__75824\
        );

    \I__18616\ : Span4Mux_h
    port map (
            O => \N__75827\,
            I => \N__75820\
        );

    \I__18615\ : InMux
    port map (
            O => \N__75824\,
            I => \N__75815\
        );

    \I__18614\ : InMux
    port map (
            O => \N__75823\,
            I => \N__75815\
        );

    \I__18613\ : Odrv4
    port map (
            O => \N__75820\,
            I => \c0.data_in_frame_23_6\
        );

    \I__18612\ : LocalMux
    port map (
            O => \N__75815\,
            I => \c0.data_in_frame_23_6\
        );

    \I__18611\ : InMux
    port map (
            O => \N__75810\,
            I => \N__75807\
        );

    \I__18610\ : LocalMux
    port map (
            O => \N__75807\,
            I => \N__75804\
        );

    \I__18609\ : Span4Mux_h
    port map (
            O => \N__75804\,
            I => \N__75801\
        );

    \I__18608\ : Span4Mux_h
    port map (
            O => \N__75801\,
            I => \N__75798\
        );

    \I__18607\ : Odrv4
    port map (
            O => \N__75798\,
            I => \c0.n4_adj_4464\
        );

    \I__18606\ : InMux
    port map (
            O => \N__75795\,
            I => \N__75792\
        );

    \I__18605\ : LocalMux
    port map (
            O => \N__75792\,
            I => \N__75789\
        );

    \I__18604\ : Odrv12
    port map (
            O => \N__75789\,
            I => \c0.n14_adj_4465\
        );

    \I__18603\ : InMux
    port map (
            O => \N__75786\,
            I => \N__75779\
        );

    \I__18602\ : InMux
    port map (
            O => \N__75785\,
            I => \N__75779\
        );

    \I__18601\ : InMux
    port map (
            O => \N__75784\,
            I => \N__75775\
        );

    \I__18600\ : LocalMux
    port map (
            O => \N__75779\,
            I => \N__75772\
        );

    \I__18599\ : InMux
    port map (
            O => \N__75778\,
            I => \N__75769\
        );

    \I__18598\ : LocalMux
    port map (
            O => \N__75775\,
            I => \N__75766\
        );

    \I__18597\ : Span4Mux_h
    port map (
            O => \N__75772\,
            I => \N__75762\
        );

    \I__18596\ : LocalMux
    port map (
            O => \N__75769\,
            I => \N__75757\
        );

    \I__18595\ : Span4Mux_h
    port map (
            O => \N__75766\,
            I => \N__75757\
        );

    \I__18594\ : CascadeMux
    port map (
            O => \N__75765\,
            I => \N__75754\
        );

    \I__18593\ : Sp12to4
    port map (
            O => \N__75762\,
            I => \N__75751\
        );

    \I__18592\ : Span4Mux_v
    port map (
            O => \N__75757\,
            I => \N__75748\
        );

    \I__18591\ : InMux
    port map (
            O => \N__75754\,
            I => \N__75745\
        );

    \I__18590\ : Span12Mux_v
    port map (
            O => \N__75751\,
            I => \N__75742\
        );

    \I__18589\ : Span4Mux_v
    port map (
            O => \N__75748\,
            I => \N__75739\
        );

    \I__18588\ : LocalMux
    port map (
            O => \N__75745\,
            I => \c0.data_in_frame_20_3\
        );

    \I__18587\ : Odrv12
    port map (
            O => \N__75742\,
            I => \c0.data_in_frame_20_3\
        );

    \I__18586\ : Odrv4
    port map (
            O => \N__75739\,
            I => \c0.data_in_frame_20_3\
        );

    \I__18585\ : InMux
    port map (
            O => \N__75732\,
            I => \N__75726\
        );

    \I__18584\ : InMux
    port map (
            O => \N__75731\,
            I => \N__75719\
        );

    \I__18583\ : InMux
    port map (
            O => \N__75730\,
            I => \N__75719\
        );

    \I__18582\ : InMux
    port map (
            O => \N__75729\,
            I => \N__75719\
        );

    \I__18581\ : LocalMux
    port map (
            O => \N__75726\,
            I => \N__75716\
        );

    \I__18580\ : LocalMux
    port map (
            O => \N__75719\,
            I => \N__75713\
        );

    \I__18579\ : Odrv12
    port map (
            O => \N__75716\,
            I => \c0.n21412\
        );

    \I__18578\ : Odrv4
    port map (
            O => \N__75713\,
            I => \c0.n21412\
        );

    \I__18577\ : InMux
    port map (
            O => \N__75708\,
            I => \N__75705\
        );

    \I__18576\ : LocalMux
    port map (
            O => \N__75705\,
            I => \c0.n4_adj_4369\
        );

    \I__18575\ : CascadeMux
    port map (
            O => \N__75702\,
            I => \N__75697\
        );

    \I__18574\ : CascadeMux
    port map (
            O => \N__75701\,
            I => \N__75694\
        );

    \I__18573\ : CascadeMux
    port map (
            O => \N__75700\,
            I => \N__75691\
        );

    \I__18572\ : InMux
    port map (
            O => \N__75697\,
            I => \N__75688\
        );

    \I__18571\ : InMux
    port map (
            O => \N__75694\,
            I => \N__75685\
        );

    \I__18570\ : InMux
    port map (
            O => \N__75691\,
            I => \N__75682\
        );

    \I__18569\ : LocalMux
    port map (
            O => \N__75688\,
            I => \N__75679\
        );

    \I__18568\ : LocalMux
    port map (
            O => \N__75685\,
            I => \N__75675\
        );

    \I__18567\ : LocalMux
    port map (
            O => \N__75682\,
            I => \N__75672\
        );

    \I__18566\ : Span4Mux_h
    port map (
            O => \N__75679\,
            I => \N__75669\
        );

    \I__18565\ : CascadeMux
    port map (
            O => \N__75678\,
            I => \N__75666\
        );

    \I__18564\ : Span4Mux_h
    port map (
            O => \N__75675\,
            I => \N__75663\
        );

    \I__18563\ : Span4Mux_h
    port map (
            O => \N__75672\,
            I => \N__75660\
        );

    \I__18562\ : Span4Mux_h
    port map (
            O => \N__75669\,
            I => \N__75657\
        );

    \I__18561\ : InMux
    port map (
            O => \N__75666\,
            I => \N__75654\
        );

    \I__18560\ : Span4Mux_h
    port map (
            O => \N__75663\,
            I => \N__75649\
        );

    \I__18559\ : Span4Mux_h
    port map (
            O => \N__75660\,
            I => \N__75649\
        );

    \I__18558\ : Span4Mux_v
    port map (
            O => \N__75657\,
            I => \N__75646\
        );

    \I__18557\ : LocalMux
    port map (
            O => \N__75654\,
            I => \N__75641\
        );

    \I__18556\ : Span4Mux_v
    port map (
            O => \N__75649\,
            I => \N__75641\
        );

    \I__18555\ : Odrv4
    port map (
            O => \N__75646\,
            I => \c0.data_in_frame_27_0\
        );

    \I__18554\ : Odrv4
    port map (
            O => \N__75641\,
            I => \c0.data_in_frame_27_0\
        );

    \I__18553\ : CascadeMux
    port map (
            O => \N__75636\,
            I => \N__75633\
        );

    \I__18552\ : InMux
    port map (
            O => \N__75633\,
            I => \N__75630\
        );

    \I__18551\ : LocalMux
    port map (
            O => \N__75630\,
            I => \N__75627\
        );

    \I__18550\ : Span4Mux_h
    port map (
            O => \N__75627\,
            I => \N__75624\
        );

    \I__18549\ : Odrv4
    port map (
            O => \N__75624\,
            I => \c0.n73\
        );

    \I__18548\ : InMux
    port map (
            O => \N__75621\,
            I => \N__75615\
        );

    \I__18547\ : InMux
    port map (
            O => \N__75620\,
            I => \N__75615\
        );

    \I__18546\ : LocalMux
    port map (
            O => \N__75615\,
            I => \N__75608\
        );

    \I__18545\ : InMux
    port map (
            O => \N__75614\,
            I => \N__75605\
        );

    \I__18544\ : InMux
    port map (
            O => \N__75613\,
            I => \N__75600\
        );

    \I__18543\ : InMux
    port map (
            O => \N__75612\,
            I => \N__75600\
        );

    \I__18542\ : InMux
    port map (
            O => \N__75611\,
            I => \N__75597\
        );

    \I__18541\ : Span4Mux_v
    port map (
            O => \N__75608\,
            I => \N__75590\
        );

    \I__18540\ : LocalMux
    port map (
            O => \N__75605\,
            I => \N__75590\
        );

    \I__18539\ : LocalMux
    port map (
            O => \N__75600\,
            I => \N__75590\
        );

    \I__18538\ : LocalMux
    port map (
            O => \N__75597\,
            I => \N__75587\
        );

    \I__18537\ : Span4Mux_h
    port map (
            O => \N__75590\,
            I => \N__75584\
        );

    \I__18536\ : Span4Mux_v
    port map (
            O => \N__75587\,
            I => \N__75579\
        );

    \I__18535\ : Span4Mux_h
    port map (
            O => \N__75584\,
            I => \N__75579\
        );

    \I__18534\ : Odrv4
    port map (
            O => \N__75579\,
            I => \c0.n20409\
        );

    \I__18533\ : CascadeMux
    port map (
            O => \N__75576\,
            I => \N__75573\
        );

    \I__18532\ : InMux
    port map (
            O => \N__75573\,
            I => \N__75570\
        );

    \I__18531\ : LocalMux
    port map (
            O => \N__75570\,
            I => \N__75567\
        );

    \I__18530\ : Span4Mux_h
    port map (
            O => \N__75567\,
            I => \N__75563\
        );

    \I__18529\ : InMux
    port map (
            O => \N__75566\,
            I => \N__75559\
        );

    \I__18528\ : Sp12to4
    port map (
            O => \N__75563\,
            I => \N__75555\
        );

    \I__18527\ : CascadeMux
    port map (
            O => \N__75562\,
            I => \N__75550\
        );

    \I__18526\ : LocalMux
    port map (
            O => \N__75559\,
            I => \N__75545\
        );

    \I__18525\ : InMux
    port map (
            O => \N__75558\,
            I => \N__75542\
        );

    \I__18524\ : Span12Mux_v
    port map (
            O => \N__75555\,
            I => \N__75539\
        );

    \I__18523\ : InMux
    port map (
            O => \N__75554\,
            I => \N__75536\
        );

    \I__18522\ : InMux
    port map (
            O => \N__75553\,
            I => \N__75533\
        );

    \I__18521\ : InMux
    port map (
            O => \N__75550\,
            I => \N__75528\
        );

    \I__18520\ : InMux
    port map (
            O => \N__75549\,
            I => \N__75528\
        );

    \I__18519\ : InMux
    port map (
            O => \N__75548\,
            I => \N__75525\
        );

    \I__18518\ : Span4Mux_v
    port map (
            O => \N__75545\,
            I => \N__75522\
        );

    \I__18517\ : LocalMux
    port map (
            O => \N__75542\,
            I => data_in_frame_22_4
        );

    \I__18516\ : Odrv12
    port map (
            O => \N__75539\,
            I => data_in_frame_22_4
        );

    \I__18515\ : LocalMux
    port map (
            O => \N__75536\,
            I => data_in_frame_22_4
        );

    \I__18514\ : LocalMux
    port map (
            O => \N__75533\,
            I => data_in_frame_22_4
        );

    \I__18513\ : LocalMux
    port map (
            O => \N__75528\,
            I => data_in_frame_22_4
        );

    \I__18512\ : LocalMux
    port map (
            O => \N__75525\,
            I => data_in_frame_22_4
        );

    \I__18511\ : Odrv4
    port map (
            O => \N__75522\,
            I => data_in_frame_22_4
        );

    \I__18510\ : InMux
    port map (
            O => \N__75507\,
            I => \N__75501\
        );

    \I__18509\ : InMux
    port map (
            O => \N__75506\,
            I => \N__75501\
        );

    \I__18508\ : LocalMux
    port map (
            O => \N__75501\,
            I => \N__75495\
        );

    \I__18507\ : InMux
    port map (
            O => \N__75500\,
            I => \N__75489\
        );

    \I__18506\ : InMux
    port map (
            O => \N__75499\,
            I => \N__75484\
        );

    \I__18505\ : InMux
    port map (
            O => \N__75498\,
            I => \N__75484\
        );

    \I__18504\ : Span4Mux_h
    port map (
            O => \N__75495\,
            I => \N__75481\
        );

    \I__18503\ : InMux
    port map (
            O => \N__75494\,
            I => \N__75476\
        );

    \I__18502\ : InMux
    port map (
            O => \N__75493\,
            I => \N__75476\
        );

    \I__18501\ : InMux
    port map (
            O => \N__75492\,
            I => \N__75473\
        );

    \I__18500\ : LocalMux
    port map (
            O => \N__75489\,
            I => \N__75470\
        );

    \I__18499\ : LocalMux
    port map (
            O => \N__75484\,
            I => \N__75467\
        );

    \I__18498\ : Span4Mux_v
    port map (
            O => \N__75481\,
            I => \N__75464\
        );

    \I__18497\ : LocalMux
    port map (
            O => \N__75476\,
            I => \N__75461\
        );

    \I__18496\ : LocalMux
    port map (
            O => \N__75473\,
            I => \N__75458\
        );

    \I__18495\ : Span4Mux_h
    port map (
            O => \N__75470\,
            I => \N__75455\
        );

    \I__18494\ : Span4Mux_v
    port map (
            O => \N__75467\,
            I => \N__75452\
        );

    \I__18493\ : Span4Mux_v
    port map (
            O => \N__75464\,
            I => \N__75449\
        );

    \I__18492\ : Span4Mux_h
    port map (
            O => \N__75461\,
            I => \N__75442\
        );

    \I__18491\ : Span4Mux_h
    port map (
            O => \N__75458\,
            I => \N__75442\
        );

    \I__18490\ : Span4Mux_v
    port map (
            O => \N__75455\,
            I => \N__75442\
        );

    \I__18489\ : Span4Mux_v
    port map (
            O => \N__75452\,
            I => \N__75439\
        );

    \I__18488\ : Span4Mux_h
    port map (
            O => \N__75449\,
            I => \N__75436\
        );

    \I__18487\ : Span4Mux_v
    port map (
            O => \N__75442\,
            I => \N__75433\
        );

    \I__18486\ : Odrv4
    port map (
            O => \N__75439\,
            I => \c0.n12_adj_4672\
        );

    \I__18485\ : Odrv4
    port map (
            O => \N__75436\,
            I => \c0.n12_adj_4672\
        );

    \I__18484\ : Odrv4
    port map (
            O => \N__75433\,
            I => \c0.n12_adj_4672\
        );

    \I__18483\ : CascadeMux
    port map (
            O => \N__75426\,
            I => \N__75423\
        );

    \I__18482\ : InMux
    port map (
            O => \N__75423\,
            I => \N__75417\
        );

    \I__18481\ : InMux
    port map (
            O => \N__75422\,
            I => \N__75408\
        );

    \I__18480\ : InMux
    port map (
            O => \N__75421\,
            I => \N__75408\
        );

    \I__18479\ : InMux
    port map (
            O => \N__75420\,
            I => \N__75408\
        );

    \I__18478\ : LocalMux
    port map (
            O => \N__75417\,
            I => \N__75403\
        );

    \I__18477\ : InMux
    port map (
            O => \N__75416\,
            I => \N__75400\
        );

    \I__18476\ : InMux
    port map (
            O => \N__75415\,
            I => \N__75394\
        );

    \I__18475\ : LocalMux
    port map (
            O => \N__75408\,
            I => \N__75390\
        );

    \I__18474\ : InMux
    port map (
            O => \N__75407\,
            I => \N__75385\
        );

    \I__18473\ : InMux
    port map (
            O => \N__75406\,
            I => \N__75385\
        );

    \I__18472\ : Span4Mux_h
    port map (
            O => \N__75403\,
            I => \N__75380\
        );

    \I__18471\ : LocalMux
    port map (
            O => \N__75400\,
            I => \N__75380\
        );

    \I__18470\ : InMux
    port map (
            O => \N__75399\,
            I => \N__75375\
        );

    \I__18469\ : InMux
    port map (
            O => \N__75398\,
            I => \N__75375\
        );

    \I__18468\ : InMux
    port map (
            O => \N__75397\,
            I => \N__75370\
        );

    \I__18467\ : LocalMux
    port map (
            O => \N__75394\,
            I => \N__75367\
        );

    \I__18466\ : InMux
    port map (
            O => \N__75393\,
            I => \N__75364\
        );

    \I__18465\ : Span4Mux_h
    port map (
            O => \N__75390\,
            I => \N__75359\
        );

    \I__18464\ : LocalMux
    port map (
            O => \N__75385\,
            I => \N__75359\
        );

    \I__18463\ : Span4Mux_h
    port map (
            O => \N__75380\,
            I => \N__75356\
        );

    \I__18462\ : LocalMux
    port map (
            O => \N__75375\,
            I => \N__75353\
        );

    \I__18461\ : InMux
    port map (
            O => \N__75374\,
            I => \N__75350\
        );

    \I__18460\ : InMux
    port map (
            O => \N__75373\,
            I => \N__75347\
        );

    \I__18459\ : LocalMux
    port map (
            O => \N__75370\,
            I => \N__75344\
        );

    \I__18458\ : Span4Mux_h
    port map (
            O => \N__75367\,
            I => \N__75341\
        );

    \I__18457\ : LocalMux
    port map (
            O => \N__75364\,
            I => \N__75338\
        );

    \I__18456\ : Span4Mux_v
    port map (
            O => \N__75359\,
            I => \N__75334\
        );

    \I__18455\ : Sp12to4
    port map (
            O => \N__75356\,
            I => \N__75331\
        );

    \I__18454\ : Span4Mux_v
    port map (
            O => \N__75353\,
            I => \N__75328\
        );

    \I__18453\ : LocalMux
    port map (
            O => \N__75350\,
            I => \N__75321\
        );

    \I__18452\ : LocalMux
    port map (
            O => \N__75347\,
            I => \N__75321\
        );

    \I__18451\ : Span4Mux_v
    port map (
            O => \N__75344\,
            I => \N__75318\
        );

    \I__18450\ : Span4Mux_h
    port map (
            O => \N__75341\,
            I => \N__75313\
        );

    \I__18449\ : Span4Mux_v
    port map (
            O => \N__75338\,
            I => \N__75313\
        );

    \I__18448\ : InMux
    port map (
            O => \N__75337\,
            I => \N__75310\
        );

    \I__18447\ : Sp12to4
    port map (
            O => \N__75334\,
            I => \N__75307\
        );

    \I__18446\ : Span12Mux_v
    port map (
            O => \N__75331\,
            I => \N__75302\
        );

    \I__18445\ : Sp12to4
    port map (
            O => \N__75328\,
            I => \N__75302\
        );

    \I__18444\ : InMux
    port map (
            O => \N__75327\,
            I => \N__75298\
        );

    \I__18443\ : InMux
    port map (
            O => \N__75326\,
            I => \N__75295\
        );

    \I__18442\ : Span4Mux_h
    port map (
            O => \N__75321\,
            I => \N__75290\
        );

    \I__18441\ : Span4Mux_v
    port map (
            O => \N__75318\,
            I => \N__75290\
        );

    \I__18440\ : Span4Mux_v
    port map (
            O => \N__75313\,
            I => \N__75287\
        );

    \I__18439\ : LocalMux
    port map (
            O => \N__75310\,
            I => \N__75280\
        );

    \I__18438\ : Span12Mux_h
    port map (
            O => \N__75307\,
            I => \N__75280\
        );

    \I__18437\ : Span12Mux_h
    port map (
            O => \N__75302\,
            I => \N__75280\
        );

    \I__18436\ : InMux
    port map (
            O => \N__75301\,
            I => \N__75277\
        );

    \I__18435\ : LocalMux
    port map (
            O => \N__75298\,
            I => \N__75274\
        );

    \I__18434\ : LocalMux
    port map (
            O => \N__75295\,
            I => \c0.n22099\
        );

    \I__18433\ : Odrv4
    port map (
            O => \N__75290\,
            I => \c0.n22099\
        );

    \I__18432\ : Odrv4
    port map (
            O => \N__75287\,
            I => \c0.n22099\
        );

    \I__18431\ : Odrv12
    port map (
            O => \N__75280\,
            I => \c0.n22099\
        );

    \I__18430\ : LocalMux
    port map (
            O => \N__75277\,
            I => \c0.n22099\
        );

    \I__18429\ : Odrv12
    port map (
            O => \N__75274\,
            I => \c0.n22099\
        );

    \I__18428\ : InMux
    port map (
            O => \N__75261\,
            I => \N__75258\
        );

    \I__18427\ : LocalMux
    port map (
            O => \N__75258\,
            I => \N__75245\
        );

    \I__18426\ : InMux
    port map (
            O => \N__75257\,
            I => \N__75239\
        );

    \I__18425\ : InMux
    port map (
            O => \N__75256\,
            I => \N__75236\
        );

    \I__18424\ : InMux
    port map (
            O => \N__75255\,
            I => \N__75233\
        );

    \I__18423\ : CascadeMux
    port map (
            O => \N__75254\,
            I => \N__75230\
        );

    \I__18422\ : InMux
    port map (
            O => \N__75253\,
            I => \N__75225\
        );

    \I__18421\ : InMux
    port map (
            O => \N__75252\,
            I => \N__75219\
        );

    \I__18420\ : InMux
    port map (
            O => \N__75251\,
            I => \N__75219\
        );

    \I__18419\ : InMux
    port map (
            O => \N__75250\,
            I => \N__75216\
        );

    \I__18418\ : InMux
    port map (
            O => \N__75249\,
            I => \N__75211\
        );

    \I__18417\ : InMux
    port map (
            O => \N__75248\,
            I => \N__75211\
        );

    \I__18416\ : Span4Mux_v
    port map (
            O => \N__75245\,
            I => \N__75208\
        );

    \I__18415\ : InMux
    port map (
            O => \N__75244\,
            I => \N__75205\
        );

    \I__18414\ : InMux
    port map (
            O => \N__75243\,
            I => \N__75202\
        );

    \I__18413\ : InMux
    port map (
            O => \N__75242\,
            I => \N__75199\
        );

    \I__18412\ : LocalMux
    port map (
            O => \N__75239\,
            I => \N__75196\
        );

    \I__18411\ : LocalMux
    port map (
            O => \N__75236\,
            I => \N__75190\
        );

    \I__18410\ : LocalMux
    port map (
            O => \N__75233\,
            I => \N__75190\
        );

    \I__18409\ : InMux
    port map (
            O => \N__75230\,
            I => \N__75187\
        );

    \I__18408\ : CascadeMux
    port map (
            O => \N__75229\,
            I => \N__75182\
        );

    \I__18407\ : CascadeMux
    port map (
            O => \N__75228\,
            I => \N__75179\
        );

    \I__18406\ : LocalMux
    port map (
            O => \N__75225\,
            I => \N__75174\
        );

    \I__18405\ : InMux
    port map (
            O => \N__75224\,
            I => \N__75171\
        );

    \I__18404\ : LocalMux
    port map (
            O => \N__75219\,
            I => \N__75166\
        );

    \I__18403\ : LocalMux
    port map (
            O => \N__75216\,
            I => \N__75166\
        );

    \I__18402\ : LocalMux
    port map (
            O => \N__75211\,
            I => \N__75163\
        );

    \I__18401\ : Span4Mux_h
    port map (
            O => \N__75208\,
            I => \N__75160\
        );

    \I__18400\ : LocalMux
    port map (
            O => \N__75205\,
            I => \N__75153\
        );

    \I__18399\ : LocalMux
    port map (
            O => \N__75202\,
            I => \N__75153\
        );

    \I__18398\ : LocalMux
    port map (
            O => \N__75199\,
            I => \N__75153\
        );

    \I__18397\ : Span4Mux_h
    port map (
            O => \N__75196\,
            I => \N__75150\
        );

    \I__18396\ : InMux
    port map (
            O => \N__75195\,
            I => \N__75147\
        );

    \I__18395\ : Span4Mux_v
    port map (
            O => \N__75190\,
            I => \N__75142\
        );

    \I__18394\ : LocalMux
    port map (
            O => \N__75187\,
            I => \N__75142\
        );

    \I__18393\ : InMux
    port map (
            O => \N__75186\,
            I => \N__75139\
        );

    \I__18392\ : InMux
    port map (
            O => \N__75185\,
            I => \N__75134\
        );

    \I__18391\ : InMux
    port map (
            O => \N__75182\,
            I => \N__75131\
        );

    \I__18390\ : InMux
    port map (
            O => \N__75179\,
            I => \N__75128\
        );

    \I__18389\ : InMux
    port map (
            O => \N__75178\,
            I => \N__75125\
        );

    \I__18388\ : InMux
    port map (
            O => \N__75177\,
            I => \N__75122\
        );

    \I__18387\ : Span4Mux_v
    port map (
            O => \N__75174\,
            I => \N__75117\
        );

    \I__18386\ : LocalMux
    port map (
            O => \N__75171\,
            I => \N__75117\
        );

    \I__18385\ : Span4Mux_h
    port map (
            O => \N__75166\,
            I => \N__75114\
        );

    \I__18384\ : Span4Mux_v
    port map (
            O => \N__75163\,
            I => \N__75103\
        );

    \I__18383\ : Span4Mux_h
    port map (
            O => \N__75160\,
            I => \N__75103\
        );

    \I__18382\ : Span4Mux_v
    port map (
            O => \N__75153\,
            I => \N__75103\
        );

    \I__18381\ : Span4Mux_h
    port map (
            O => \N__75150\,
            I => \N__75098\
        );

    \I__18380\ : LocalMux
    port map (
            O => \N__75147\,
            I => \N__75098\
        );

    \I__18379\ : Span4Mux_v
    port map (
            O => \N__75142\,
            I => \N__75093\
        );

    \I__18378\ : LocalMux
    port map (
            O => \N__75139\,
            I => \N__75093\
        );

    \I__18377\ : InMux
    port map (
            O => \N__75138\,
            I => \N__75088\
        );

    \I__18376\ : InMux
    port map (
            O => \N__75137\,
            I => \N__75088\
        );

    \I__18375\ : LocalMux
    port map (
            O => \N__75134\,
            I => \N__75085\
        );

    \I__18374\ : LocalMux
    port map (
            O => \N__75131\,
            I => \N__75080\
        );

    \I__18373\ : LocalMux
    port map (
            O => \N__75128\,
            I => \N__75080\
        );

    \I__18372\ : LocalMux
    port map (
            O => \N__75125\,
            I => \N__75077\
        );

    \I__18371\ : LocalMux
    port map (
            O => \N__75122\,
            I => \N__75074\
        );

    \I__18370\ : Span4Mux_v
    port map (
            O => \N__75117\,
            I => \N__75071\
        );

    \I__18369\ : Span4Mux_v
    port map (
            O => \N__75114\,
            I => \N__75068\
        );

    \I__18368\ : InMux
    port map (
            O => \N__75113\,
            I => \N__75065\
        );

    \I__18367\ : InMux
    port map (
            O => \N__75112\,
            I => \N__75062\
        );

    \I__18366\ : InMux
    port map (
            O => \N__75111\,
            I => \N__75057\
        );

    \I__18365\ : InMux
    port map (
            O => \N__75110\,
            I => \N__75057\
        );

    \I__18364\ : Sp12to4
    port map (
            O => \N__75103\,
            I => \N__75054\
        );

    \I__18363\ : Span4Mux_h
    port map (
            O => \N__75098\,
            I => \N__75051\
        );

    \I__18362\ : Span4Mux_h
    port map (
            O => \N__75093\,
            I => \N__75048\
        );

    \I__18361\ : LocalMux
    port map (
            O => \N__75088\,
            I => \N__75041\
        );

    \I__18360\ : Span4Mux_h
    port map (
            O => \N__75085\,
            I => \N__75041\
        );

    \I__18359\ : Span4Mux_v
    port map (
            O => \N__75080\,
            I => \N__75034\
        );

    \I__18358\ : Span4Mux_v
    port map (
            O => \N__75077\,
            I => \N__75034\
        );

    \I__18357\ : Span4Mux_v
    port map (
            O => \N__75074\,
            I => \N__75034\
        );

    \I__18356\ : Span4Mux_h
    port map (
            O => \N__75071\,
            I => \N__75029\
        );

    \I__18355\ : Span4Mux_v
    port map (
            O => \N__75068\,
            I => \N__75029\
        );

    \I__18354\ : LocalMux
    port map (
            O => \N__75065\,
            I => \N__75022\
        );

    \I__18353\ : LocalMux
    port map (
            O => \N__75062\,
            I => \N__75022\
        );

    \I__18352\ : LocalMux
    port map (
            O => \N__75057\,
            I => \N__75019\
        );

    \I__18351\ : Span12Mux_h
    port map (
            O => \N__75054\,
            I => \N__75012\
        );

    \I__18350\ : Sp12to4
    port map (
            O => \N__75051\,
            I => \N__75012\
        );

    \I__18349\ : Sp12to4
    port map (
            O => \N__75048\,
            I => \N__75012\
        );

    \I__18348\ : InMux
    port map (
            O => \N__75047\,
            I => \N__75007\
        );

    \I__18347\ : InMux
    port map (
            O => \N__75046\,
            I => \N__75007\
        );

    \I__18346\ : Span4Mux_v
    port map (
            O => \N__75041\,
            I => \N__75002\
        );

    \I__18345\ : Span4Mux_h
    port map (
            O => \N__75034\,
            I => \N__75002\
        );

    \I__18344\ : Sp12to4
    port map (
            O => \N__75029\,
            I => \N__74999\
        );

    \I__18343\ : InMux
    port map (
            O => \N__75028\,
            I => \N__74996\
        );

    \I__18342\ : InMux
    port map (
            O => \N__75027\,
            I => \N__74993\
        );

    \I__18341\ : Span4Mux_v
    port map (
            O => \N__75022\,
            I => \N__74990\
        );

    \I__18340\ : Span4Mux_h
    port map (
            O => \N__75019\,
            I => \N__74987\
        );

    \I__18339\ : Span12Mux_v
    port map (
            O => \N__75012\,
            I => \N__74984\
        );

    \I__18338\ : LocalMux
    port map (
            O => \N__75007\,
            I => \N__74977\
        );

    \I__18337\ : Sp12to4
    port map (
            O => \N__75002\,
            I => \N__74977\
        );

    \I__18336\ : Span12Mux_s6_h
    port map (
            O => \N__74999\,
            I => \N__74977\
        );

    \I__18335\ : LocalMux
    port map (
            O => \N__74996\,
            I => rx_data_1
        );

    \I__18334\ : LocalMux
    port map (
            O => \N__74993\,
            I => rx_data_1
        );

    \I__18333\ : Odrv4
    port map (
            O => \N__74990\,
            I => rx_data_1
        );

    \I__18332\ : Odrv4
    port map (
            O => \N__74987\,
            I => rx_data_1
        );

    \I__18331\ : Odrv12
    port map (
            O => \N__74984\,
            I => rx_data_1
        );

    \I__18330\ : Odrv12
    port map (
            O => \N__74977\,
            I => rx_data_1
        );

    \I__18329\ : CascadeMux
    port map (
            O => \N__74964\,
            I => \N__74958\
        );

    \I__18328\ : CascadeMux
    port map (
            O => \N__74963\,
            I => \N__74955\
        );

    \I__18327\ : InMux
    port map (
            O => \N__74962\,
            I => \N__74952\
        );

    \I__18326\ : InMux
    port map (
            O => \N__74961\,
            I => \N__74949\
        );

    \I__18325\ : InMux
    port map (
            O => \N__74958\,
            I => \N__74946\
        );

    \I__18324\ : InMux
    port map (
            O => \N__74955\,
            I => \N__74943\
        );

    \I__18323\ : LocalMux
    port map (
            O => \N__74952\,
            I => \N__74940\
        );

    \I__18322\ : LocalMux
    port map (
            O => \N__74949\,
            I => \N__74937\
        );

    \I__18321\ : LocalMux
    port map (
            O => \N__74946\,
            I => \N__74934\
        );

    \I__18320\ : LocalMux
    port map (
            O => \N__74943\,
            I => \N__74930\
        );

    \I__18319\ : Span4Mux_h
    port map (
            O => \N__74940\,
            I => \N__74927\
        );

    \I__18318\ : Span4Mux_v
    port map (
            O => \N__74937\,
            I => \N__74922\
        );

    \I__18317\ : Span4Mux_v
    port map (
            O => \N__74934\,
            I => \N__74922\
        );

    \I__18316\ : InMux
    port map (
            O => \N__74933\,
            I => \N__74919\
        );

    \I__18315\ : Span4Mux_h
    port map (
            O => \N__74930\,
            I => \N__74914\
        );

    \I__18314\ : Span4Mux_v
    port map (
            O => \N__74927\,
            I => \N__74914\
        );

    \I__18313\ : Span4Mux_h
    port map (
            O => \N__74922\,
            I => \N__74911\
        );

    \I__18312\ : LocalMux
    port map (
            O => \N__74919\,
            I => \c0.data_in_frame_13_1\
        );

    \I__18311\ : Odrv4
    port map (
            O => \N__74914\,
            I => \c0.data_in_frame_13_1\
        );

    \I__18310\ : Odrv4
    port map (
            O => \N__74911\,
            I => \c0.data_in_frame_13_1\
        );

    \I__18309\ : InMux
    port map (
            O => \N__74904\,
            I => \N__74900\
        );

    \I__18308\ : InMux
    port map (
            O => \N__74903\,
            I => \N__74897\
        );

    \I__18307\ : LocalMux
    port map (
            O => \N__74900\,
            I => \N__74894\
        );

    \I__18306\ : LocalMux
    port map (
            O => \N__74897\,
            I => \N__74890\
        );

    \I__18305\ : Span4Mux_v
    port map (
            O => \N__74894\,
            I => \N__74887\
        );

    \I__18304\ : InMux
    port map (
            O => \N__74893\,
            I => \N__74884\
        );

    \I__18303\ : Span4Mux_h
    port map (
            O => \N__74890\,
            I => \N__74881\
        );

    \I__18302\ : Odrv4
    port map (
            O => \N__74887\,
            I => \c0.n13490\
        );

    \I__18301\ : LocalMux
    port map (
            O => \N__74884\,
            I => \c0.n13490\
        );

    \I__18300\ : Odrv4
    port map (
            O => \N__74881\,
            I => \c0.n13490\
        );

    \I__18299\ : InMux
    port map (
            O => \N__74874\,
            I => \N__74871\
        );

    \I__18298\ : LocalMux
    port map (
            O => \N__74871\,
            I => \N__74867\
        );

    \I__18297\ : CascadeMux
    port map (
            O => \N__74870\,
            I => \N__74863\
        );

    \I__18296\ : Span4Mux_h
    port map (
            O => \N__74867\,
            I => \N__74860\
        );

    \I__18295\ : CascadeMux
    port map (
            O => \N__74866\,
            I => \N__74857\
        );

    \I__18294\ : InMux
    port map (
            O => \N__74863\,
            I => \N__74854\
        );

    \I__18293\ : Span4Mux_h
    port map (
            O => \N__74860\,
            I => \N__74851\
        );

    \I__18292\ : InMux
    port map (
            O => \N__74857\,
            I => \N__74848\
        );

    \I__18291\ : LocalMux
    port map (
            O => \N__74854\,
            I => \c0.data_in_frame_24_5\
        );

    \I__18290\ : Odrv4
    port map (
            O => \N__74851\,
            I => \c0.data_in_frame_24_5\
        );

    \I__18289\ : LocalMux
    port map (
            O => \N__74848\,
            I => \c0.data_in_frame_24_5\
        );

    \I__18288\ : InMux
    port map (
            O => \N__74841\,
            I => \N__74838\
        );

    \I__18287\ : LocalMux
    port map (
            O => \N__74838\,
            I => \N__74834\
        );

    \I__18286\ : InMux
    port map (
            O => \N__74837\,
            I => \N__74831\
        );

    \I__18285\ : Span4Mux_h
    port map (
            O => \N__74834\,
            I => \N__74828\
        );

    \I__18284\ : LocalMux
    port map (
            O => \N__74831\,
            I => \N__74825\
        );

    \I__18283\ : Span4Mux_h
    port map (
            O => \N__74828\,
            I => \N__74822\
        );

    \I__18282\ : Odrv4
    port map (
            O => \N__74825\,
            I => \c0.n22505\
        );

    \I__18281\ : Odrv4
    port map (
            O => \N__74822\,
            I => \c0.n22505\
        );

    \I__18280\ : InMux
    port map (
            O => \N__74817\,
            I => \N__74812\
        );

    \I__18279\ : InMux
    port map (
            O => \N__74816\,
            I => \N__74808\
        );

    \I__18278\ : InMux
    port map (
            O => \N__74815\,
            I => \N__74805\
        );

    \I__18277\ : LocalMux
    port map (
            O => \N__74812\,
            I => \N__74802\
        );

    \I__18276\ : InMux
    port map (
            O => \N__74811\,
            I => \N__74799\
        );

    \I__18275\ : LocalMux
    port map (
            O => \N__74808\,
            I => \N__74794\
        );

    \I__18274\ : LocalMux
    port map (
            O => \N__74805\,
            I => \N__74794\
        );

    \I__18273\ : Span4Mux_v
    port map (
            O => \N__74802\,
            I => \N__74789\
        );

    \I__18272\ : LocalMux
    port map (
            O => \N__74799\,
            I => \N__74789\
        );

    \I__18271\ : Span4Mux_v
    port map (
            O => \N__74794\,
            I => \N__74786\
        );

    \I__18270\ : Span4Mux_h
    port map (
            O => \N__74789\,
            I => \N__74783\
        );

    \I__18269\ : Odrv4
    port map (
            O => \N__74786\,
            I => \c0.n6718\
        );

    \I__18268\ : Odrv4
    port map (
            O => \N__74783\,
            I => \c0.n6718\
        );

    \I__18267\ : InMux
    port map (
            O => \N__74778\,
            I => \N__74775\
        );

    \I__18266\ : LocalMux
    port map (
            O => \N__74775\,
            I => \N__74769\
        );

    \I__18265\ : CascadeMux
    port map (
            O => \N__74774\,
            I => \N__74765\
        );

    \I__18264\ : InMux
    port map (
            O => \N__74773\,
            I => \N__74760\
        );

    \I__18263\ : InMux
    port map (
            O => \N__74772\,
            I => \N__74760\
        );

    \I__18262\ : Span4Mux_h
    port map (
            O => \N__74769\,
            I => \N__74757\
        );

    \I__18261\ : InMux
    port map (
            O => \N__74768\,
            I => \N__74752\
        );

    \I__18260\ : InMux
    port map (
            O => \N__74765\,
            I => \N__74752\
        );

    \I__18259\ : LocalMux
    port map (
            O => \N__74760\,
            I => \c0.n13963\
        );

    \I__18258\ : Odrv4
    port map (
            O => \N__74757\,
            I => \c0.n13963\
        );

    \I__18257\ : LocalMux
    port map (
            O => \N__74752\,
            I => \c0.n13963\
        );

    \I__18256\ : InMux
    port map (
            O => \N__74745\,
            I => \N__74742\
        );

    \I__18255\ : LocalMux
    port map (
            O => \N__74742\,
            I => \N__74739\
        );

    \I__18254\ : Span4Mux_v
    port map (
            O => \N__74739\,
            I => \N__74736\
        );

    \I__18253\ : Odrv4
    port map (
            O => \N__74736\,
            I => \c0.n21295\
        );

    \I__18252\ : InMux
    port map (
            O => \N__74733\,
            I => \N__74730\
        );

    \I__18251\ : LocalMux
    port map (
            O => \N__74730\,
            I => \N__74727\
        );

    \I__18250\ : Span4Mux_h
    port map (
            O => \N__74727\,
            I => \N__74724\
        );

    \I__18249\ : Span4Mux_h
    port map (
            O => \N__74724\,
            I => \N__74721\
        );

    \I__18248\ : Odrv4
    port map (
            O => \N__74721\,
            I => \c0.n20239\
        );

    \I__18247\ : CascadeMux
    port map (
            O => \N__74718\,
            I => \N__74715\
        );

    \I__18246\ : InMux
    port map (
            O => \N__74715\,
            I => \N__74709\
        );

    \I__18245\ : InMux
    port map (
            O => \N__74714\,
            I => \N__74704\
        );

    \I__18244\ : InMux
    port map (
            O => \N__74713\,
            I => \N__74704\
        );

    \I__18243\ : CascadeMux
    port map (
            O => \N__74712\,
            I => \N__74701\
        );

    \I__18242\ : LocalMux
    port map (
            O => \N__74709\,
            I => \N__74698\
        );

    \I__18241\ : LocalMux
    port map (
            O => \N__74704\,
            I => \N__74695\
        );

    \I__18240\ : InMux
    port map (
            O => \N__74701\,
            I => \N__74692\
        );

    \I__18239\ : Span12Mux_h
    port map (
            O => \N__74698\,
            I => \N__74689\
        );

    \I__18238\ : Span4Mux_h
    port map (
            O => \N__74695\,
            I => \N__74686\
        );

    \I__18237\ : LocalMux
    port map (
            O => \N__74692\,
            I => \c0.data_in_frame_17_1\
        );

    \I__18236\ : Odrv12
    port map (
            O => \N__74689\,
            I => \c0.data_in_frame_17_1\
        );

    \I__18235\ : Odrv4
    port map (
            O => \N__74686\,
            I => \c0.data_in_frame_17_1\
        );

    \I__18234\ : InMux
    port map (
            O => \N__74679\,
            I => \N__74675\
        );

    \I__18233\ : InMux
    port map (
            O => \N__74678\,
            I => \N__74670\
        );

    \I__18232\ : LocalMux
    port map (
            O => \N__74675\,
            I => \N__74667\
        );

    \I__18231\ : CascadeMux
    port map (
            O => \N__74674\,
            I => \N__74663\
        );

    \I__18230\ : InMux
    port map (
            O => \N__74673\,
            I => \N__74660\
        );

    \I__18229\ : LocalMux
    port map (
            O => \N__74670\,
            I => \N__74655\
        );

    \I__18228\ : Span4Mux_v
    port map (
            O => \N__74667\,
            I => \N__74652\
        );

    \I__18227\ : InMux
    port map (
            O => \N__74666\,
            I => \N__74647\
        );

    \I__18226\ : InMux
    port map (
            O => \N__74663\,
            I => \N__74647\
        );

    \I__18225\ : LocalMux
    port map (
            O => \N__74660\,
            I => \N__74644\
        );

    \I__18224\ : InMux
    port map (
            O => \N__74659\,
            I => \N__74637\
        );

    \I__18223\ : InMux
    port map (
            O => \N__74658\,
            I => \N__74637\
        );

    \I__18222\ : Span4Mux_h
    port map (
            O => \N__74655\,
            I => \N__74633\
        );

    \I__18221\ : Sp12to4
    port map (
            O => \N__74652\,
            I => \N__74626\
        );

    \I__18220\ : LocalMux
    port map (
            O => \N__74647\,
            I => \N__74626\
        );

    \I__18219\ : Span4Mux_h
    port map (
            O => \N__74644\,
            I => \N__74622\
        );

    \I__18218\ : InMux
    port map (
            O => \N__74643\,
            I => \N__74619\
        );

    \I__18217\ : InMux
    port map (
            O => \N__74642\,
            I => \N__74616\
        );

    \I__18216\ : LocalMux
    port map (
            O => \N__74637\,
            I => \N__74613\
        );

    \I__18215\ : InMux
    port map (
            O => \N__74636\,
            I => \N__74610\
        );

    \I__18214\ : Sp12to4
    port map (
            O => \N__74633\,
            I => \N__74607\
        );

    \I__18213\ : InMux
    port map (
            O => \N__74632\,
            I => \N__74604\
        );

    \I__18212\ : InMux
    port map (
            O => \N__74631\,
            I => \N__74601\
        );

    \I__18211\ : Span12Mux_h
    port map (
            O => \N__74626\,
            I => \N__74598\
        );

    \I__18210\ : InMux
    port map (
            O => \N__74625\,
            I => \N__74595\
        );

    \I__18209\ : Span4Mux_v
    port map (
            O => \N__74622\,
            I => \N__74592\
        );

    \I__18208\ : LocalMux
    port map (
            O => \N__74619\,
            I => \N__74589\
        );

    \I__18207\ : LocalMux
    port map (
            O => \N__74616\,
            I => \N__74586\
        );

    \I__18206\ : Span4Mux_v
    port map (
            O => \N__74613\,
            I => \N__74581\
        );

    \I__18205\ : LocalMux
    port map (
            O => \N__74610\,
            I => \N__74581\
        );

    \I__18204\ : Span12Mux_v
    port map (
            O => \N__74607\,
            I => \N__74578\
        );

    \I__18203\ : LocalMux
    port map (
            O => \N__74604\,
            I => \N__74573\
        );

    \I__18202\ : LocalMux
    port map (
            O => \N__74601\,
            I => \N__74573\
        );

    \I__18201\ : Span12Mux_v
    port map (
            O => \N__74598\,
            I => \N__74570\
        );

    \I__18200\ : LocalMux
    port map (
            O => \N__74595\,
            I => \N__74563\
        );

    \I__18199\ : Span4Mux_v
    port map (
            O => \N__74592\,
            I => \N__74563\
        );

    \I__18198\ : Span4Mux_h
    port map (
            O => \N__74589\,
            I => \N__74563\
        );

    \I__18197\ : Span4Mux_v
    port map (
            O => \N__74586\,
            I => \N__74559\
        );

    \I__18196\ : Span4Mux_v
    port map (
            O => \N__74581\,
            I => \N__74556\
        );

    \I__18195\ : Span12Mux_v
    port map (
            O => \N__74578\,
            I => \N__74553\
        );

    \I__18194\ : Span12Mux_h
    port map (
            O => \N__74573\,
            I => \N__74548\
        );

    \I__18193\ : Span12Mux_h
    port map (
            O => \N__74570\,
            I => \N__74548\
        );

    \I__18192\ : Span4Mux_v
    port map (
            O => \N__74563\,
            I => \N__74545\
        );

    \I__18191\ : InMux
    port map (
            O => \N__74562\,
            I => \N__74542\
        );

    \I__18190\ : Odrv4
    port map (
            O => \N__74559\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__18189\ : Odrv4
    port map (
            O => \N__74556\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__18188\ : Odrv12
    port map (
            O => \N__74553\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__18187\ : Odrv12
    port map (
            O => \N__74548\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__18186\ : Odrv4
    port map (
            O => \N__74545\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__18185\ : LocalMux
    port map (
            O => \N__74542\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__18184\ : InMux
    port map (
            O => \N__74529\,
            I => \N__74526\
        );

    \I__18183\ : LocalMux
    port map (
            O => \N__74526\,
            I => \N__74521\
        );

    \I__18182\ : InMux
    port map (
            O => \N__74525\,
            I => \N__74517\
        );

    \I__18181\ : InMux
    port map (
            O => \N__74524\,
            I => \N__74514\
        );

    \I__18180\ : Span4Mux_v
    port map (
            O => \N__74521\,
            I => \N__74511\
        );

    \I__18179\ : InMux
    port map (
            O => \N__74520\,
            I => \N__74508\
        );

    \I__18178\ : LocalMux
    port map (
            O => \N__74517\,
            I => \N__74504\
        );

    \I__18177\ : LocalMux
    port map (
            O => \N__74514\,
            I => \N__74501\
        );

    \I__18176\ : Span4Mux_h
    port map (
            O => \N__74511\,
            I => \N__74493\
        );

    \I__18175\ : LocalMux
    port map (
            O => \N__74508\,
            I => \N__74493\
        );

    \I__18174\ : InMux
    port map (
            O => \N__74507\,
            I => \N__74490\
        );

    \I__18173\ : Span4Mux_v
    port map (
            O => \N__74504\,
            I => \N__74487\
        );

    \I__18172\ : Span4Mux_v
    port map (
            O => \N__74501\,
            I => \N__74484\
        );

    \I__18171\ : InMux
    port map (
            O => \N__74500\,
            I => \N__74481\
        );

    \I__18170\ : InMux
    port map (
            O => \N__74499\,
            I => \N__74477\
        );

    \I__18169\ : InMux
    port map (
            O => \N__74498\,
            I => \N__74474\
        );

    \I__18168\ : Span4Mux_v
    port map (
            O => \N__74493\,
            I => \N__74471\
        );

    \I__18167\ : LocalMux
    port map (
            O => \N__74490\,
            I => \N__74466\
        );

    \I__18166\ : Span4Mux_h
    port map (
            O => \N__74487\,
            I => \N__74459\
        );

    \I__18165\ : Span4Mux_v
    port map (
            O => \N__74484\,
            I => \N__74459\
        );

    \I__18164\ : LocalMux
    port map (
            O => \N__74481\,
            I => \N__74459\
        );

    \I__18163\ : InMux
    port map (
            O => \N__74480\,
            I => \N__74456\
        );

    \I__18162\ : LocalMux
    port map (
            O => \N__74477\,
            I => \N__74453\
        );

    \I__18161\ : LocalMux
    port map (
            O => \N__74474\,
            I => \N__74448\
        );

    \I__18160\ : Span4Mux_v
    port map (
            O => \N__74471\,
            I => \N__74448\
        );

    \I__18159\ : InMux
    port map (
            O => \N__74470\,
            I => \N__74442\
        );

    \I__18158\ : InMux
    port map (
            O => \N__74469\,
            I => \N__74442\
        );

    \I__18157\ : Span4Mux_v
    port map (
            O => \N__74466\,
            I => \N__74436\
        );

    \I__18156\ : Span4Mux_v
    port map (
            O => \N__74459\,
            I => \N__74436\
        );

    \I__18155\ : LocalMux
    port map (
            O => \N__74456\,
            I => \N__74429\
        );

    \I__18154\ : Span4Mux_h
    port map (
            O => \N__74453\,
            I => \N__74429\
        );

    \I__18153\ : Span4Mux_v
    port map (
            O => \N__74448\,
            I => \N__74429\
        );

    \I__18152\ : InMux
    port map (
            O => \N__74447\,
            I => \N__74426\
        );

    \I__18151\ : LocalMux
    port map (
            O => \N__74442\,
            I => \N__74423\
        );

    \I__18150\ : InMux
    port map (
            O => \N__74441\,
            I => \N__74420\
        );

    \I__18149\ : Span4Mux_h
    port map (
            O => \N__74436\,
            I => \N__74417\
        );

    \I__18148\ : Span4Mux_v
    port map (
            O => \N__74429\,
            I => \N__74414\
        );

    \I__18147\ : LocalMux
    port map (
            O => \N__74426\,
            I => \N__74407\
        );

    \I__18146\ : Span12Mux_v
    port map (
            O => \N__74423\,
            I => \N__74407\
        );

    \I__18145\ : LocalMux
    port map (
            O => \N__74420\,
            I => \N__74407\
        );

    \I__18144\ : Span4Mux_v
    port map (
            O => \N__74417\,
            I => \N__74403\
        );

    \I__18143\ : Sp12to4
    port map (
            O => \N__74414\,
            I => \N__74398\
        );

    \I__18142\ : Span12Mux_v
    port map (
            O => \N__74407\,
            I => \N__74398\
        );

    \I__18141\ : InMux
    port map (
            O => \N__74406\,
            I => \N__74395\
        );

    \I__18140\ : Odrv4
    port map (
            O => \N__74403\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__18139\ : Odrv12
    port map (
            O => \N__74398\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__18138\ : LocalMux
    port map (
            O => \N__74395\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__18137\ : CascadeMux
    port map (
            O => \N__74388\,
            I => \N__74383\
        );

    \I__18136\ : CascadeMux
    port map (
            O => \N__74387\,
            I => \N__74378\
        );

    \I__18135\ : CascadeMux
    port map (
            O => \N__74386\,
            I => \N__74375\
        );

    \I__18134\ : InMux
    port map (
            O => \N__74383\,
            I => \N__74372\
        );

    \I__18133\ : InMux
    port map (
            O => \N__74382\,
            I => \N__74369\
        );

    \I__18132\ : CascadeMux
    port map (
            O => \N__74381\,
            I => \N__74366\
        );

    \I__18131\ : InMux
    port map (
            O => \N__74378\,
            I => \N__74362\
        );

    \I__18130\ : InMux
    port map (
            O => \N__74375\,
            I => \N__74359\
        );

    \I__18129\ : LocalMux
    port map (
            O => \N__74372\,
            I => \N__74355\
        );

    \I__18128\ : LocalMux
    port map (
            O => \N__74369\,
            I => \N__74352\
        );

    \I__18127\ : InMux
    port map (
            O => \N__74366\,
            I => \N__74349\
        );

    \I__18126\ : InMux
    port map (
            O => \N__74365\,
            I => \N__74345\
        );

    \I__18125\ : LocalMux
    port map (
            O => \N__74362\,
            I => \N__74341\
        );

    \I__18124\ : LocalMux
    port map (
            O => \N__74359\,
            I => \N__74338\
        );

    \I__18123\ : InMux
    port map (
            O => \N__74358\,
            I => \N__74335\
        );

    \I__18122\ : Span4Mux_h
    port map (
            O => \N__74355\,
            I => \N__74332\
        );

    \I__18121\ : Span4Mux_v
    port map (
            O => \N__74352\,
            I => \N__74329\
        );

    \I__18120\ : LocalMux
    port map (
            O => \N__74349\,
            I => \N__74326\
        );

    \I__18119\ : InMux
    port map (
            O => \N__74348\,
            I => \N__74323\
        );

    \I__18118\ : LocalMux
    port map (
            O => \N__74345\,
            I => \N__74320\
        );

    \I__18117\ : InMux
    port map (
            O => \N__74344\,
            I => \N__74317\
        );

    \I__18116\ : Span4Mux_v
    port map (
            O => \N__74341\,
            I => \N__74312\
        );

    \I__18115\ : Span4Mux_h
    port map (
            O => \N__74338\,
            I => \N__74312\
        );

    \I__18114\ : LocalMux
    port map (
            O => \N__74335\,
            I => \N__74309\
        );

    \I__18113\ : Span4Mux_h
    port map (
            O => \N__74332\,
            I => \N__74306\
        );

    \I__18112\ : Span4Mux_v
    port map (
            O => \N__74329\,
            I => \N__74303\
        );

    \I__18111\ : Span4Mux_v
    port map (
            O => \N__74326\,
            I => \N__74297\
        );

    \I__18110\ : LocalMux
    port map (
            O => \N__74323\,
            I => \N__74297\
        );

    \I__18109\ : Span4Mux_v
    port map (
            O => \N__74320\,
            I => \N__74292\
        );

    \I__18108\ : LocalMux
    port map (
            O => \N__74317\,
            I => \N__74292\
        );

    \I__18107\ : Span4Mux_v
    port map (
            O => \N__74312\,
            I => \N__74289\
        );

    \I__18106\ : Span4Mux_h
    port map (
            O => \N__74309\,
            I => \N__74285\
        );

    \I__18105\ : Span4Mux_v
    port map (
            O => \N__74306\,
            I => \N__74280\
        );

    \I__18104\ : Span4Mux_h
    port map (
            O => \N__74303\,
            I => \N__74280\
        );

    \I__18103\ : InMux
    port map (
            O => \N__74302\,
            I => \N__74276\
        );

    \I__18102\ : Span4Mux_v
    port map (
            O => \N__74297\,
            I => \N__74273\
        );

    \I__18101\ : Span4Mux_v
    port map (
            O => \N__74292\,
            I => \N__74270\
        );

    \I__18100\ : Span4Mux_v
    port map (
            O => \N__74289\,
            I => \N__74267\
        );

    \I__18099\ : InMux
    port map (
            O => \N__74288\,
            I => \N__74264\
        );

    \I__18098\ : Span4Mux_h
    port map (
            O => \N__74285\,
            I => \N__74259\
        );

    \I__18097\ : Span4Mux_v
    port map (
            O => \N__74280\,
            I => \N__74259\
        );

    \I__18096\ : InMux
    port map (
            O => \N__74279\,
            I => \N__74256\
        );

    \I__18095\ : LocalMux
    port map (
            O => \N__74276\,
            I => \N__74247\
        );

    \I__18094\ : Span4Mux_h
    port map (
            O => \N__74273\,
            I => \N__74247\
        );

    \I__18093\ : Span4Mux_h
    port map (
            O => \N__74270\,
            I => \N__74247\
        );

    \I__18092\ : Span4Mux_v
    port map (
            O => \N__74267\,
            I => \N__74247\
        );

    \I__18091\ : LocalMux
    port map (
            O => \N__74264\,
            I => \N__74242\
        );

    \I__18090\ : Span4Mux_v
    port map (
            O => \N__74259\,
            I => \N__74242\
        );

    \I__18089\ : LocalMux
    port map (
            O => \N__74256\,
            I => \N__74239\
        );

    \I__18088\ : Span4Mux_v
    port map (
            O => \N__74247\,
            I => \N__74235\
        );

    \I__18087\ : Sp12to4
    port map (
            O => \N__74242\,
            I => \N__74230\
        );

    \I__18086\ : Span12Mux_h
    port map (
            O => \N__74239\,
            I => \N__74230\
        );

    \I__18085\ : InMux
    port map (
            O => \N__74238\,
            I => \N__74227\
        );

    \I__18084\ : Odrv4
    port map (
            O => \N__74235\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__18083\ : Odrv12
    port map (
            O => \N__74230\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__18082\ : LocalMux
    port map (
            O => \N__74227\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__18081\ : InMux
    port map (
            O => \N__74220\,
            I => \N__74217\
        );

    \I__18080\ : LocalMux
    port map (
            O => \N__74217\,
            I => \N__74213\
        );

    \I__18079\ : InMux
    port map (
            O => \N__74216\,
            I => \N__74210\
        );

    \I__18078\ : Span4Mux_h
    port map (
            O => \N__74213\,
            I => \N__74197\
        );

    \I__18077\ : LocalMux
    port map (
            O => \N__74210\,
            I => \N__74197\
        );

    \I__18076\ : InMux
    port map (
            O => \N__74209\,
            I => \N__74194\
        );

    \I__18075\ : InMux
    port map (
            O => \N__74208\,
            I => \N__74189\
        );

    \I__18074\ : InMux
    port map (
            O => \N__74207\,
            I => \N__74189\
        );

    \I__18073\ : InMux
    port map (
            O => \N__74206\,
            I => \N__74184\
        );

    \I__18072\ : InMux
    port map (
            O => \N__74205\,
            I => \N__74181\
        );

    \I__18071\ : InMux
    port map (
            O => \N__74204\,
            I => \N__74171\
        );

    \I__18070\ : InMux
    port map (
            O => \N__74203\,
            I => \N__74171\
        );

    \I__18069\ : InMux
    port map (
            O => \N__74202\,
            I => \N__74171\
        );

    \I__18068\ : Span4Mux_v
    port map (
            O => \N__74197\,
            I => \N__74166\
        );

    \I__18067\ : LocalMux
    port map (
            O => \N__74194\,
            I => \N__74166\
        );

    \I__18066\ : LocalMux
    port map (
            O => \N__74189\,
            I => \N__74163\
        );

    \I__18065\ : InMux
    port map (
            O => \N__74188\,
            I => \N__74158\
        );

    \I__18064\ : InMux
    port map (
            O => \N__74187\,
            I => \N__74158\
        );

    \I__18063\ : LocalMux
    port map (
            O => \N__74184\,
            I => \N__74151\
        );

    \I__18062\ : LocalMux
    port map (
            O => \N__74181\,
            I => \N__74151\
        );

    \I__18061\ : InMux
    port map (
            O => \N__74180\,
            I => \N__74147\
        );

    \I__18060\ : InMux
    port map (
            O => \N__74179\,
            I => \N__74142\
        );

    \I__18059\ : InMux
    port map (
            O => \N__74178\,
            I => \N__74139\
        );

    \I__18058\ : LocalMux
    port map (
            O => \N__74171\,
            I => \N__74136\
        );

    \I__18057\ : Span4Mux_h
    port map (
            O => \N__74166\,
            I => \N__74132\
        );

    \I__18056\ : Span4Mux_v
    port map (
            O => \N__74163\,
            I => \N__74127\
        );

    \I__18055\ : LocalMux
    port map (
            O => \N__74158\,
            I => \N__74127\
        );

    \I__18054\ : InMux
    port map (
            O => \N__74157\,
            I => \N__74124\
        );

    \I__18053\ : InMux
    port map (
            O => \N__74156\,
            I => \N__74121\
        );

    \I__18052\ : Span4Mux_h
    port map (
            O => \N__74151\,
            I => \N__74118\
        );

    \I__18051\ : InMux
    port map (
            O => \N__74150\,
            I => \N__74112\
        );

    \I__18050\ : LocalMux
    port map (
            O => \N__74147\,
            I => \N__74108\
        );

    \I__18049\ : InMux
    port map (
            O => \N__74146\,
            I => \N__74105\
        );

    \I__18048\ : InMux
    port map (
            O => \N__74145\,
            I => \N__74101\
        );

    \I__18047\ : LocalMux
    port map (
            O => \N__74142\,
            I => \N__74098\
        );

    \I__18046\ : LocalMux
    port map (
            O => \N__74139\,
            I => \N__74095\
        );

    \I__18045\ : Span4Mux_v
    port map (
            O => \N__74136\,
            I => \N__74092\
        );

    \I__18044\ : InMux
    port map (
            O => \N__74135\,
            I => \N__74089\
        );

    \I__18043\ : Span4Mux_h
    port map (
            O => \N__74132\,
            I => \N__74086\
        );

    \I__18042\ : Span4Mux_h
    port map (
            O => \N__74127\,
            I => \N__74081\
        );

    \I__18041\ : LocalMux
    port map (
            O => \N__74124\,
            I => \N__74081\
        );

    \I__18040\ : LocalMux
    port map (
            O => \N__74121\,
            I => \N__74076\
        );

    \I__18039\ : Span4Mux_h
    port map (
            O => \N__74118\,
            I => \N__74076\
        );

    \I__18038\ : InMux
    port map (
            O => \N__74117\,
            I => \N__74073\
        );

    \I__18037\ : InMux
    port map (
            O => \N__74116\,
            I => \N__74070\
        );

    \I__18036\ : InMux
    port map (
            O => \N__74115\,
            I => \N__74063\
        );

    \I__18035\ : LocalMux
    port map (
            O => \N__74112\,
            I => \N__74060\
        );

    \I__18034\ : InMux
    port map (
            O => \N__74111\,
            I => \N__74057\
        );

    \I__18033\ : Span4Mux_v
    port map (
            O => \N__74108\,
            I => \N__74052\
        );

    \I__18032\ : LocalMux
    port map (
            O => \N__74105\,
            I => \N__74052\
        );

    \I__18031\ : InMux
    port map (
            O => \N__74104\,
            I => \N__74048\
        );

    \I__18030\ : LocalMux
    port map (
            O => \N__74101\,
            I => \N__74045\
        );

    \I__18029\ : Span4Mux_v
    port map (
            O => \N__74098\,
            I => \N__74040\
        );

    \I__18028\ : Span4Mux_v
    port map (
            O => \N__74095\,
            I => \N__74040\
        );

    \I__18027\ : Sp12to4
    port map (
            O => \N__74092\,
            I => \N__74035\
        );

    \I__18026\ : LocalMux
    port map (
            O => \N__74089\,
            I => \N__74035\
        );

    \I__18025\ : Span4Mux_v
    port map (
            O => \N__74086\,
            I => \N__74030\
        );

    \I__18024\ : Span4Mux_v
    port map (
            O => \N__74081\,
            I => \N__74030\
        );

    \I__18023\ : Span4Mux_v
    port map (
            O => \N__74076\,
            I => \N__74025\
        );

    \I__18022\ : LocalMux
    port map (
            O => \N__74073\,
            I => \N__74025\
        );

    \I__18021\ : LocalMux
    port map (
            O => \N__74070\,
            I => \N__74022\
        );

    \I__18020\ : InMux
    port map (
            O => \N__74069\,
            I => \N__74018\
        );

    \I__18019\ : InMux
    port map (
            O => \N__74068\,
            I => \N__74015\
        );

    \I__18018\ : InMux
    port map (
            O => \N__74067\,
            I => \N__74010\
        );

    \I__18017\ : InMux
    port map (
            O => \N__74066\,
            I => \N__74010\
        );

    \I__18016\ : LocalMux
    port map (
            O => \N__74063\,
            I => \N__74003\
        );

    \I__18015\ : Span4Mux_h
    port map (
            O => \N__74060\,
            I => \N__74003\
        );

    \I__18014\ : LocalMux
    port map (
            O => \N__74057\,
            I => \N__74003\
        );

    \I__18013\ : Span4Mux_h
    port map (
            O => \N__74052\,
            I => \N__74000\
        );

    \I__18012\ : InMux
    port map (
            O => \N__74051\,
            I => \N__73997\
        );

    \I__18011\ : LocalMux
    port map (
            O => \N__74048\,
            I => \N__73990\
        );

    \I__18010\ : Span4Mux_v
    port map (
            O => \N__74045\,
            I => \N__73990\
        );

    \I__18009\ : Span4Mux_h
    port map (
            O => \N__74040\,
            I => \N__73990\
        );

    \I__18008\ : Span12Mux_h
    port map (
            O => \N__74035\,
            I => \N__73981\
        );

    \I__18007\ : Sp12to4
    port map (
            O => \N__74030\,
            I => \N__73981\
        );

    \I__18006\ : Sp12to4
    port map (
            O => \N__74025\,
            I => \N__73981\
        );

    \I__18005\ : Sp12to4
    port map (
            O => \N__74022\,
            I => \N__73981\
        );

    \I__18004\ : InMux
    port map (
            O => \N__74021\,
            I => \N__73978\
        );

    \I__18003\ : LocalMux
    port map (
            O => \N__74018\,
            I => \N__73975\
        );

    \I__18002\ : LocalMux
    port map (
            O => \N__74015\,
            I => \N__73972\
        );

    \I__18001\ : LocalMux
    port map (
            O => \N__74010\,
            I => \N__73967\
        );

    \I__18000\ : Span4Mux_h
    port map (
            O => \N__74003\,
            I => \N__73967\
        );

    \I__17999\ : Span4Mux_v
    port map (
            O => \N__74000\,
            I => \N__73964\
        );

    \I__17998\ : LocalMux
    port map (
            O => \N__73997\,
            I => \N__73957\
        );

    \I__17997\ : Sp12to4
    port map (
            O => \N__73990\,
            I => \N__73957\
        );

    \I__17996\ : Span12Mux_v
    port map (
            O => \N__73981\,
            I => \N__73957\
        );

    \I__17995\ : LocalMux
    port map (
            O => \N__73978\,
            I => \c0.n9_adj_4601\
        );

    \I__17994\ : Odrv4
    port map (
            O => \N__73975\,
            I => \c0.n9_adj_4601\
        );

    \I__17993\ : Odrv4
    port map (
            O => \N__73972\,
            I => \c0.n9_adj_4601\
        );

    \I__17992\ : Odrv4
    port map (
            O => \N__73967\,
            I => \c0.n9_adj_4601\
        );

    \I__17991\ : Odrv4
    port map (
            O => \N__73964\,
            I => \c0.n9_adj_4601\
        );

    \I__17990\ : Odrv12
    port map (
            O => \N__73957\,
            I => \c0.n9_adj_4601\
        );

    \I__17989\ : InMux
    port map (
            O => \N__73944\,
            I => \N__73940\
        );

    \I__17988\ : InMux
    port map (
            O => \N__73943\,
            I => \N__73936\
        );

    \I__17987\ : LocalMux
    port map (
            O => \N__73940\,
            I => \N__73933\
        );

    \I__17986\ : CascadeMux
    port map (
            O => \N__73939\,
            I => \N__73930\
        );

    \I__17985\ : LocalMux
    port map (
            O => \N__73936\,
            I => \N__73927\
        );

    \I__17984\ : Span4Mux_v
    port map (
            O => \N__73933\,
            I => \N__73924\
        );

    \I__17983\ : InMux
    port map (
            O => \N__73930\,
            I => \N__73921\
        );

    \I__17982\ : Span4Mux_h
    port map (
            O => \N__73927\,
            I => \N__73918\
        );

    \I__17981\ : Span4Mux_h
    port map (
            O => \N__73924\,
            I => \N__73915\
        );

    \I__17980\ : LocalMux
    port map (
            O => \N__73921\,
            I => \c0.data_in_frame_25_1\
        );

    \I__17979\ : Odrv4
    port map (
            O => \N__73918\,
            I => \c0.data_in_frame_25_1\
        );

    \I__17978\ : Odrv4
    port map (
            O => \N__73915\,
            I => \c0.data_in_frame_25_1\
        );

    \I__17977\ : CascadeMux
    port map (
            O => \N__73908\,
            I => \N__73905\
        );

    \I__17976\ : InMux
    port map (
            O => \N__73905\,
            I => \N__73902\
        );

    \I__17975\ : LocalMux
    port map (
            O => \N__73902\,
            I => \N__73896\
        );

    \I__17974\ : CascadeMux
    port map (
            O => \N__73901\,
            I => \N__73893\
        );

    \I__17973\ : InMux
    port map (
            O => \N__73900\,
            I => \N__73890\
        );

    \I__17972\ : InMux
    port map (
            O => \N__73899\,
            I => \N__73887\
        );

    \I__17971\ : Span4Mux_h
    port map (
            O => \N__73896\,
            I => \N__73884\
        );

    \I__17970\ : InMux
    port map (
            O => \N__73893\,
            I => \N__73881\
        );

    \I__17969\ : LocalMux
    port map (
            O => \N__73890\,
            I => \N__73876\
        );

    \I__17968\ : LocalMux
    port map (
            O => \N__73887\,
            I => \N__73876\
        );

    \I__17967\ : Span4Mux_v
    port map (
            O => \N__73884\,
            I => \N__73873\
        );

    \I__17966\ : LocalMux
    port map (
            O => \N__73881\,
            I => \N__73868\
        );

    \I__17965\ : Span4Mux_v
    port map (
            O => \N__73876\,
            I => \N__73868\
        );

    \I__17964\ : Odrv4
    port map (
            O => \N__73873\,
            I => \c0.data_in_frame_20_0\
        );

    \I__17963\ : Odrv4
    port map (
            O => \N__73868\,
            I => \c0.data_in_frame_20_0\
        );

    \I__17962\ : CascadeMux
    port map (
            O => \N__73863\,
            I => \N__73858\
        );

    \I__17961\ : CascadeMux
    port map (
            O => \N__73862\,
            I => \N__73855\
        );

    \I__17960\ : CascadeMux
    port map (
            O => \N__73861\,
            I => \N__73851\
        );

    \I__17959\ : InMux
    port map (
            O => \N__73858\,
            I => \N__73848\
        );

    \I__17958\ : InMux
    port map (
            O => \N__73855\,
            I => \N__73843\
        );

    \I__17957\ : InMux
    port map (
            O => \N__73854\,
            I => \N__73843\
        );

    \I__17956\ : InMux
    port map (
            O => \N__73851\,
            I => \N__73840\
        );

    \I__17955\ : LocalMux
    port map (
            O => \N__73848\,
            I => \N__73837\
        );

    \I__17954\ : LocalMux
    port map (
            O => \N__73843\,
            I => \N__73834\
        );

    \I__17953\ : LocalMux
    port map (
            O => \N__73840\,
            I => \N__73831\
        );

    \I__17952\ : Span4Mux_v
    port map (
            O => \N__73837\,
            I => \N__73828\
        );

    \I__17951\ : Span4Mux_h
    port map (
            O => \N__73834\,
            I => \N__73825\
        );

    \I__17950\ : Span4Mux_h
    port map (
            O => \N__73831\,
            I => \N__73822\
        );

    \I__17949\ : Span4Mux_h
    port map (
            O => \N__73828\,
            I => \N__73817\
        );

    \I__17948\ : Span4Mux_h
    port map (
            O => \N__73825\,
            I => \N__73817\
        );

    \I__17947\ : Span4Mux_h
    port map (
            O => \N__73822\,
            I => \N__73814\
        );

    \I__17946\ : Odrv4
    port map (
            O => \N__73817\,
            I => \c0.data_in_frame_19_0\
        );

    \I__17945\ : Odrv4
    port map (
            O => \N__73814\,
            I => \c0.data_in_frame_19_0\
        );

    \I__17944\ : InMux
    port map (
            O => \N__73809\,
            I => \N__73806\
        );

    \I__17943\ : LocalMux
    port map (
            O => \N__73806\,
            I => \N__73803\
        );

    \I__17942\ : Span4Mux_h
    port map (
            O => \N__73803\,
            I => \N__73800\
        );

    \I__17941\ : Odrv4
    port map (
            O => \N__73800\,
            I => \c0.n12_adj_4564\
        );

    \I__17940\ : InMux
    port map (
            O => \N__73797\,
            I => \N__73793\
        );

    \I__17939\ : InMux
    port map (
            O => \N__73796\,
            I => \N__73790\
        );

    \I__17938\ : LocalMux
    port map (
            O => \N__73793\,
            I => \N__73787\
        );

    \I__17937\ : LocalMux
    port map (
            O => \N__73790\,
            I => \N__73784\
        );

    \I__17936\ : Span4Mux_v
    port map (
            O => \N__73787\,
            I => \N__73779\
        );

    \I__17935\ : Span4Mux_h
    port map (
            O => \N__73784\,
            I => \N__73779\
        );

    \I__17934\ : Odrv4
    port map (
            O => \N__73779\,
            I => \c0.n21404\
        );

    \I__17933\ : CascadeMux
    port map (
            O => \N__73776\,
            I => \c0.n6_adj_4462_cascade_\
        );

    \I__17932\ : InMux
    port map (
            O => \N__73773\,
            I => \N__73769\
        );

    \I__17931\ : InMux
    port map (
            O => \N__73772\,
            I => \N__73766\
        );

    \I__17930\ : LocalMux
    port map (
            O => \N__73769\,
            I => \N__73763\
        );

    \I__17929\ : LocalMux
    port map (
            O => \N__73766\,
            I => \N__73760\
        );

    \I__17928\ : Span4Mux_v
    port map (
            O => \N__73763\,
            I => \N__73755\
        );

    \I__17927\ : Span4Mux_h
    port map (
            O => \N__73760\,
            I => \N__73755\
        );

    \I__17926\ : Odrv4
    port map (
            O => \N__73755\,
            I => \c0.n22562\
        );

    \I__17925\ : CascadeMux
    port map (
            O => \N__73752\,
            I => \N__73747\
        );

    \I__17924\ : InMux
    port map (
            O => \N__73751\,
            I => \N__73744\
        );

    \I__17923\ : InMux
    port map (
            O => \N__73750\,
            I => \N__73741\
        );

    \I__17922\ : InMux
    port map (
            O => \N__73747\,
            I => \N__73738\
        );

    \I__17921\ : LocalMux
    port map (
            O => \N__73744\,
            I => \N__73735\
        );

    \I__17920\ : LocalMux
    port map (
            O => \N__73741\,
            I => \N__73727\
        );

    \I__17919\ : LocalMux
    port map (
            O => \N__73738\,
            I => \N__73727\
        );

    \I__17918\ : Span4Mux_v
    port map (
            O => \N__73735\,
            I => \N__73727\
        );

    \I__17917\ : InMux
    port map (
            O => \N__73734\,
            I => \N__73724\
        );

    \I__17916\ : Odrv4
    port map (
            O => \N__73727\,
            I => data_in_frame_22_3
        );

    \I__17915\ : LocalMux
    port map (
            O => \N__73724\,
            I => data_in_frame_22_3
        );

    \I__17914\ : CascadeMux
    port map (
            O => \N__73719\,
            I => \N__73711\
        );

    \I__17913\ : InMux
    port map (
            O => \N__73718\,
            I => \N__73697\
        );

    \I__17912\ : InMux
    port map (
            O => \N__73717\,
            I => \N__73697\
        );

    \I__17911\ : InMux
    port map (
            O => \N__73716\,
            I => \N__73681\
        );

    \I__17910\ : InMux
    port map (
            O => \N__73715\,
            I => \N__73670\
        );

    \I__17909\ : InMux
    port map (
            O => \N__73714\,
            I => \N__73670\
        );

    \I__17908\ : InMux
    port map (
            O => \N__73711\,
            I => \N__73670\
        );

    \I__17907\ : InMux
    port map (
            O => \N__73710\,
            I => \N__73670\
        );

    \I__17906\ : InMux
    port map (
            O => \N__73709\,
            I => \N__73670\
        );

    \I__17905\ : InMux
    port map (
            O => \N__73708\,
            I => \N__73662\
        );

    \I__17904\ : InMux
    port map (
            O => \N__73707\,
            I => \N__73659\
        );

    \I__17903\ : InMux
    port map (
            O => \N__73706\,
            I => \N__73655\
        );

    \I__17902\ : InMux
    port map (
            O => \N__73705\,
            I => \N__73652\
        );

    \I__17901\ : InMux
    port map (
            O => \N__73704\,
            I => \N__73644\
        );

    \I__17900\ : InMux
    port map (
            O => \N__73703\,
            I => \N__73644\
        );

    \I__17899\ : InMux
    port map (
            O => \N__73702\,
            I => \N__73644\
        );

    \I__17898\ : LocalMux
    port map (
            O => \N__73697\,
            I => \N__73641\
        );

    \I__17897\ : InMux
    port map (
            O => \N__73696\,
            I => \N__73630\
        );

    \I__17896\ : InMux
    port map (
            O => \N__73695\,
            I => \N__73630\
        );

    \I__17895\ : InMux
    port map (
            O => \N__73694\,
            I => \N__73630\
        );

    \I__17894\ : InMux
    port map (
            O => \N__73693\,
            I => \N__73630\
        );

    \I__17893\ : InMux
    port map (
            O => \N__73692\,
            I => \N__73630\
        );

    \I__17892\ : InMux
    port map (
            O => \N__73691\,
            I => \N__73623\
        );

    \I__17891\ : InMux
    port map (
            O => \N__73690\,
            I => \N__73623\
        );

    \I__17890\ : InMux
    port map (
            O => \N__73689\,
            I => \N__73623\
        );

    \I__17889\ : InMux
    port map (
            O => \N__73688\,
            I => \N__73620\
        );

    \I__17888\ : InMux
    port map (
            O => \N__73687\,
            I => \N__73615\
        );

    \I__17887\ : InMux
    port map (
            O => \N__73686\,
            I => \N__73615\
        );

    \I__17886\ : CascadeMux
    port map (
            O => \N__73685\,
            I => \N__73612\
        );

    \I__17885\ : CascadeMux
    port map (
            O => \N__73684\,
            I => \N__73605\
        );

    \I__17884\ : LocalMux
    port map (
            O => \N__73681\,
            I => \N__73602\
        );

    \I__17883\ : LocalMux
    port map (
            O => \N__73670\,
            I => \N__73599\
        );

    \I__17882\ : InMux
    port map (
            O => \N__73669\,
            I => \N__73590\
        );

    \I__17881\ : InMux
    port map (
            O => \N__73668\,
            I => \N__73590\
        );

    \I__17880\ : InMux
    port map (
            O => \N__73667\,
            I => \N__73587\
        );

    \I__17879\ : InMux
    port map (
            O => \N__73666\,
            I => \N__73582\
        );

    \I__17878\ : InMux
    port map (
            O => \N__73665\,
            I => \N__73582\
        );

    \I__17877\ : LocalMux
    port map (
            O => \N__73662\,
            I => \N__73579\
        );

    \I__17876\ : LocalMux
    port map (
            O => \N__73659\,
            I => \N__73576\
        );

    \I__17875\ : InMux
    port map (
            O => \N__73658\,
            I => \N__73573\
        );

    \I__17874\ : LocalMux
    port map (
            O => \N__73655\,
            I => \N__73570\
        );

    \I__17873\ : LocalMux
    port map (
            O => \N__73652\,
            I => \N__73567\
        );

    \I__17872\ : InMux
    port map (
            O => \N__73651\,
            I => \N__73564\
        );

    \I__17871\ : LocalMux
    port map (
            O => \N__73644\,
            I => \N__73561\
        );

    \I__17870\ : Span4Mux_v
    port map (
            O => \N__73641\,
            I => \N__73558\
        );

    \I__17869\ : LocalMux
    port map (
            O => \N__73630\,
            I => \N__73551\
        );

    \I__17868\ : LocalMux
    port map (
            O => \N__73623\,
            I => \N__73551\
        );

    \I__17867\ : LocalMux
    port map (
            O => \N__73620\,
            I => \N__73551\
        );

    \I__17866\ : LocalMux
    port map (
            O => \N__73615\,
            I => \N__73548\
        );

    \I__17865\ : InMux
    port map (
            O => \N__73612\,
            I => \N__73543\
        );

    \I__17864\ : InMux
    port map (
            O => \N__73611\,
            I => \N__73543\
        );

    \I__17863\ : InMux
    port map (
            O => \N__73610\,
            I => \N__73534\
        );

    \I__17862\ : InMux
    port map (
            O => \N__73609\,
            I => \N__73534\
        );

    \I__17861\ : InMux
    port map (
            O => \N__73608\,
            I => \N__73534\
        );

    \I__17860\ : InMux
    port map (
            O => \N__73605\,
            I => \N__73534\
        );

    \I__17859\ : Span4Mux_h
    port map (
            O => \N__73602\,
            I => \N__73529\
        );

    \I__17858\ : Span4Mux_v
    port map (
            O => \N__73599\,
            I => \N__73529\
        );

    \I__17857\ : InMux
    port map (
            O => \N__73598\,
            I => \N__73526\
        );

    \I__17856\ : InMux
    port map (
            O => \N__73597\,
            I => \N__73523\
        );

    \I__17855\ : InMux
    port map (
            O => \N__73596\,
            I => \N__73513\
        );

    \I__17854\ : InMux
    port map (
            O => \N__73595\,
            I => \N__73513\
        );

    \I__17853\ : LocalMux
    port map (
            O => \N__73590\,
            I => \N__73506\
        );

    \I__17852\ : LocalMux
    port map (
            O => \N__73587\,
            I => \N__73506\
        );

    \I__17851\ : LocalMux
    port map (
            O => \N__73582\,
            I => \N__73506\
        );

    \I__17850\ : Span4Mux_v
    port map (
            O => \N__73579\,
            I => \N__73503\
        );

    \I__17849\ : Span4Mux_h
    port map (
            O => \N__73576\,
            I => \N__73500\
        );

    \I__17848\ : LocalMux
    port map (
            O => \N__73573\,
            I => \N__73497\
        );

    \I__17847\ : Span4Mux_h
    port map (
            O => \N__73570\,
            I => \N__73492\
        );

    \I__17846\ : Span4Mux_v
    port map (
            O => \N__73567\,
            I => \N__73492\
        );

    \I__17845\ : LocalMux
    port map (
            O => \N__73564\,
            I => \N__73489\
        );

    \I__17844\ : Span4Mux_h
    port map (
            O => \N__73561\,
            I => \N__73484\
        );

    \I__17843\ : Span4Mux_v
    port map (
            O => \N__73558\,
            I => \N__73484\
        );

    \I__17842\ : Span4Mux_v
    port map (
            O => \N__73551\,
            I => \N__73479\
        );

    \I__17841\ : Span4Mux_h
    port map (
            O => \N__73548\,
            I => \N__73479\
        );

    \I__17840\ : LocalMux
    port map (
            O => \N__73543\,
            I => \N__73472\
        );

    \I__17839\ : LocalMux
    port map (
            O => \N__73534\,
            I => \N__73472\
        );

    \I__17838\ : Span4Mux_v
    port map (
            O => \N__73529\,
            I => \N__73472\
        );

    \I__17837\ : LocalMux
    port map (
            O => \N__73526\,
            I => \N__73467\
        );

    \I__17836\ : LocalMux
    port map (
            O => \N__73523\,
            I => \N__73467\
        );

    \I__17835\ : InMux
    port map (
            O => \N__73522\,
            I => \N__73464\
        );

    \I__17834\ : InMux
    port map (
            O => \N__73521\,
            I => \N__73461\
        );

    \I__17833\ : InMux
    port map (
            O => \N__73520\,
            I => \N__73458\
        );

    \I__17832\ : InMux
    port map (
            O => \N__73519\,
            I => \N__73453\
        );

    \I__17831\ : InMux
    port map (
            O => \N__73518\,
            I => \N__73453\
        );

    \I__17830\ : LocalMux
    port map (
            O => \N__73513\,
            I => \N__73450\
        );

    \I__17829\ : Span12Mux_h
    port map (
            O => \N__73506\,
            I => \N__73447\
        );

    \I__17828\ : Span4Mux_h
    port map (
            O => \N__73503\,
            I => \N__73444\
        );

    \I__17827\ : Span4Mux_v
    port map (
            O => \N__73500\,
            I => \N__73441\
        );

    \I__17826\ : Span4Mux_v
    port map (
            O => \N__73497\,
            I => \N__73436\
        );

    \I__17825\ : Span4Mux_h
    port map (
            O => \N__73492\,
            I => \N__73436\
        );

    \I__17824\ : Span4Mux_h
    port map (
            O => \N__73489\,
            I => \N__73431\
        );

    \I__17823\ : Span4Mux_h
    port map (
            O => \N__73484\,
            I => \N__73431\
        );

    \I__17822\ : Span4Mux_h
    port map (
            O => \N__73479\,
            I => \N__73424\
        );

    \I__17821\ : Span4Mux_v
    port map (
            O => \N__73472\,
            I => \N__73424\
        );

    \I__17820\ : Span4Mux_v
    port map (
            O => \N__73467\,
            I => \N__73424\
        );

    \I__17819\ : LocalMux
    port map (
            O => \N__73464\,
            I => \c0.n22112\
        );

    \I__17818\ : LocalMux
    port map (
            O => \N__73461\,
            I => \c0.n22112\
        );

    \I__17817\ : LocalMux
    port map (
            O => \N__73458\,
            I => \c0.n22112\
        );

    \I__17816\ : LocalMux
    port map (
            O => \N__73453\,
            I => \c0.n22112\
        );

    \I__17815\ : Odrv12
    port map (
            O => \N__73450\,
            I => \c0.n22112\
        );

    \I__17814\ : Odrv12
    port map (
            O => \N__73447\,
            I => \c0.n22112\
        );

    \I__17813\ : Odrv4
    port map (
            O => \N__73444\,
            I => \c0.n22112\
        );

    \I__17812\ : Odrv4
    port map (
            O => \N__73441\,
            I => \c0.n22112\
        );

    \I__17811\ : Odrv4
    port map (
            O => \N__73436\,
            I => \c0.n22112\
        );

    \I__17810\ : Odrv4
    port map (
            O => \N__73431\,
            I => \c0.n22112\
        );

    \I__17809\ : Odrv4
    port map (
            O => \N__73424\,
            I => \c0.n22112\
        );

    \I__17808\ : CascadeMux
    port map (
            O => \N__73401\,
            I => \N__73397\
        );

    \I__17807\ : InMux
    port map (
            O => \N__73400\,
            I => \N__73393\
        );

    \I__17806\ : InMux
    port map (
            O => \N__73397\,
            I => \N__73389\
        );

    \I__17805\ : CascadeMux
    port map (
            O => \N__73396\,
            I => \N__73386\
        );

    \I__17804\ : LocalMux
    port map (
            O => \N__73393\,
            I => \N__73383\
        );

    \I__17803\ : InMux
    port map (
            O => \N__73392\,
            I => \N__73380\
        );

    \I__17802\ : LocalMux
    port map (
            O => \N__73389\,
            I => \N__73377\
        );

    \I__17801\ : InMux
    port map (
            O => \N__73386\,
            I => \N__73374\
        );

    \I__17800\ : Span4Mux_h
    port map (
            O => \N__73383\,
            I => \N__73369\
        );

    \I__17799\ : LocalMux
    port map (
            O => \N__73380\,
            I => \N__73369\
        );

    \I__17798\ : Span4Mux_h
    port map (
            O => \N__73377\,
            I => \N__73366\
        );

    \I__17797\ : LocalMux
    port map (
            O => \N__73374\,
            I => \N__73361\
        );

    \I__17796\ : Span4Mux_v
    port map (
            O => \N__73369\,
            I => \N__73361\
        );

    \I__17795\ : Odrv4
    port map (
            O => \N__73366\,
            I => \c0.data_in_frame_15_0\
        );

    \I__17794\ : Odrv4
    port map (
            O => \N__73361\,
            I => \c0.data_in_frame_15_0\
        );

    \I__17793\ : CascadeMux
    port map (
            O => \N__73356\,
            I => \N__73353\
        );

    \I__17792\ : InMux
    port map (
            O => \N__73353\,
            I => \N__73350\
        );

    \I__17791\ : LocalMux
    port map (
            O => \N__73350\,
            I => \N__73343\
        );

    \I__17790\ : InMux
    port map (
            O => \N__73349\,
            I => \N__73338\
        );

    \I__17789\ : InMux
    port map (
            O => \N__73348\,
            I => \N__73338\
        );

    \I__17788\ : CascadeMux
    port map (
            O => \N__73347\,
            I => \N__73332\
        );

    \I__17787\ : InMux
    port map (
            O => \N__73346\,
            I => \N__73327\
        );

    \I__17786\ : Span4Mux_v
    port map (
            O => \N__73343\,
            I => \N__73321\
        );

    \I__17785\ : LocalMux
    port map (
            O => \N__73338\,
            I => \N__73321\
        );

    \I__17784\ : InMux
    port map (
            O => \N__73337\,
            I => \N__73316\
        );

    \I__17783\ : InMux
    port map (
            O => \N__73336\,
            I => \N__73316\
        );

    \I__17782\ : InMux
    port map (
            O => \N__73335\,
            I => \N__73313\
        );

    \I__17781\ : InMux
    port map (
            O => \N__73332\,
            I => \N__73308\
        );

    \I__17780\ : InMux
    port map (
            O => \N__73331\,
            I => \N__73308\
        );

    \I__17779\ : InMux
    port map (
            O => \N__73330\,
            I => \N__73304\
        );

    \I__17778\ : LocalMux
    port map (
            O => \N__73327\,
            I => \N__73301\
        );

    \I__17777\ : InMux
    port map (
            O => \N__73326\,
            I => \N__73295\
        );

    \I__17776\ : Span4Mux_v
    port map (
            O => \N__73321\,
            I => \N__73286\
        );

    \I__17775\ : LocalMux
    port map (
            O => \N__73316\,
            I => \N__73283\
        );

    \I__17774\ : LocalMux
    port map (
            O => \N__73313\,
            I => \N__73280\
        );

    \I__17773\ : LocalMux
    port map (
            O => \N__73308\,
            I => \N__73277\
        );

    \I__17772\ : CascadeMux
    port map (
            O => \N__73307\,
            I => \N__73273\
        );

    \I__17771\ : LocalMux
    port map (
            O => \N__73304\,
            I => \N__73270\
        );

    \I__17770\ : Span4Mux_h
    port map (
            O => \N__73301\,
            I => \N__73267\
        );

    \I__17769\ : InMux
    port map (
            O => \N__73300\,
            I => \N__73264\
        );

    \I__17768\ : InMux
    port map (
            O => \N__73299\,
            I => \N__73261\
        );

    \I__17767\ : InMux
    port map (
            O => \N__73298\,
            I => \N__73258\
        );

    \I__17766\ : LocalMux
    port map (
            O => \N__73295\,
            I => \N__73255\
        );

    \I__17765\ : InMux
    port map (
            O => \N__73294\,
            I => \N__73250\
        );

    \I__17764\ : InMux
    port map (
            O => \N__73293\,
            I => \N__73250\
        );

    \I__17763\ : InMux
    port map (
            O => \N__73292\,
            I => \N__73245\
        );

    \I__17762\ : InMux
    port map (
            O => \N__73291\,
            I => \N__73245\
        );

    \I__17761\ : InMux
    port map (
            O => \N__73290\,
            I => \N__73242\
        );

    \I__17760\ : InMux
    port map (
            O => \N__73289\,
            I => \N__73239\
        );

    \I__17759\ : Span4Mux_h
    port map (
            O => \N__73286\,
            I => \N__73234\
        );

    \I__17758\ : Span4Mux_v
    port map (
            O => \N__73283\,
            I => \N__73234\
        );

    \I__17757\ : Span4Mux_h
    port map (
            O => \N__73280\,
            I => \N__73229\
        );

    \I__17756\ : Span4Mux_v
    port map (
            O => \N__73277\,
            I => \N__73229\
        );

    \I__17755\ : InMux
    port map (
            O => \N__73276\,
            I => \N__73226\
        );

    \I__17754\ : InMux
    port map (
            O => \N__73273\,
            I => \N__73223\
        );

    \I__17753\ : Span4Mux_h
    port map (
            O => \N__73270\,
            I => \N__73220\
        );

    \I__17752\ : Span4Mux_v
    port map (
            O => \N__73267\,
            I => \N__73215\
        );

    \I__17751\ : LocalMux
    port map (
            O => \N__73264\,
            I => \N__73215\
        );

    \I__17750\ : LocalMux
    port map (
            O => \N__73261\,
            I => \N__73211\
        );

    \I__17749\ : LocalMux
    port map (
            O => \N__73258\,
            I => \N__73202\
        );

    \I__17748\ : Span4Mux_h
    port map (
            O => \N__73255\,
            I => \N__73202\
        );

    \I__17747\ : LocalMux
    port map (
            O => \N__73250\,
            I => \N__73196\
        );

    \I__17746\ : LocalMux
    port map (
            O => \N__73245\,
            I => \N__73196\
        );

    \I__17745\ : LocalMux
    port map (
            O => \N__73242\,
            I => \N__73187\
        );

    \I__17744\ : LocalMux
    port map (
            O => \N__73239\,
            I => \N__73187\
        );

    \I__17743\ : Span4Mux_h
    port map (
            O => \N__73234\,
            I => \N__73187\
        );

    \I__17742\ : Span4Mux_v
    port map (
            O => \N__73229\,
            I => \N__73187\
        );

    \I__17741\ : LocalMux
    port map (
            O => \N__73226\,
            I => \N__73182\
        );

    \I__17740\ : LocalMux
    port map (
            O => \N__73223\,
            I => \N__73182\
        );

    \I__17739\ : Span4Mux_v
    port map (
            O => \N__73220\,
            I => \N__73179\
        );

    \I__17738\ : Span4Mux_h
    port map (
            O => \N__73215\,
            I => \N__73176\
        );

    \I__17737\ : InMux
    port map (
            O => \N__73214\,
            I => \N__73173\
        );

    \I__17736\ : Span4Mux_h
    port map (
            O => \N__73211\,
            I => \N__73170\
        );

    \I__17735\ : InMux
    port map (
            O => \N__73210\,
            I => \N__73167\
        );

    \I__17734\ : InMux
    port map (
            O => \N__73209\,
            I => \N__73160\
        );

    \I__17733\ : InMux
    port map (
            O => \N__73208\,
            I => \N__73160\
        );

    \I__17732\ : InMux
    port map (
            O => \N__73207\,
            I => \N__73160\
        );

    \I__17731\ : Span4Mux_h
    port map (
            O => \N__73202\,
            I => \N__73157\
        );

    \I__17730\ : InMux
    port map (
            O => \N__73201\,
            I => \N__73150\
        );

    \I__17729\ : Span4Mux_v
    port map (
            O => \N__73196\,
            I => \N__73147\
        );

    \I__17728\ : Span4Mux_v
    port map (
            O => \N__73187\,
            I => \N__73144\
        );

    \I__17727\ : Sp12to4
    port map (
            O => \N__73182\,
            I => \N__73137\
        );

    \I__17726\ : Sp12to4
    port map (
            O => \N__73179\,
            I => \N__73137\
        );

    \I__17725\ : Sp12to4
    port map (
            O => \N__73176\,
            I => \N__73137\
        );

    \I__17724\ : LocalMux
    port map (
            O => \N__73173\,
            I => \N__73134\
        );

    \I__17723\ : Span4Mux_h
    port map (
            O => \N__73170\,
            I => \N__73131\
        );

    \I__17722\ : LocalMux
    port map (
            O => \N__73167\,
            I => \N__73124\
        );

    \I__17721\ : LocalMux
    port map (
            O => \N__73160\,
            I => \N__73124\
        );

    \I__17720\ : Sp12to4
    port map (
            O => \N__73157\,
            I => \N__73124\
        );

    \I__17719\ : InMux
    port map (
            O => \N__73156\,
            I => \N__73121\
        );

    \I__17718\ : InMux
    port map (
            O => \N__73155\,
            I => \N__73118\
        );

    \I__17717\ : InMux
    port map (
            O => \N__73154\,
            I => \N__73113\
        );

    \I__17716\ : InMux
    port map (
            O => \N__73153\,
            I => \N__73113\
        );

    \I__17715\ : LocalMux
    port map (
            O => \N__73150\,
            I => \N__73110\
        );

    \I__17714\ : Sp12to4
    port map (
            O => \N__73147\,
            I => \N__73103\
        );

    \I__17713\ : Sp12to4
    port map (
            O => \N__73144\,
            I => \N__73103\
        );

    \I__17712\ : Span12Mux_v
    port map (
            O => \N__73137\,
            I => \N__73103\
        );

    \I__17711\ : Span12Mux_h
    port map (
            O => \N__73134\,
            I => \N__73096\
        );

    \I__17710\ : Sp12to4
    port map (
            O => \N__73131\,
            I => \N__73096\
        );

    \I__17709\ : Span12Mux_v
    port map (
            O => \N__73124\,
            I => \N__73096\
        );

    \I__17708\ : LocalMux
    port map (
            O => \N__73121\,
            I => rx_data_6
        );

    \I__17707\ : LocalMux
    port map (
            O => \N__73118\,
            I => rx_data_6
        );

    \I__17706\ : LocalMux
    port map (
            O => \N__73113\,
            I => rx_data_6
        );

    \I__17705\ : Odrv4
    port map (
            O => \N__73110\,
            I => rx_data_6
        );

    \I__17704\ : Odrv12
    port map (
            O => \N__73103\,
            I => rx_data_6
        );

    \I__17703\ : Odrv12
    port map (
            O => \N__73096\,
            I => rx_data_6
        );

    \I__17702\ : CascadeMux
    port map (
            O => \N__73083\,
            I => \N__73078\
        );

    \I__17701\ : CascadeMux
    port map (
            O => \N__73082\,
            I => \N__73075\
        );

    \I__17700\ : InMux
    port map (
            O => \N__73081\,
            I => \N__73072\
        );

    \I__17699\ : InMux
    port map (
            O => \N__73078\,
            I => \N__73067\
        );

    \I__17698\ : InMux
    port map (
            O => \N__73075\,
            I => \N__73067\
        );

    \I__17697\ : LocalMux
    port map (
            O => \N__73072\,
            I => \N__73064\
        );

    \I__17696\ : LocalMux
    port map (
            O => \N__73067\,
            I => data_in_frame_22_1
        );

    \I__17695\ : Odrv4
    port map (
            O => \N__73064\,
            I => data_in_frame_22_1
        );

    \I__17694\ : CascadeMux
    port map (
            O => \N__73059\,
            I => \N__73056\
        );

    \I__17693\ : InMux
    port map (
            O => \N__73056\,
            I => \N__73052\
        );

    \I__17692\ : InMux
    port map (
            O => \N__73055\,
            I => \N__73049\
        );

    \I__17691\ : LocalMux
    port map (
            O => \N__73052\,
            I => \N__73046\
        );

    \I__17690\ : LocalMux
    port map (
            O => \N__73049\,
            I => \N__73043\
        );

    \I__17689\ : Odrv4
    port map (
            O => \N__73046\,
            I => \c0.data_in_frame_20_2\
        );

    \I__17688\ : Odrv4
    port map (
            O => \N__73043\,
            I => \c0.data_in_frame_20_2\
        );

    \I__17687\ : CascadeMux
    port map (
            O => \N__73038\,
            I => \N__73035\
        );

    \I__17686\ : InMux
    port map (
            O => \N__73035\,
            I => \N__73030\
        );

    \I__17685\ : InMux
    port map (
            O => \N__73034\,
            I => \N__73027\
        );

    \I__17684\ : InMux
    port map (
            O => \N__73033\,
            I => \N__73024\
        );

    \I__17683\ : LocalMux
    port map (
            O => \N__73030\,
            I => \N__73021\
        );

    \I__17682\ : LocalMux
    port map (
            O => \N__73027\,
            I => \N__73015\
        );

    \I__17681\ : LocalMux
    port map (
            O => \N__73024\,
            I => \N__73015\
        );

    \I__17680\ : Span4Mux_h
    port map (
            O => \N__73021\,
            I => \N__73012\
        );

    \I__17679\ : InMux
    port map (
            O => \N__73020\,
            I => \N__73009\
        );

    \I__17678\ : Span4Mux_h
    port map (
            O => \N__73015\,
            I => \N__73006\
        );

    \I__17677\ : Span4Mux_v
    port map (
            O => \N__73012\,
            I => \N__73003\
        );

    \I__17676\ : LocalMux
    port map (
            O => \N__73009\,
            I => \c0.data_in_frame_23_5\
        );

    \I__17675\ : Odrv4
    port map (
            O => \N__73006\,
            I => \c0.data_in_frame_23_5\
        );

    \I__17674\ : Odrv4
    port map (
            O => \N__73003\,
            I => \c0.data_in_frame_23_5\
        );

    \I__17673\ : CascadeMux
    port map (
            O => \N__72996\,
            I => \N__72993\
        );

    \I__17672\ : InMux
    port map (
            O => \N__72993\,
            I => \N__72986\
        );

    \I__17671\ : CascadeMux
    port map (
            O => \N__72992\,
            I => \N__72983\
        );

    \I__17670\ : InMux
    port map (
            O => \N__72991\,
            I => \N__72974\
        );

    \I__17669\ : InMux
    port map (
            O => \N__72990\,
            I => \N__72971\
        );

    \I__17668\ : InMux
    port map (
            O => \N__72989\,
            I => \N__72968\
        );

    \I__17667\ : LocalMux
    port map (
            O => \N__72986\,
            I => \N__72961\
        );

    \I__17666\ : InMux
    port map (
            O => \N__72983\,
            I => \N__72956\
        );

    \I__17665\ : InMux
    port map (
            O => \N__72982\,
            I => \N__72956\
        );

    \I__17664\ : InMux
    port map (
            O => \N__72981\,
            I => \N__72949\
        );

    \I__17663\ : InMux
    port map (
            O => \N__72980\,
            I => \N__72949\
        );

    \I__17662\ : InMux
    port map (
            O => \N__72979\,
            I => \N__72949\
        );

    \I__17661\ : CascadeMux
    port map (
            O => \N__72978\,
            I => \N__72946\
        );

    \I__17660\ : CascadeMux
    port map (
            O => \N__72977\,
            I => \N__72943\
        );

    \I__17659\ : LocalMux
    port map (
            O => \N__72974\,
            I => \N__72932\
        );

    \I__17658\ : LocalMux
    port map (
            O => \N__72971\,
            I => \N__72929\
        );

    \I__17657\ : LocalMux
    port map (
            O => \N__72968\,
            I => \N__72926\
        );

    \I__17656\ : CascadeMux
    port map (
            O => \N__72967\,
            I => \N__72920\
        );

    \I__17655\ : CascadeMux
    port map (
            O => \N__72966\,
            I => \N__72917\
        );

    \I__17654\ : InMux
    port map (
            O => \N__72965\,
            I => \N__72912\
        );

    \I__17653\ : InMux
    port map (
            O => \N__72964\,
            I => \N__72912\
        );

    \I__17652\ : Span4Mux_h
    port map (
            O => \N__72961\,
            I => \N__72909\
        );

    \I__17651\ : LocalMux
    port map (
            O => \N__72956\,
            I => \N__72906\
        );

    \I__17650\ : LocalMux
    port map (
            O => \N__72949\,
            I => \N__72903\
        );

    \I__17649\ : InMux
    port map (
            O => \N__72946\,
            I => \N__72900\
        );

    \I__17648\ : InMux
    port map (
            O => \N__72943\,
            I => \N__72893\
        );

    \I__17647\ : InMux
    port map (
            O => \N__72942\,
            I => \N__72893\
        );

    \I__17646\ : InMux
    port map (
            O => \N__72941\,
            I => \N__72890\
        );

    \I__17645\ : InMux
    port map (
            O => \N__72940\,
            I => \N__72887\
        );

    \I__17644\ : InMux
    port map (
            O => \N__72939\,
            I => \N__72884\
        );

    \I__17643\ : InMux
    port map (
            O => \N__72938\,
            I => \N__72881\
        );

    \I__17642\ : InMux
    port map (
            O => \N__72937\,
            I => \N__72875\
        );

    \I__17641\ : InMux
    port map (
            O => \N__72936\,
            I => \N__72875\
        );

    \I__17640\ : InMux
    port map (
            O => \N__72935\,
            I => \N__72872\
        );

    \I__17639\ : Span4Mux_v
    port map (
            O => \N__72932\,
            I => \N__72869\
        );

    \I__17638\ : Span4Mux_h
    port map (
            O => \N__72929\,
            I => \N__72866\
        );

    \I__17637\ : Span4Mux_h
    port map (
            O => \N__72926\,
            I => \N__72863\
        );

    \I__17636\ : InMux
    port map (
            O => \N__72925\,
            I => \N__72857\
        );

    \I__17635\ : InMux
    port map (
            O => \N__72924\,
            I => \N__72848\
        );

    \I__17634\ : InMux
    port map (
            O => \N__72923\,
            I => \N__72848\
        );

    \I__17633\ : InMux
    port map (
            O => \N__72920\,
            I => \N__72848\
        );

    \I__17632\ : InMux
    port map (
            O => \N__72917\,
            I => \N__72848\
        );

    \I__17631\ : LocalMux
    port map (
            O => \N__72912\,
            I => \N__72845\
        );

    \I__17630\ : Span4Mux_h
    port map (
            O => \N__72909\,
            I => \N__72838\
        );

    \I__17629\ : Span4Mux_h
    port map (
            O => \N__72906\,
            I => \N__72838\
        );

    \I__17628\ : Span4Mux_h
    port map (
            O => \N__72903\,
            I => \N__72838\
        );

    \I__17627\ : LocalMux
    port map (
            O => \N__72900\,
            I => \N__72835\
        );

    \I__17626\ : InMux
    port map (
            O => \N__72899\,
            I => \N__72832\
        );

    \I__17625\ : InMux
    port map (
            O => \N__72898\,
            I => \N__72829\
        );

    \I__17624\ : LocalMux
    port map (
            O => \N__72893\,
            I => \N__72826\
        );

    \I__17623\ : LocalMux
    port map (
            O => \N__72890\,
            I => \N__72821\
        );

    \I__17622\ : LocalMux
    port map (
            O => \N__72887\,
            I => \N__72821\
        );

    \I__17621\ : LocalMux
    port map (
            O => \N__72884\,
            I => \N__72816\
        );

    \I__17620\ : LocalMux
    port map (
            O => \N__72881\,
            I => \N__72816\
        );

    \I__17619\ : InMux
    port map (
            O => \N__72880\,
            I => \N__72813\
        );

    \I__17618\ : LocalMux
    port map (
            O => \N__72875\,
            I => \N__72810\
        );

    \I__17617\ : LocalMux
    port map (
            O => \N__72872\,
            I => \N__72805\
        );

    \I__17616\ : Span4Mux_v
    port map (
            O => \N__72869\,
            I => \N__72805\
        );

    \I__17615\ : Span4Mux_v
    port map (
            O => \N__72866\,
            I => \N__72800\
        );

    \I__17614\ : Span4Mux_v
    port map (
            O => \N__72863\,
            I => \N__72800\
        );

    \I__17613\ : InMux
    port map (
            O => \N__72862\,
            I => \N__72797\
        );

    \I__17612\ : InMux
    port map (
            O => \N__72861\,
            I => \N__72792\
        );

    \I__17611\ : InMux
    port map (
            O => \N__72860\,
            I => \N__72792\
        );

    \I__17610\ : LocalMux
    port map (
            O => \N__72857\,
            I => \N__72789\
        );

    \I__17609\ : LocalMux
    port map (
            O => \N__72848\,
            I => \N__72786\
        );

    \I__17608\ : Span4Mux_h
    port map (
            O => \N__72845\,
            I => \N__72781\
        );

    \I__17607\ : Span4Mux_v
    port map (
            O => \N__72838\,
            I => \N__72781\
        );

    \I__17606\ : Span4Mux_v
    port map (
            O => \N__72835\,
            I => \N__72774\
        );

    \I__17605\ : LocalMux
    port map (
            O => \N__72832\,
            I => \N__72774\
        );

    \I__17604\ : LocalMux
    port map (
            O => \N__72829\,
            I => \N__72774\
        );

    \I__17603\ : Span4Mux_h
    port map (
            O => \N__72826\,
            I => \N__72771\
        );

    \I__17602\ : Span4Mux_v
    port map (
            O => \N__72821\,
            I => \N__72768\
        );

    \I__17601\ : Span4Mux_v
    port map (
            O => \N__72816\,
            I => \N__72765\
        );

    \I__17600\ : LocalMux
    port map (
            O => \N__72813\,
            I => \N__72762\
        );

    \I__17599\ : Span4Mux_v
    port map (
            O => \N__72810\,
            I => \N__72759\
        );

    \I__17598\ : Span4Mux_h
    port map (
            O => \N__72805\,
            I => \N__72754\
        );

    \I__17597\ : Span4Mux_v
    port map (
            O => \N__72800\,
            I => \N__72754\
        );

    \I__17596\ : LocalMux
    port map (
            O => \N__72797\,
            I => \N__72751\
        );

    \I__17595\ : LocalMux
    port map (
            O => \N__72792\,
            I => \N__72748\
        );

    \I__17594\ : Span4Mux_h
    port map (
            O => \N__72789\,
            I => \N__72745\
        );

    \I__17593\ : Span4Mux_h
    port map (
            O => \N__72786\,
            I => \N__72740\
        );

    \I__17592\ : Span4Mux_v
    port map (
            O => \N__72781\,
            I => \N__72740\
        );

    \I__17591\ : Span4Mux_h
    port map (
            O => \N__72774\,
            I => \N__72737\
        );

    \I__17590\ : Sp12to4
    port map (
            O => \N__72771\,
            I => \N__72734\
        );

    \I__17589\ : Sp12to4
    port map (
            O => \N__72768\,
            I => \N__72729\
        );

    \I__17588\ : Sp12to4
    port map (
            O => \N__72765\,
            I => \N__72729\
        );

    \I__17587\ : Span4Mux_h
    port map (
            O => \N__72762\,
            I => \N__72722\
        );

    \I__17586\ : Span4Mux_h
    port map (
            O => \N__72759\,
            I => \N__72722\
        );

    \I__17585\ : Span4Mux_v
    port map (
            O => \N__72754\,
            I => \N__72722\
        );

    \I__17584\ : Span12Mux_h
    port map (
            O => \N__72751\,
            I => \N__72717\
        );

    \I__17583\ : Span12Mux_h
    port map (
            O => \N__72748\,
            I => \N__72717\
        );

    \I__17582\ : Span4Mux_h
    port map (
            O => \N__72745\,
            I => \N__72712\
        );

    \I__17581\ : Span4Mux_v
    port map (
            O => \N__72740\,
            I => \N__72712\
        );

    \I__17580\ : Sp12to4
    port map (
            O => \N__72737\,
            I => \N__72705\
        );

    \I__17579\ : Span12Mux_v
    port map (
            O => \N__72734\,
            I => \N__72705\
        );

    \I__17578\ : Span12Mux_h
    port map (
            O => \N__72729\,
            I => \N__72705\
        );

    \I__17577\ : Span4Mux_v
    port map (
            O => \N__72722\,
            I => \N__72702\
        );

    \I__17576\ : Odrv12
    port map (
            O => \N__72717\,
            I => \c0.n9_adj_4563\
        );

    \I__17575\ : Odrv4
    port map (
            O => \N__72712\,
            I => \c0.n9_adj_4563\
        );

    \I__17574\ : Odrv12
    port map (
            O => \N__72705\,
            I => \c0.n9_adj_4563\
        );

    \I__17573\ : Odrv4
    port map (
            O => \N__72702\,
            I => \c0.n9_adj_4563\
        );

    \I__17572\ : CascadeMux
    port map (
            O => \N__72693\,
            I => \N__72690\
        );

    \I__17571\ : InMux
    port map (
            O => \N__72690\,
            I => \N__72686\
        );

    \I__17570\ : InMux
    port map (
            O => \N__72689\,
            I => \N__72683\
        );

    \I__17569\ : LocalMux
    port map (
            O => \N__72686\,
            I => \N__72678\
        );

    \I__17568\ : LocalMux
    port map (
            O => \N__72683\,
            I => \N__72675\
        );

    \I__17567\ : CascadeMux
    port map (
            O => \N__72682\,
            I => \N__72672\
        );

    \I__17566\ : InMux
    port map (
            O => \N__72681\,
            I => \N__72669\
        );

    \I__17565\ : Span4Mux_h
    port map (
            O => \N__72678\,
            I => \N__72666\
        );

    \I__17564\ : Span4Mux_h
    port map (
            O => \N__72675\,
            I => \N__72663\
        );

    \I__17563\ : InMux
    port map (
            O => \N__72672\,
            I => \N__72660\
        );

    \I__17562\ : LocalMux
    port map (
            O => \N__72669\,
            I => \N__72657\
        );

    \I__17561\ : Span4Mux_h
    port map (
            O => \N__72666\,
            I => \N__72654\
        );

    \I__17560\ : Span4Mux_h
    port map (
            O => \N__72663\,
            I => \N__72651\
        );

    \I__17559\ : LocalMux
    port map (
            O => \N__72660\,
            I => \c0.data_in_frame_16_7\
        );

    \I__17558\ : Odrv12
    port map (
            O => \N__72657\,
            I => \c0.data_in_frame_16_7\
        );

    \I__17557\ : Odrv4
    port map (
            O => \N__72654\,
            I => \c0.data_in_frame_16_7\
        );

    \I__17556\ : Odrv4
    port map (
            O => \N__72651\,
            I => \c0.data_in_frame_16_7\
        );

    \I__17555\ : InMux
    port map (
            O => \N__72642\,
            I => \N__72639\
        );

    \I__17554\ : LocalMux
    port map (
            O => \N__72639\,
            I => \N__72635\
        );

    \I__17553\ : InMux
    port map (
            O => \N__72638\,
            I => \N__72632\
        );

    \I__17552\ : Span4Mux_v
    port map (
            O => \N__72635\,
            I => \N__72626\
        );

    \I__17551\ : LocalMux
    port map (
            O => \N__72632\,
            I => \N__72626\
        );

    \I__17550\ : InMux
    port map (
            O => \N__72631\,
            I => \N__72623\
        );

    \I__17549\ : Span4Mux_v
    port map (
            O => \N__72626\,
            I => \N__72620\
        );

    \I__17548\ : LocalMux
    port map (
            O => \N__72623\,
            I => \N__72617\
        );

    \I__17547\ : Odrv4
    port map (
            O => \N__72620\,
            I => \c0.n22_adj_4244\
        );

    \I__17546\ : Odrv4
    port map (
            O => \N__72617\,
            I => \c0.n22_adj_4244\
        );

    \I__17545\ : InMux
    port map (
            O => \N__72612\,
            I => \N__72609\
        );

    \I__17544\ : LocalMux
    port map (
            O => \N__72609\,
            I => \c0.n24_adj_4618\
        );

    \I__17543\ : CascadeMux
    port map (
            O => \N__72606\,
            I => \N__72603\
        );

    \I__17542\ : InMux
    port map (
            O => \N__72603\,
            I => \N__72600\
        );

    \I__17541\ : LocalMux
    port map (
            O => \N__72600\,
            I => \N__72597\
        );

    \I__17540\ : Odrv4
    port map (
            O => \N__72597\,
            I => \c0.n14_adj_4619\
        );

    \I__17539\ : CascadeMux
    port map (
            O => \N__72594\,
            I => \N__72591\
        );

    \I__17538\ : InMux
    port map (
            O => \N__72591\,
            I => \N__72588\
        );

    \I__17537\ : LocalMux
    port map (
            O => \N__72588\,
            I => \N__72582\
        );

    \I__17536\ : InMux
    port map (
            O => \N__72587\,
            I => \N__72578\
        );

    \I__17535\ : CascadeMux
    port map (
            O => \N__72586\,
            I => \N__72574\
        );

    \I__17534\ : CascadeMux
    port map (
            O => \N__72585\,
            I => \N__72571\
        );

    \I__17533\ : Span4Mux_v
    port map (
            O => \N__72582\,
            I => \N__72567\
        );

    \I__17532\ : InMux
    port map (
            O => \N__72581\,
            I => \N__72564\
        );

    \I__17531\ : LocalMux
    port map (
            O => \N__72578\,
            I => \N__72560\
        );

    \I__17530\ : InMux
    port map (
            O => \N__72577\,
            I => \N__72556\
        );

    \I__17529\ : InMux
    port map (
            O => \N__72574\,
            I => \N__72553\
        );

    \I__17528\ : InMux
    port map (
            O => \N__72571\,
            I => \N__72550\
        );

    \I__17527\ : InMux
    port map (
            O => \N__72570\,
            I => \N__72547\
        );

    \I__17526\ : Span4Mux_v
    port map (
            O => \N__72567\,
            I => \N__72542\
        );

    \I__17525\ : LocalMux
    port map (
            O => \N__72564\,
            I => \N__72542\
        );

    \I__17524\ : InMux
    port map (
            O => \N__72563\,
            I => \N__72539\
        );

    \I__17523\ : Span4Mux_v
    port map (
            O => \N__72560\,
            I => \N__72536\
        );

    \I__17522\ : InMux
    port map (
            O => \N__72559\,
            I => \N__72533\
        );

    \I__17521\ : LocalMux
    port map (
            O => \N__72556\,
            I => \N__72530\
        );

    \I__17520\ : LocalMux
    port map (
            O => \N__72553\,
            I => \N__72521\
        );

    \I__17519\ : LocalMux
    port map (
            O => \N__72550\,
            I => \N__72521\
        );

    \I__17518\ : LocalMux
    port map (
            O => \N__72547\,
            I => \N__72521\
        );

    \I__17517\ : Span4Mux_v
    port map (
            O => \N__72542\,
            I => \N__72518\
        );

    \I__17516\ : LocalMux
    port map (
            O => \N__72539\,
            I => \N__72515\
        );

    \I__17515\ : Span4Mux_v
    port map (
            O => \N__72536\,
            I => \N__72508\
        );

    \I__17514\ : LocalMux
    port map (
            O => \N__72533\,
            I => \N__72508\
        );

    \I__17513\ : Span4Mux_h
    port map (
            O => \N__72530\,
            I => \N__72508\
        );

    \I__17512\ : InMux
    port map (
            O => \N__72529\,
            I => \N__72503\
        );

    \I__17511\ : InMux
    port map (
            O => \N__72528\,
            I => \N__72503\
        );

    \I__17510\ : Span4Mux_h
    port map (
            O => \N__72521\,
            I => \N__72500\
        );

    \I__17509\ : Odrv4
    port map (
            O => \N__72518\,
            I => \c0.data_in_frame_2_1\
        );

    \I__17508\ : Odrv4
    port map (
            O => \N__72515\,
            I => \c0.data_in_frame_2_1\
        );

    \I__17507\ : Odrv4
    port map (
            O => \N__72508\,
            I => \c0.data_in_frame_2_1\
        );

    \I__17506\ : LocalMux
    port map (
            O => \N__72503\,
            I => \c0.data_in_frame_2_1\
        );

    \I__17505\ : Odrv4
    port map (
            O => \N__72500\,
            I => \c0.data_in_frame_2_1\
        );

    \I__17504\ : InMux
    port map (
            O => \N__72489\,
            I => \N__72486\
        );

    \I__17503\ : LocalMux
    port map (
            O => \N__72486\,
            I => \c0.n22288\
        );

    \I__17502\ : CascadeMux
    port map (
            O => \N__72483\,
            I => \N__72479\
        );

    \I__17501\ : CascadeMux
    port map (
            O => \N__72482\,
            I => \N__72476\
        );

    \I__17500\ : InMux
    port map (
            O => \N__72479\,
            I => \N__72473\
        );

    \I__17499\ : InMux
    port map (
            O => \N__72476\,
            I => \N__72469\
        );

    \I__17498\ : LocalMux
    port map (
            O => \N__72473\,
            I => \N__72465\
        );

    \I__17497\ : InMux
    port map (
            O => \N__72472\,
            I => \N__72460\
        );

    \I__17496\ : LocalMux
    port map (
            O => \N__72469\,
            I => \N__72457\
        );

    \I__17495\ : InMux
    port map (
            O => \N__72468\,
            I => \N__72454\
        );

    \I__17494\ : Span4Mux_h
    port map (
            O => \N__72465\,
            I => \N__72451\
        );

    \I__17493\ : CascadeMux
    port map (
            O => \N__72464\,
            I => \N__72448\
        );

    \I__17492\ : InMux
    port map (
            O => \N__72463\,
            I => \N__72445\
        );

    \I__17491\ : LocalMux
    port map (
            O => \N__72460\,
            I => \N__72442\
        );

    \I__17490\ : Span4Mux_v
    port map (
            O => \N__72457\,
            I => \N__72439\
        );

    \I__17489\ : LocalMux
    port map (
            O => \N__72454\,
            I => \N__72436\
        );

    \I__17488\ : Span4Mux_h
    port map (
            O => \N__72451\,
            I => \N__72433\
        );

    \I__17487\ : InMux
    port map (
            O => \N__72448\,
            I => \N__72430\
        );

    \I__17486\ : LocalMux
    port map (
            O => \N__72445\,
            I => \c0.data_in_frame_13_2\
        );

    \I__17485\ : Odrv4
    port map (
            O => \N__72442\,
            I => \c0.data_in_frame_13_2\
        );

    \I__17484\ : Odrv4
    port map (
            O => \N__72439\,
            I => \c0.data_in_frame_13_2\
        );

    \I__17483\ : Odrv4
    port map (
            O => \N__72436\,
            I => \c0.data_in_frame_13_2\
        );

    \I__17482\ : Odrv4
    port map (
            O => \N__72433\,
            I => \c0.data_in_frame_13_2\
        );

    \I__17481\ : LocalMux
    port map (
            O => \N__72430\,
            I => \c0.data_in_frame_13_2\
        );

    \I__17480\ : CascadeMux
    port map (
            O => \N__72417\,
            I => \c0.n22288_cascade_\
        );

    \I__17479\ : CascadeMux
    port map (
            O => \N__72414\,
            I => \N__72410\
        );

    \I__17478\ : InMux
    port map (
            O => \N__72413\,
            I => \N__72407\
        );

    \I__17477\ : InMux
    port map (
            O => \N__72410\,
            I => \N__72404\
        );

    \I__17476\ : LocalMux
    port map (
            O => \N__72407\,
            I => \N__72401\
        );

    \I__17475\ : LocalMux
    port map (
            O => \N__72404\,
            I => \N__72398\
        );

    \I__17474\ : Span4Mux_h
    port map (
            O => \N__72401\,
            I => \N__72393\
        );

    \I__17473\ : Span4Mux_v
    port map (
            O => \N__72398\,
            I => \N__72390\
        );

    \I__17472\ : InMux
    port map (
            O => \N__72397\,
            I => \N__72387\
        );

    \I__17471\ : InMux
    port map (
            O => \N__72396\,
            I => \N__72384\
        );

    \I__17470\ : Span4Mux_v
    port map (
            O => \N__72393\,
            I => \N__72377\
        );

    \I__17469\ : Span4Mux_h
    port map (
            O => \N__72390\,
            I => \N__72377\
        );

    \I__17468\ : LocalMux
    port map (
            O => \N__72387\,
            I => \N__72377\
        );

    \I__17467\ : LocalMux
    port map (
            O => \N__72384\,
            I => \c0.n5807\
        );

    \I__17466\ : Odrv4
    port map (
            O => \N__72377\,
            I => \c0.n5807\
        );

    \I__17465\ : InMux
    port map (
            O => \N__72372\,
            I => \N__72367\
        );

    \I__17464\ : InMux
    port map (
            O => \N__72371\,
            I => \N__72361\
        );

    \I__17463\ : InMux
    port map (
            O => \N__72370\,
            I => \N__72361\
        );

    \I__17462\ : LocalMux
    port map (
            O => \N__72367\,
            I => \N__72357\
        );

    \I__17461\ : InMux
    port map (
            O => \N__72366\,
            I => \N__72354\
        );

    \I__17460\ : LocalMux
    port map (
            O => \N__72361\,
            I => \N__72351\
        );

    \I__17459\ : InMux
    port map (
            O => \N__72360\,
            I => \N__72348\
        );

    \I__17458\ : Span4Mux_v
    port map (
            O => \N__72357\,
            I => \N__72342\
        );

    \I__17457\ : LocalMux
    port map (
            O => \N__72354\,
            I => \N__72342\
        );

    \I__17456\ : Span4Mux_v
    port map (
            O => \N__72351\,
            I => \N__72337\
        );

    \I__17455\ : LocalMux
    port map (
            O => \N__72348\,
            I => \N__72337\
        );

    \I__17454\ : InMux
    port map (
            O => \N__72347\,
            I => \N__72334\
        );

    \I__17453\ : Span4Mux_v
    port map (
            O => \N__72342\,
            I => \N__72329\
        );

    \I__17452\ : Span4Mux_h
    port map (
            O => \N__72337\,
            I => \N__72329\
        );

    \I__17451\ : LocalMux
    port map (
            O => \N__72334\,
            I => \N__72326\
        );

    \I__17450\ : Odrv4
    port map (
            O => \N__72329\,
            I => \c0.n14160\
        );

    \I__17449\ : Odrv12
    port map (
            O => \N__72326\,
            I => \c0.n14160\
        );

    \I__17448\ : InMux
    port map (
            O => \N__72321\,
            I => \N__72315\
        );

    \I__17447\ : InMux
    port map (
            O => \N__72320\,
            I => \N__72310\
        );

    \I__17446\ : InMux
    port map (
            O => \N__72319\,
            I => \N__72310\
        );

    \I__17445\ : InMux
    port map (
            O => \N__72318\,
            I => \N__72306\
        );

    \I__17444\ : LocalMux
    port map (
            O => \N__72315\,
            I => \N__72303\
        );

    \I__17443\ : LocalMux
    port map (
            O => \N__72310\,
            I => \N__72300\
        );

    \I__17442\ : CascadeMux
    port map (
            O => \N__72309\,
            I => \N__72296\
        );

    \I__17441\ : LocalMux
    port map (
            O => \N__72306\,
            I => \N__72293\
        );

    \I__17440\ : Span4Mux_v
    port map (
            O => \N__72303\,
            I => \N__72288\
        );

    \I__17439\ : Span4Mux_h
    port map (
            O => \N__72300\,
            I => \N__72288\
        );

    \I__17438\ : InMux
    port map (
            O => \N__72299\,
            I => \N__72285\
        );

    \I__17437\ : InMux
    port map (
            O => \N__72296\,
            I => \N__72280\
        );

    \I__17436\ : Span4Mux_h
    port map (
            O => \N__72293\,
            I => \N__72277\
        );

    \I__17435\ : Span4Mux_v
    port map (
            O => \N__72288\,
            I => \N__72274\
        );

    \I__17434\ : LocalMux
    port map (
            O => \N__72285\,
            I => \N__72271\
        );

    \I__17433\ : InMux
    port map (
            O => \N__72284\,
            I => \N__72268\
        );

    \I__17432\ : InMux
    port map (
            O => \N__72283\,
            I => \N__72265\
        );

    \I__17431\ : LocalMux
    port map (
            O => \N__72280\,
            I => \c0.data_in_frame_8_3\
        );

    \I__17430\ : Odrv4
    port map (
            O => \N__72277\,
            I => \c0.data_in_frame_8_3\
        );

    \I__17429\ : Odrv4
    port map (
            O => \N__72274\,
            I => \c0.data_in_frame_8_3\
        );

    \I__17428\ : Odrv12
    port map (
            O => \N__72271\,
            I => \c0.data_in_frame_8_3\
        );

    \I__17427\ : LocalMux
    port map (
            O => \N__72268\,
            I => \c0.data_in_frame_8_3\
        );

    \I__17426\ : LocalMux
    port map (
            O => \N__72265\,
            I => \c0.data_in_frame_8_3\
        );

    \I__17425\ : InMux
    port map (
            O => \N__72252\,
            I => \N__72246\
        );

    \I__17424\ : InMux
    port map (
            O => \N__72251\,
            I => \N__72246\
        );

    \I__17423\ : LocalMux
    port map (
            O => \N__72246\,
            I => \N__72243\
        );

    \I__17422\ : Span4Mux_v
    port map (
            O => \N__72243\,
            I => \N__72239\
        );

    \I__17421\ : InMux
    port map (
            O => \N__72242\,
            I => \N__72234\
        );

    \I__17420\ : Span4Mux_h
    port map (
            O => \N__72239\,
            I => \N__72231\
        );

    \I__17419\ : InMux
    port map (
            O => \N__72238\,
            I => \N__72226\
        );

    \I__17418\ : InMux
    port map (
            O => \N__72237\,
            I => \N__72226\
        );

    \I__17417\ : LocalMux
    port map (
            O => \N__72234\,
            I => \c0.data_in_frame_17_4\
        );

    \I__17416\ : Odrv4
    port map (
            O => \N__72231\,
            I => \c0.data_in_frame_17_4\
        );

    \I__17415\ : LocalMux
    port map (
            O => \N__72226\,
            I => \c0.data_in_frame_17_4\
        );

    \I__17414\ : InMux
    port map (
            O => \N__72219\,
            I => \N__72216\
        );

    \I__17413\ : LocalMux
    port map (
            O => \N__72216\,
            I => \N__72211\
        );

    \I__17412\ : CascadeMux
    port map (
            O => \N__72215\,
            I => \N__72207\
        );

    \I__17411\ : CascadeMux
    port map (
            O => \N__72214\,
            I => \N__72203\
        );

    \I__17410\ : Span4Mux_v
    port map (
            O => \N__72211\,
            I => \N__72200\
        );

    \I__17409\ : InMux
    port map (
            O => \N__72210\,
            I => \N__72197\
        );

    \I__17408\ : InMux
    port map (
            O => \N__72207\,
            I => \N__72192\
        );

    \I__17407\ : InMux
    port map (
            O => \N__72206\,
            I => \N__72187\
        );

    \I__17406\ : InMux
    port map (
            O => \N__72203\,
            I => \N__72187\
        );

    \I__17405\ : Span4Mux_h
    port map (
            O => \N__72200\,
            I => \N__72182\
        );

    \I__17404\ : LocalMux
    port map (
            O => \N__72197\,
            I => \N__72182\
        );

    \I__17403\ : InMux
    port map (
            O => \N__72196\,
            I => \N__72179\
        );

    \I__17402\ : InMux
    port map (
            O => \N__72195\,
            I => \N__72176\
        );

    \I__17401\ : LocalMux
    port map (
            O => \N__72192\,
            I => \c0.data_in_frame_13_3\
        );

    \I__17400\ : LocalMux
    port map (
            O => \N__72187\,
            I => \c0.data_in_frame_13_3\
        );

    \I__17399\ : Odrv4
    port map (
            O => \N__72182\,
            I => \c0.data_in_frame_13_3\
        );

    \I__17398\ : LocalMux
    port map (
            O => \N__72179\,
            I => \c0.data_in_frame_13_3\
        );

    \I__17397\ : LocalMux
    port map (
            O => \N__72176\,
            I => \c0.data_in_frame_13_3\
        );

    \I__17396\ : InMux
    port map (
            O => \N__72165\,
            I => \N__72162\
        );

    \I__17395\ : LocalMux
    port map (
            O => \N__72162\,
            I => \N__72158\
        );

    \I__17394\ : InMux
    port map (
            O => \N__72161\,
            I => \N__72155\
        );

    \I__17393\ : Span4Mux_h
    port map (
            O => \N__72158\,
            I => \N__72149\
        );

    \I__17392\ : LocalMux
    port map (
            O => \N__72155\,
            I => \N__72146\
        );

    \I__17391\ : InMux
    port map (
            O => \N__72154\,
            I => \N__72143\
        );

    \I__17390\ : InMux
    port map (
            O => \N__72153\,
            I => \N__72138\
        );

    \I__17389\ : InMux
    port map (
            O => \N__72152\,
            I => \N__72138\
        );

    \I__17388\ : Span4Mux_h
    port map (
            O => \N__72149\,
            I => \N__72135\
        );

    \I__17387\ : Span12Mux_v
    port map (
            O => \N__72146\,
            I => \N__72130\
        );

    \I__17386\ : LocalMux
    port map (
            O => \N__72143\,
            I => \N__72130\
        );

    \I__17385\ : LocalMux
    port map (
            O => \N__72138\,
            I => \c0.n22319\
        );

    \I__17384\ : Odrv4
    port map (
            O => \N__72135\,
            I => \c0.n22319\
        );

    \I__17383\ : Odrv12
    port map (
            O => \N__72130\,
            I => \c0.n22319\
        );

    \I__17382\ : InMux
    port map (
            O => \N__72123\,
            I => \N__72120\
        );

    \I__17381\ : LocalMux
    port map (
            O => \N__72120\,
            I => \N__72117\
        );

    \I__17380\ : Span4Mux_h
    port map (
            O => \N__72117\,
            I => \N__72114\
        );

    \I__17379\ : Odrv4
    port map (
            O => \N__72114\,
            I => \c0.n4_adj_4586\
        );

    \I__17378\ : InMux
    port map (
            O => \N__72111\,
            I => \N__72107\
        );

    \I__17377\ : CascadeMux
    port map (
            O => \N__72110\,
            I => \N__72104\
        );

    \I__17376\ : LocalMux
    port map (
            O => \N__72107\,
            I => \N__72100\
        );

    \I__17375\ : InMux
    port map (
            O => \N__72104\,
            I => \N__72095\
        );

    \I__17374\ : InMux
    port map (
            O => \N__72103\,
            I => \N__72095\
        );

    \I__17373\ : Odrv4
    port map (
            O => \N__72100\,
            I => \c0.data_in_frame_16_0\
        );

    \I__17372\ : LocalMux
    port map (
            O => \N__72095\,
            I => \c0.data_in_frame_16_0\
        );

    \I__17371\ : InMux
    port map (
            O => \N__72090\,
            I => \N__72085\
        );

    \I__17370\ : InMux
    port map (
            O => \N__72089\,
            I => \N__72082\
        );

    \I__17369\ : CascadeMux
    port map (
            O => \N__72088\,
            I => \N__72079\
        );

    \I__17368\ : LocalMux
    port map (
            O => \N__72085\,
            I => \N__72075\
        );

    \I__17367\ : LocalMux
    port map (
            O => \N__72082\,
            I => \N__72072\
        );

    \I__17366\ : InMux
    port map (
            O => \N__72079\,
            I => \N__72067\
        );

    \I__17365\ : InMux
    port map (
            O => \N__72078\,
            I => \N__72067\
        );

    \I__17364\ : Odrv12
    port map (
            O => \N__72075\,
            I => \c0.data_in_frame_13_6\
        );

    \I__17363\ : Odrv4
    port map (
            O => \N__72072\,
            I => \c0.data_in_frame_13_6\
        );

    \I__17362\ : LocalMux
    port map (
            O => \N__72067\,
            I => \c0.data_in_frame_13_6\
        );

    \I__17361\ : CascadeMux
    port map (
            O => \N__72060\,
            I => \N__72057\
        );

    \I__17360\ : InMux
    port map (
            O => \N__72057\,
            I => \N__72054\
        );

    \I__17359\ : LocalMux
    port map (
            O => \N__72054\,
            I => \N__72051\
        );

    \I__17358\ : Span12Mux_s11_h
    port map (
            O => \N__72051\,
            I => \N__72046\
        );

    \I__17357\ : InMux
    port map (
            O => \N__72050\,
            I => \N__72041\
        );

    \I__17356\ : InMux
    port map (
            O => \N__72049\,
            I => \N__72041\
        );

    \I__17355\ : Odrv12
    port map (
            O => \N__72046\,
            I => \c0.data_in_frame_18_1\
        );

    \I__17354\ : LocalMux
    port map (
            O => \N__72041\,
            I => \c0.data_in_frame_18_1\
        );

    \I__17353\ : InMux
    port map (
            O => \N__72036\,
            I => \N__72033\
        );

    \I__17352\ : LocalMux
    port map (
            O => \N__72033\,
            I => \N__72029\
        );

    \I__17351\ : InMux
    port map (
            O => \N__72032\,
            I => \N__72026\
        );

    \I__17350\ : Odrv4
    port map (
            O => \N__72029\,
            I => \c0.n14081\
        );

    \I__17349\ : LocalMux
    port map (
            O => \N__72026\,
            I => \c0.n14081\
        );

    \I__17348\ : InMux
    port map (
            O => \N__72021\,
            I => \N__72018\
        );

    \I__17347\ : LocalMux
    port map (
            O => \N__72018\,
            I => \N__72014\
        );

    \I__17346\ : InMux
    port map (
            O => \N__72017\,
            I => \N__72011\
        );

    \I__17345\ : Odrv12
    port map (
            O => \N__72014\,
            I => \c0.n10_adj_4250\
        );

    \I__17344\ : LocalMux
    port map (
            O => \N__72011\,
            I => \c0.n10_adj_4250\
        );

    \I__17343\ : CascadeMux
    port map (
            O => \N__72006\,
            I => \N__72003\
        );

    \I__17342\ : InMux
    port map (
            O => \N__72003\,
            I => \N__71998\
        );

    \I__17341\ : InMux
    port map (
            O => \N__72002\,
            I => \N__71995\
        );

    \I__17340\ : InMux
    port map (
            O => \N__72001\,
            I => \N__71992\
        );

    \I__17339\ : LocalMux
    port map (
            O => \N__71998\,
            I => \N__71989\
        );

    \I__17338\ : LocalMux
    port map (
            O => \N__71995\,
            I => \N__71981\
        );

    \I__17337\ : LocalMux
    port map (
            O => \N__71992\,
            I => \N__71981\
        );

    \I__17336\ : Span4Mux_v
    port map (
            O => \N__71989\,
            I => \N__71981\
        );

    \I__17335\ : InMux
    port map (
            O => \N__71988\,
            I => \N__71978\
        );

    \I__17334\ : Span4Mux_h
    port map (
            O => \N__71981\,
            I => \N__71975\
        );

    \I__17333\ : LocalMux
    port map (
            O => \N__71978\,
            I => \c0.data_in_frame_16_4\
        );

    \I__17332\ : Odrv4
    port map (
            O => \N__71975\,
            I => \c0.data_in_frame_16_4\
        );

    \I__17331\ : CascadeMux
    port map (
            O => \N__71970\,
            I => \N__71963\
        );

    \I__17330\ : CascadeMux
    port map (
            O => \N__71969\,
            I => \N__71960\
        );

    \I__17329\ : InMux
    port map (
            O => \N__71968\,
            I => \N__71954\
        );

    \I__17328\ : CascadeMux
    port map (
            O => \N__71967\,
            I => \N__71950\
        );

    \I__17327\ : CascadeMux
    port map (
            O => \N__71966\,
            I => \N__71947\
        );

    \I__17326\ : InMux
    port map (
            O => \N__71963\,
            I => \N__71940\
        );

    \I__17325\ : InMux
    port map (
            O => \N__71960\,
            I => \N__71931\
        );

    \I__17324\ : InMux
    port map (
            O => \N__71959\,
            I => \N__71931\
        );

    \I__17323\ : InMux
    port map (
            O => \N__71958\,
            I => \N__71928\
        );

    \I__17322\ : InMux
    port map (
            O => \N__71957\,
            I => \N__71925\
        );

    \I__17321\ : LocalMux
    port map (
            O => \N__71954\,
            I => \N__71922\
        );

    \I__17320\ : InMux
    port map (
            O => \N__71953\,
            I => \N__71918\
        );

    \I__17319\ : InMux
    port map (
            O => \N__71950\,
            I => \N__71910\
        );

    \I__17318\ : InMux
    port map (
            O => \N__71947\,
            I => \N__71907\
        );

    \I__17317\ : CascadeMux
    port map (
            O => \N__71946\,
            I => \N__71903\
        );

    \I__17316\ : InMux
    port map (
            O => \N__71945\,
            I => \N__71897\
        );

    \I__17315\ : InMux
    port map (
            O => \N__71944\,
            I => \N__71897\
        );

    \I__17314\ : InMux
    port map (
            O => \N__71943\,
            I => \N__71894\
        );

    \I__17313\ : LocalMux
    port map (
            O => \N__71940\,
            I => \N__71891\
        );

    \I__17312\ : InMux
    port map (
            O => \N__71939\,
            I => \N__71888\
        );

    \I__17311\ : CascadeMux
    port map (
            O => \N__71938\,
            I => \N__71884\
        );

    \I__17310\ : InMux
    port map (
            O => \N__71937\,
            I => \N__71879\
        );

    \I__17309\ : InMux
    port map (
            O => \N__71936\,
            I => \N__71879\
        );

    \I__17308\ : LocalMux
    port map (
            O => \N__71931\,
            I => \N__71876\
        );

    \I__17307\ : LocalMux
    port map (
            O => \N__71928\,
            I => \N__71872\
        );

    \I__17306\ : LocalMux
    port map (
            O => \N__71925\,
            I => \N__71867\
        );

    \I__17305\ : Span4Mux_h
    port map (
            O => \N__71922\,
            I => \N__71867\
        );

    \I__17304\ : CascadeMux
    port map (
            O => \N__71921\,
            I => \N__71863\
        );

    \I__17303\ : LocalMux
    port map (
            O => \N__71918\,
            I => \N__71860\
        );

    \I__17302\ : InMux
    port map (
            O => \N__71917\,
            I => \N__71855\
        );

    \I__17301\ : InMux
    port map (
            O => \N__71916\,
            I => \N__71855\
        );

    \I__17300\ : InMux
    port map (
            O => \N__71915\,
            I => \N__71850\
        );

    \I__17299\ : InMux
    port map (
            O => \N__71914\,
            I => \N__71850\
        );

    \I__17298\ : InMux
    port map (
            O => \N__71913\,
            I => \N__71847\
        );

    \I__17297\ : LocalMux
    port map (
            O => \N__71910\,
            I => \N__71842\
        );

    \I__17296\ : LocalMux
    port map (
            O => \N__71907\,
            I => \N__71842\
        );

    \I__17295\ : InMux
    port map (
            O => \N__71906\,
            I => \N__71837\
        );

    \I__17294\ : InMux
    port map (
            O => \N__71903\,
            I => \N__71837\
        );

    \I__17293\ : InMux
    port map (
            O => \N__71902\,
            I => \N__71834\
        );

    \I__17292\ : LocalMux
    port map (
            O => \N__71897\,
            I => \N__71831\
        );

    \I__17291\ : LocalMux
    port map (
            O => \N__71894\,
            I => \N__71828\
        );

    \I__17290\ : Span4Mux_h
    port map (
            O => \N__71891\,
            I => \N__71825\
        );

    \I__17289\ : LocalMux
    port map (
            O => \N__71888\,
            I => \N__71822\
        );

    \I__17288\ : InMux
    port map (
            O => \N__71887\,
            I => \N__71817\
        );

    \I__17287\ : InMux
    port map (
            O => \N__71884\,
            I => \N__71817\
        );

    \I__17286\ : LocalMux
    port map (
            O => \N__71879\,
            I => \N__71811\
        );

    \I__17285\ : Span4Mux_v
    port map (
            O => \N__71876\,
            I => \N__71811\
        );

    \I__17284\ : InMux
    port map (
            O => \N__71875\,
            I => \N__71808\
        );

    \I__17283\ : Span4Mux_h
    port map (
            O => \N__71872\,
            I => \N__71805\
        );

    \I__17282\ : Sp12to4
    port map (
            O => \N__71867\,
            I => \N__71802\
        );

    \I__17281\ : InMux
    port map (
            O => \N__71866\,
            I => \N__71799\
        );

    \I__17280\ : InMux
    port map (
            O => \N__71863\,
            I => \N__71796\
        );

    \I__17279\ : Span4Mux_v
    port map (
            O => \N__71860\,
            I => \N__71793\
        );

    \I__17278\ : LocalMux
    port map (
            O => \N__71855\,
            I => \N__71790\
        );

    \I__17277\ : LocalMux
    port map (
            O => \N__71850\,
            I => \N__71787\
        );

    \I__17276\ : LocalMux
    port map (
            O => \N__71847\,
            I => \N__71782\
        );

    \I__17275\ : Span4Mux_h
    port map (
            O => \N__71842\,
            I => \N__71782\
        );

    \I__17274\ : LocalMux
    port map (
            O => \N__71837\,
            I => \N__71778\
        );

    \I__17273\ : LocalMux
    port map (
            O => \N__71834\,
            I => \N__71773\
        );

    \I__17272\ : Span4Mux_v
    port map (
            O => \N__71831\,
            I => \N__71773\
        );

    \I__17271\ : Span4Mux_h
    port map (
            O => \N__71828\,
            I => \N__71768\
        );

    \I__17270\ : Span4Mux_v
    port map (
            O => \N__71825\,
            I => \N__71768\
        );

    \I__17269\ : Span4Mux_h
    port map (
            O => \N__71822\,
            I => \N__71763\
        );

    \I__17268\ : LocalMux
    port map (
            O => \N__71817\,
            I => \N__71763\
        );

    \I__17267\ : InMux
    port map (
            O => \N__71816\,
            I => \N__71758\
        );

    \I__17266\ : Span4Mux_v
    port map (
            O => \N__71811\,
            I => \N__71753\
        );

    \I__17265\ : LocalMux
    port map (
            O => \N__71808\,
            I => \N__71753\
        );

    \I__17264\ : Sp12to4
    port map (
            O => \N__71805\,
            I => \N__71744\
        );

    \I__17263\ : Span12Mux_v
    port map (
            O => \N__71802\,
            I => \N__71744\
        );

    \I__17262\ : LocalMux
    port map (
            O => \N__71799\,
            I => \N__71744\
        );

    \I__17261\ : LocalMux
    port map (
            O => \N__71796\,
            I => \N__71744\
        );

    \I__17260\ : Span4Mux_v
    port map (
            O => \N__71793\,
            I => \N__71741\
        );

    \I__17259\ : Span4Mux_h
    port map (
            O => \N__71790\,
            I => \N__71734\
        );

    \I__17258\ : Span4Mux_v
    port map (
            O => \N__71787\,
            I => \N__71734\
        );

    \I__17257\ : Span4Mux_v
    port map (
            O => \N__71782\,
            I => \N__71734\
        );

    \I__17256\ : InMux
    port map (
            O => \N__71781\,
            I => \N__71731\
        );

    \I__17255\ : Span4Mux_v
    port map (
            O => \N__71778\,
            I => \N__71726\
        );

    \I__17254\ : Span4Mux_v
    port map (
            O => \N__71773\,
            I => \N__71726\
        );

    \I__17253\ : Sp12to4
    port map (
            O => \N__71768\,
            I => \N__71723\
        );

    \I__17252\ : Sp12to4
    port map (
            O => \N__71763\,
            I => \N__71720\
        );

    \I__17251\ : InMux
    port map (
            O => \N__71762\,
            I => \N__71715\
        );

    \I__17250\ : InMux
    port map (
            O => \N__71761\,
            I => \N__71715\
        );

    \I__17249\ : LocalMux
    port map (
            O => \N__71758\,
            I => \N__71712\
        );

    \I__17248\ : Span4Mux_h
    port map (
            O => \N__71753\,
            I => \N__71709\
        );

    \I__17247\ : Span12Mux_v
    port map (
            O => \N__71744\,
            I => \N__71706\
        );

    \I__17246\ : Span4Mux_h
    port map (
            O => \N__71741\,
            I => \N__71701\
        );

    \I__17245\ : Span4Mux_v
    port map (
            O => \N__71734\,
            I => \N__71701\
        );

    \I__17244\ : LocalMux
    port map (
            O => \N__71731\,
            I => \N__71692\
        );

    \I__17243\ : Sp12to4
    port map (
            O => \N__71726\,
            I => \N__71692\
        );

    \I__17242\ : Span12Mux_v
    port map (
            O => \N__71723\,
            I => \N__71692\
        );

    \I__17241\ : Span12Mux_v
    port map (
            O => \N__71720\,
            I => \N__71692\
        );

    \I__17240\ : LocalMux
    port map (
            O => \N__71715\,
            I => rx_data_4
        );

    \I__17239\ : Odrv4
    port map (
            O => \N__71712\,
            I => rx_data_4
        );

    \I__17238\ : Odrv4
    port map (
            O => \N__71709\,
            I => rx_data_4
        );

    \I__17237\ : Odrv12
    port map (
            O => \N__71706\,
            I => rx_data_4
        );

    \I__17236\ : Odrv4
    port map (
            O => \N__71701\,
            I => rx_data_4
        );

    \I__17235\ : Odrv12
    port map (
            O => \N__71692\,
            I => rx_data_4
        );

    \I__17234\ : CascadeMux
    port map (
            O => \N__71679\,
            I => \N__71676\
        );

    \I__17233\ : InMux
    port map (
            O => \N__71676\,
            I => \N__71670\
        );

    \I__17232\ : InMux
    port map (
            O => \N__71675\,
            I => \N__71667\
        );

    \I__17231\ : InMux
    port map (
            O => \N__71674\,
            I => \N__71662\
        );

    \I__17230\ : InMux
    port map (
            O => \N__71673\,
            I => \N__71662\
        );

    \I__17229\ : LocalMux
    port map (
            O => \N__71670\,
            I => \N__71659\
        );

    \I__17228\ : LocalMux
    port map (
            O => \N__71667\,
            I => \N__71656\
        );

    \I__17227\ : LocalMux
    port map (
            O => \N__71662\,
            I => \N__71653\
        );

    \I__17226\ : Odrv4
    port map (
            O => \N__71659\,
            I => \c0.data_in_frame_13_4\
        );

    \I__17225\ : Odrv4
    port map (
            O => \N__71656\,
            I => \c0.data_in_frame_13_4\
        );

    \I__17224\ : Odrv4
    port map (
            O => \N__71653\,
            I => \c0.data_in_frame_13_4\
        );

    \I__17223\ : InMux
    port map (
            O => \N__71646\,
            I => \N__71642\
        );

    \I__17222\ : InMux
    port map (
            O => \N__71645\,
            I => \N__71639\
        );

    \I__17221\ : LocalMux
    port map (
            O => \N__71642\,
            I => \N__71636\
        );

    \I__17220\ : LocalMux
    port map (
            O => \N__71639\,
            I => \N__71632\
        );

    \I__17219\ : Span4Mux_v
    port map (
            O => \N__71636\,
            I => \N__71628\
        );

    \I__17218\ : CascadeMux
    port map (
            O => \N__71635\,
            I => \N__71624\
        );

    \I__17217\ : Span4Mux_v
    port map (
            O => \N__71632\,
            I => \N__71621\
        );

    \I__17216\ : CascadeMux
    port map (
            O => \N__71631\,
            I => \N__71618\
        );

    \I__17215\ : Span4Mux_h
    port map (
            O => \N__71628\,
            I => \N__71615\
        );

    \I__17214\ : InMux
    port map (
            O => \N__71627\,
            I => \N__71612\
        );

    \I__17213\ : InMux
    port map (
            O => \N__71624\,
            I => \N__71609\
        );

    \I__17212\ : Span4Mux_h
    port map (
            O => \N__71621\,
            I => \N__71606\
        );

    \I__17211\ : InMux
    port map (
            O => \N__71618\,
            I => \N__71603\
        );

    \I__17210\ : Sp12to4
    port map (
            O => \N__71615\,
            I => \N__71598\
        );

    \I__17209\ : LocalMux
    port map (
            O => \N__71612\,
            I => \N__71598\
        );

    \I__17208\ : LocalMux
    port map (
            O => \N__71609\,
            I => \c0.data_in_frame_19_5\
        );

    \I__17207\ : Odrv4
    port map (
            O => \N__71606\,
            I => \c0.data_in_frame_19_5\
        );

    \I__17206\ : LocalMux
    port map (
            O => \N__71603\,
            I => \c0.data_in_frame_19_5\
        );

    \I__17205\ : Odrv12
    port map (
            O => \N__71598\,
            I => \c0.data_in_frame_19_5\
        );

    \I__17204\ : InMux
    port map (
            O => \N__71589\,
            I => \N__71585\
        );

    \I__17203\ : InMux
    port map (
            O => \N__71588\,
            I => \N__71582\
        );

    \I__17202\ : LocalMux
    port map (
            O => \N__71585\,
            I => \N__71579\
        );

    \I__17201\ : LocalMux
    port map (
            O => \N__71582\,
            I => \N__71576\
        );

    \I__17200\ : Span4Mux_h
    port map (
            O => \N__71579\,
            I => \N__71573\
        );

    \I__17199\ : Span4Mux_v
    port map (
            O => \N__71576\,
            I => \N__71569\
        );

    \I__17198\ : Span4Mux_h
    port map (
            O => \N__71573\,
            I => \N__71566\
        );

    \I__17197\ : InMux
    port map (
            O => \N__71572\,
            I => \N__71563\
        );

    \I__17196\ : Span4Mux_v
    port map (
            O => \N__71569\,
            I => \N__71560\
        );

    \I__17195\ : Odrv4
    port map (
            O => \N__71566\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__17194\ : LocalMux
    port map (
            O => \N__71563\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__17193\ : Odrv4
    port map (
            O => \N__71560\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__17192\ : InMux
    port map (
            O => \N__71553\,
            I => \N__71549\
        );

    \I__17191\ : InMux
    port map (
            O => \N__71552\,
            I => \N__71546\
        );

    \I__17190\ : LocalMux
    port map (
            O => \N__71549\,
            I => \N__71539\
        );

    \I__17189\ : LocalMux
    port map (
            O => \N__71546\,
            I => \N__71533\
        );

    \I__17188\ : InMux
    port map (
            O => \N__71545\,
            I => \N__71530\
        );

    \I__17187\ : InMux
    port map (
            O => \N__71544\,
            I => \N__71526\
        );

    \I__17186\ : InMux
    port map (
            O => \N__71543\,
            I => \N__71523\
        );

    \I__17185\ : InMux
    port map (
            O => \N__71542\,
            I => \N__71520\
        );

    \I__17184\ : Span4Mux_h
    port map (
            O => \N__71539\,
            I => \N__71516\
        );

    \I__17183\ : InMux
    port map (
            O => \N__71538\,
            I => \N__71513\
        );

    \I__17182\ : InMux
    port map (
            O => \N__71537\,
            I => \N__71510\
        );

    \I__17181\ : InMux
    port map (
            O => \N__71536\,
            I => \N__71507\
        );

    \I__17180\ : Span4Mux_v
    port map (
            O => \N__71533\,
            I => \N__71499\
        );

    \I__17179\ : LocalMux
    port map (
            O => \N__71530\,
            I => \N__71499\
        );

    \I__17178\ : InMux
    port map (
            O => \N__71529\,
            I => \N__71496\
        );

    \I__17177\ : LocalMux
    port map (
            O => \N__71526\,
            I => \N__71493\
        );

    \I__17176\ : LocalMux
    port map (
            O => \N__71523\,
            I => \N__71490\
        );

    \I__17175\ : LocalMux
    port map (
            O => \N__71520\,
            I => \N__71487\
        );

    \I__17174\ : InMux
    port map (
            O => \N__71519\,
            I => \N__71484\
        );

    \I__17173\ : Span4Mux_v
    port map (
            O => \N__71516\,
            I => \N__71477\
        );

    \I__17172\ : LocalMux
    port map (
            O => \N__71513\,
            I => \N__71477\
        );

    \I__17171\ : LocalMux
    port map (
            O => \N__71510\,
            I => \N__71474\
        );

    \I__17170\ : LocalMux
    port map (
            O => \N__71507\,
            I => \N__71468\
        );

    \I__17169\ : InMux
    port map (
            O => \N__71506\,
            I => \N__71465\
        );

    \I__17168\ : InMux
    port map (
            O => \N__71505\,
            I => \N__71462\
        );

    \I__17167\ : InMux
    port map (
            O => \N__71504\,
            I => \N__71459\
        );

    \I__17166\ : Span4Mux_h
    port map (
            O => \N__71499\,
            I => \N__71451\
        );

    \I__17165\ : LocalMux
    port map (
            O => \N__71496\,
            I => \N__71448\
        );

    \I__17164\ : Span4Mux_h
    port map (
            O => \N__71493\,
            I => \N__71445\
        );

    \I__17163\ : Span4Mux_v
    port map (
            O => \N__71490\,
            I => \N__71442\
        );

    \I__17162\ : Span4Mux_v
    port map (
            O => \N__71487\,
            I => \N__71437\
        );

    \I__17161\ : LocalMux
    port map (
            O => \N__71484\,
            I => \N__71437\
        );

    \I__17160\ : InMux
    port map (
            O => \N__71483\,
            I => \N__71432\
        );

    \I__17159\ : InMux
    port map (
            O => \N__71482\,
            I => \N__71432\
        );

    \I__17158\ : Span4Mux_v
    port map (
            O => \N__71477\,
            I => \N__71429\
        );

    \I__17157\ : Span4Mux_v
    port map (
            O => \N__71474\,
            I => \N__71425\
        );

    \I__17156\ : InMux
    port map (
            O => \N__71473\,
            I => \N__71418\
        );

    \I__17155\ : InMux
    port map (
            O => \N__71472\,
            I => \N__71418\
        );

    \I__17154\ : InMux
    port map (
            O => \N__71471\,
            I => \N__71418\
        );

    \I__17153\ : Span4Mux_h
    port map (
            O => \N__71468\,
            I => \N__71409\
        );

    \I__17152\ : LocalMux
    port map (
            O => \N__71465\,
            I => \N__71409\
        );

    \I__17151\ : LocalMux
    port map (
            O => \N__71462\,
            I => \N__71409\
        );

    \I__17150\ : LocalMux
    port map (
            O => \N__71459\,
            I => \N__71409\
        );

    \I__17149\ : InMux
    port map (
            O => \N__71458\,
            I => \N__71406\
        );

    \I__17148\ : InMux
    port map (
            O => \N__71457\,
            I => \N__71403\
        );

    \I__17147\ : InMux
    port map (
            O => \N__71456\,
            I => \N__71398\
        );

    \I__17146\ : InMux
    port map (
            O => \N__71455\,
            I => \N__71398\
        );

    \I__17145\ : InMux
    port map (
            O => \N__71454\,
            I => \N__71395\
        );

    \I__17144\ : Sp12to4
    port map (
            O => \N__71451\,
            I => \N__71391\
        );

    \I__17143\ : Span12Mux_s11_h
    port map (
            O => \N__71448\,
            I => \N__71388\
        );

    \I__17142\ : Span4Mux_h
    port map (
            O => \N__71445\,
            I => \N__71379\
        );

    \I__17141\ : Span4Mux_h
    port map (
            O => \N__71442\,
            I => \N__71379\
        );

    \I__17140\ : Span4Mux_v
    port map (
            O => \N__71437\,
            I => \N__71379\
        );

    \I__17139\ : LocalMux
    port map (
            O => \N__71432\,
            I => \N__71379\
        );

    \I__17138\ : Span4Mux_v
    port map (
            O => \N__71429\,
            I => \N__71376\
        );

    \I__17137\ : InMux
    port map (
            O => \N__71428\,
            I => \N__71373\
        );

    \I__17136\ : Span4Mux_v
    port map (
            O => \N__71425\,
            I => \N__71369\
        );

    \I__17135\ : LocalMux
    port map (
            O => \N__71418\,
            I => \N__71366\
        );

    \I__17134\ : Span4Mux_v
    port map (
            O => \N__71409\,
            I => \N__71355\
        );

    \I__17133\ : LocalMux
    port map (
            O => \N__71406\,
            I => \N__71355\
        );

    \I__17132\ : LocalMux
    port map (
            O => \N__71403\,
            I => \N__71355\
        );

    \I__17131\ : LocalMux
    port map (
            O => \N__71398\,
            I => \N__71355\
        );

    \I__17130\ : LocalMux
    port map (
            O => \N__71395\,
            I => \N__71355\
        );

    \I__17129\ : InMux
    port map (
            O => \N__71394\,
            I => \N__71352\
        );

    \I__17128\ : Span12Mux_v
    port map (
            O => \N__71391\,
            I => \N__71344\
        );

    \I__17127\ : Span12Mux_v
    port map (
            O => \N__71388\,
            I => \N__71341\
        );

    \I__17126\ : Span4Mux_v
    port map (
            O => \N__71379\,
            I => \N__71338\
        );

    \I__17125\ : Span4Mux_v
    port map (
            O => \N__71376\,
            I => \N__71333\
        );

    \I__17124\ : LocalMux
    port map (
            O => \N__71373\,
            I => \N__71333\
        );

    \I__17123\ : InMux
    port map (
            O => \N__71372\,
            I => \N__71330\
        );

    \I__17122\ : Span4Mux_h
    port map (
            O => \N__71369\,
            I => \N__71321\
        );

    \I__17121\ : Span4Mux_v
    port map (
            O => \N__71366\,
            I => \N__71321\
        );

    \I__17120\ : Span4Mux_v
    port map (
            O => \N__71355\,
            I => \N__71321\
        );

    \I__17119\ : LocalMux
    port map (
            O => \N__71352\,
            I => \N__71321\
        );

    \I__17118\ : InMux
    port map (
            O => \N__71351\,
            I => \N__71310\
        );

    \I__17117\ : InMux
    port map (
            O => \N__71350\,
            I => \N__71310\
        );

    \I__17116\ : InMux
    port map (
            O => \N__71349\,
            I => \N__71310\
        );

    \I__17115\ : InMux
    port map (
            O => \N__71348\,
            I => \N__71310\
        );

    \I__17114\ : InMux
    port map (
            O => \N__71347\,
            I => \N__71310\
        );

    \I__17113\ : Odrv12
    port map (
            O => \N__71344\,
            I => \c0.n2119\
        );

    \I__17112\ : Odrv12
    port map (
            O => \N__71341\,
            I => \c0.n2119\
        );

    \I__17111\ : Odrv4
    port map (
            O => \N__71338\,
            I => \c0.n2119\
        );

    \I__17110\ : Odrv4
    port map (
            O => \N__71333\,
            I => \c0.n2119\
        );

    \I__17109\ : LocalMux
    port map (
            O => \N__71330\,
            I => \c0.n2119\
        );

    \I__17108\ : Odrv4
    port map (
            O => \N__71321\,
            I => \c0.n2119\
        );

    \I__17107\ : LocalMux
    port map (
            O => \N__71310\,
            I => \c0.n2119\
        );

    \I__17106\ : SRMux
    port map (
            O => \N__71295\,
            I => \N__71292\
        );

    \I__17105\ : LocalMux
    port map (
            O => \N__71292\,
            I => \N__71289\
        );

    \I__17104\ : Span4Mux_v
    port map (
            O => \N__71289\,
            I => \N__71286\
        );

    \I__17103\ : Span4Mux_h
    port map (
            O => \N__71286\,
            I => \N__71283\
        );

    \I__17102\ : Odrv4
    port map (
            O => \N__71283\,
            I => \c0.n3_adj_4400\
        );

    \I__17101\ : CascadeMux
    port map (
            O => \N__71280\,
            I => \N__71277\
        );

    \I__17100\ : InMux
    port map (
            O => \N__71277\,
            I => \N__71274\
        );

    \I__17099\ : LocalMux
    port map (
            O => \N__71274\,
            I => \N__71271\
        );

    \I__17098\ : Span4Mux_v
    port map (
            O => \N__71271\,
            I => \N__71265\
        );

    \I__17097\ : InMux
    port map (
            O => \N__71270\,
            I => \N__71260\
        );

    \I__17096\ : InMux
    port map (
            O => \N__71269\,
            I => \N__71260\
        );

    \I__17095\ : InMux
    port map (
            O => \N__71268\,
            I => \N__71257\
        );

    \I__17094\ : Span4Mux_h
    port map (
            O => \N__71265\,
            I => \N__71254\
        );

    \I__17093\ : LocalMux
    port map (
            O => \N__71260\,
            I => \c0.data_in_frame_17_6\
        );

    \I__17092\ : LocalMux
    port map (
            O => \N__71257\,
            I => \c0.data_in_frame_17_6\
        );

    \I__17091\ : Odrv4
    port map (
            O => \N__71254\,
            I => \c0.data_in_frame_17_6\
        );

    \I__17090\ : InMux
    port map (
            O => \N__71247\,
            I => \N__71243\
        );

    \I__17089\ : CascadeMux
    port map (
            O => \N__71246\,
            I => \N__71239\
        );

    \I__17088\ : LocalMux
    port map (
            O => \N__71243\,
            I => \N__71236\
        );

    \I__17087\ : InMux
    port map (
            O => \N__71242\,
            I => \N__71233\
        );

    \I__17086\ : InMux
    port map (
            O => \N__71239\,
            I => \N__71230\
        );

    \I__17085\ : Span4Mux_v
    port map (
            O => \N__71236\,
            I => \N__71225\
        );

    \I__17084\ : LocalMux
    port map (
            O => \N__71233\,
            I => \N__71225\
        );

    \I__17083\ : LocalMux
    port map (
            O => \N__71230\,
            I => \c0.data_in_frame_15_5\
        );

    \I__17082\ : Odrv4
    port map (
            O => \N__71225\,
            I => \c0.data_in_frame_15_5\
        );

    \I__17081\ : CascadeMux
    port map (
            O => \N__71220\,
            I => \N__71216\
        );

    \I__17080\ : InMux
    port map (
            O => \N__71219\,
            I => \N__71213\
        );

    \I__17079\ : InMux
    port map (
            O => \N__71216\,
            I => \N__71210\
        );

    \I__17078\ : LocalMux
    port map (
            O => \N__71213\,
            I => \N__71206\
        );

    \I__17077\ : LocalMux
    port map (
            O => \N__71210\,
            I => \N__71203\
        );

    \I__17076\ : InMux
    port map (
            O => \N__71209\,
            I => \N__71200\
        );

    \I__17075\ : Span4Mux_h
    port map (
            O => \N__71206\,
            I => \N__71197\
        );

    \I__17074\ : Span4Mux_v
    port map (
            O => \N__71203\,
            I => \N__71192\
        );

    \I__17073\ : LocalMux
    port map (
            O => \N__71200\,
            I => \N__71192\
        );

    \I__17072\ : Odrv4
    port map (
            O => \N__71197\,
            I => \c0.n31_adj_4701\
        );

    \I__17071\ : Odrv4
    port map (
            O => \N__71192\,
            I => \c0.n31_adj_4701\
        );

    \I__17070\ : CascadeMux
    port map (
            O => \N__71187\,
            I => \N__71184\
        );

    \I__17069\ : InMux
    port map (
            O => \N__71184\,
            I => \N__71181\
        );

    \I__17068\ : LocalMux
    port map (
            O => \N__71181\,
            I => \N__71178\
        );

    \I__17067\ : Span4Mux_h
    port map (
            O => \N__71178\,
            I => \N__71172\
        );

    \I__17066\ : InMux
    port map (
            O => \N__71177\,
            I => \N__71169\
        );

    \I__17065\ : CascadeMux
    port map (
            O => \N__71176\,
            I => \N__71166\
        );

    \I__17064\ : InMux
    port map (
            O => \N__71175\,
            I => \N__71163\
        );

    \I__17063\ : Span4Mux_h
    port map (
            O => \N__71172\,
            I => \N__71158\
        );

    \I__17062\ : LocalMux
    port map (
            O => \N__71169\,
            I => \N__71158\
        );

    \I__17061\ : InMux
    port map (
            O => \N__71166\,
            I => \N__71155\
        );

    \I__17060\ : LocalMux
    port map (
            O => \N__71163\,
            I => \c0.n13474\
        );

    \I__17059\ : Odrv4
    port map (
            O => \N__71158\,
            I => \c0.n13474\
        );

    \I__17058\ : LocalMux
    port map (
            O => \N__71155\,
            I => \c0.n13474\
        );

    \I__17057\ : CascadeMux
    port map (
            O => \N__71148\,
            I => \N__71145\
        );

    \I__17056\ : InMux
    port map (
            O => \N__71145\,
            I => \N__71142\
        );

    \I__17055\ : LocalMux
    port map (
            O => \N__71142\,
            I => \N__71139\
        );

    \I__17054\ : Span4Mux_h
    port map (
            O => \N__71139\,
            I => \N__71136\
        );

    \I__17053\ : Odrv4
    port map (
            O => \N__71136\,
            I => \c0.n22650\
        );

    \I__17052\ : InMux
    port map (
            O => \N__71133\,
            I => \N__71130\
        );

    \I__17051\ : LocalMux
    port map (
            O => \N__71130\,
            I => \N__71127\
        );

    \I__17050\ : Span4Mux_h
    port map (
            O => \N__71127\,
            I => \N__71123\
        );

    \I__17049\ : InMux
    port map (
            O => \N__71126\,
            I => \N__71120\
        );

    \I__17048\ : Span4Mux_h
    port map (
            O => \N__71123\,
            I => \N__71110\
        );

    \I__17047\ : LocalMux
    port map (
            O => \N__71120\,
            I => \N__71107\
        );

    \I__17046\ : InMux
    port map (
            O => \N__71119\,
            I => \N__71104\
        );

    \I__17045\ : InMux
    port map (
            O => \N__71118\,
            I => \N__71101\
        );

    \I__17044\ : InMux
    port map (
            O => \N__71117\,
            I => \N__71096\
        );

    \I__17043\ : InMux
    port map (
            O => \N__71116\,
            I => \N__71088\
        );

    \I__17042\ : InMux
    port map (
            O => \N__71115\,
            I => \N__71081\
        );

    \I__17041\ : InMux
    port map (
            O => \N__71114\,
            I => \N__71081\
        );

    \I__17040\ : InMux
    port map (
            O => \N__71113\,
            I => \N__71081\
        );

    \I__17039\ : Span4Mux_v
    port map (
            O => \N__71110\,
            I => \N__71068\
        );

    \I__17038\ : Span4Mux_h
    port map (
            O => \N__71107\,
            I => \N__71068\
        );

    \I__17037\ : LocalMux
    port map (
            O => \N__71104\,
            I => \N__71068\
        );

    \I__17036\ : LocalMux
    port map (
            O => \N__71101\,
            I => \N__71068\
        );

    \I__17035\ : InMux
    port map (
            O => \N__71100\,
            I => \N__71065\
        );

    \I__17034\ : InMux
    port map (
            O => \N__71099\,
            I => \N__71062\
        );

    \I__17033\ : LocalMux
    port map (
            O => \N__71096\,
            I => \N__71059\
        );

    \I__17032\ : InMux
    port map (
            O => \N__71095\,
            I => \N__71054\
        );

    \I__17031\ : InMux
    port map (
            O => \N__71094\,
            I => \N__71054\
        );

    \I__17030\ : InMux
    port map (
            O => \N__71093\,
            I => \N__71051\
        );

    \I__17029\ : InMux
    port map (
            O => \N__71092\,
            I => \N__71046\
        );

    \I__17028\ : InMux
    port map (
            O => \N__71091\,
            I => \N__71046\
        );

    \I__17027\ : LocalMux
    port map (
            O => \N__71088\,
            I => \N__71041\
        );

    \I__17026\ : LocalMux
    port map (
            O => \N__71081\,
            I => \N__71041\
        );

    \I__17025\ : InMux
    port map (
            O => \N__71080\,
            I => \N__71036\
        );

    \I__17024\ : InMux
    port map (
            O => \N__71079\,
            I => \N__71036\
        );

    \I__17023\ : CascadeMux
    port map (
            O => \N__71078\,
            I => \N__71033\
        );

    \I__17022\ : InMux
    port map (
            O => \N__71077\,
            I => \N__71027\
        );

    \I__17021\ : Span4Mux_v
    port map (
            O => \N__71068\,
            I => \N__71024\
        );

    \I__17020\ : LocalMux
    port map (
            O => \N__71065\,
            I => \N__71019\
        );

    \I__17019\ : LocalMux
    port map (
            O => \N__71062\,
            I => \N__71019\
        );

    \I__17018\ : Span4Mux_v
    port map (
            O => \N__71059\,
            I => \N__71016\
        );

    \I__17017\ : LocalMux
    port map (
            O => \N__71054\,
            I => \N__71005\
        );

    \I__17016\ : LocalMux
    port map (
            O => \N__71051\,
            I => \N__71005\
        );

    \I__17015\ : LocalMux
    port map (
            O => \N__71046\,
            I => \N__71005\
        );

    \I__17014\ : Span4Mux_v
    port map (
            O => \N__71041\,
            I => \N__71005\
        );

    \I__17013\ : LocalMux
    port map (
            O => \N__71036\,
            I => \N__71005\
        );

    \I__17012\ : InMux
    port map (
            O => \N__71033\,
            I => \N__71002\
        );

    \I__17011\ : InMux
    port map (
            O => \N__71032\,
            I => \N__70999\
        );

    \I__17010\ : InMux
    port map (
            O => \N__71031\,
            I => \N__70994\
        );

    \I__17009\ : InMux
    port map (
            O => \N__71030\,
            I => \N__70994\
        );

    \I__17008\ : LocalMux
    port map (
            O => \N__71027\,
            I => \N__70989\
        );

    \I__17007\ : Span4Mux_h
    port map (
            O => \N__71024\,
            I => \N__70989\
        );

    \I__17006\ : Span4Mux_v
    port map (
            O => \N__71019\,
            I => \N__70982\
        );

    \I__17005\ : Span4Mux_h
    port map (
            O => \N__71016\,
            I => \N__70982\
        );

    \I__17004\ : Span4Mux_v
    port map (
            O => \N__71005\,
            I => \N__70982\
        );

    \I__17003\ : LocalMux
    port map (
            O => \N__71002\,
            I => data_in_frame_1_7
        );

    \I__17002\ : LocalMux
    port map (
            O => \N__70999\,
            I => data_in_frame_1_7
        );

    \I__17001\ : LocalMux
    port map (
            O => \N__70994\,
            I => data_in_frame_1_7
        );

    \I__17000\ : Odrv4
    port map (
            O => \N__70989\,
            I => data_in_frame_1_7
        );

    \I__16999\ : Odrv4
    port map (
            O => \N__70982\,
            I => data_in_frame_1_7
        );

    \I__16998\ : CascadeMux
    port map (
            O => \N__70971\,
            I => \N__70968\
        );

    \I__16997\ : InMux
    port map (
            O => \N__70968\,
            I => \N__70965\
        );

    \I__16996\ : LocalMux
    port map (
            O => \N__70965\,
            I => \N__70962\
        );

    \I__16995\ : Odrv4
    port map (
            O => \N__70962\,
            I => \c0.n30_adj_4747\
        );

    \I__16994\ : InMux
    port map (
            O => \N__70959\,
            I => \N__70955\
        );

    \I__16993\ : InMux
    port map (
            O => \N__70958\,
            I => \N__70952\
        );

    \I__16992\ : LocalMux
    port map (
            O => \N__70955\,
            I => \N__70949\
        );

    \I__16991\ : LocalMux
    port map (
            O => \N__70952\,
            I => \N__70946\
        );

    \I__16990\ : Span4Mux_v
    port map (
            O => \N__70949\,
            I => \N__70943\
        );

    \I__16989\ : Span4Mux_v
    port map (
            O => \N__70946\,
            I => \N__70940\
        );

    \I__16988\ : Span4Mux_v
    port map (
            O => \N__70943\,
            I => \N__70937\
        );

    \I__16987\ : Odrv4
    port map (
            O => \N__70940\,
            I => \c0.n6_adj_4632\
        );

    \I__16986\ : Odrv4
    port map (
            O => \N__70937\,
            I => \c0.n6_adj_4632\
        );

    \I__16985\ : InMux
    port map (
            O => \N__70932\,
            I => \N__70929\
        );

    \I__16984\ : LocalMux
    port map (
            O => \N__70929\,
            I => \c0.n5_adj_4631\
        );

    \I__16983\ : InMux
    port map (
            O => \N__70926\,
            I => \N__70923\
        );

    \I__16982\ : LocalMux
    port map (
            O => \N__70923\,
            I => \N__70919\
        );

    \I__16981\ : InMux
    port map (
            O => \N__70922\,
            I => \N__70916\
        );

    \I__16980\ : Span4Mux_h
    port map (
            O => \N__70919\,
            I => \N__70910\
        );

    \I__16979\ : LocalMux
    port map (
            O => \N__70916\,
            I => \N__70910\
        );

    \I__16978\ : InMux
    port map (
            O => \N__70915\,
            I => \N__70907\
        );

    \I__16977\ : Span4Mux_v
    port map (
            O => \N__70910\,
            I => \N__70902\
        );

    \I__16976\ : LocalMux
    port map (
            O => \N__70907\,
            I => \N__70902\
        );

    \I__16975\ : Odrv4
    port map (
            O => \N__70902\,
            I => \c0.n23343\
        );

    \I__16974\ : InMux
    port map (
            O => \N__70899\,
            I => \N__70896\
        );

    \I__16973\ : LocalMux
    port map (
            O => \N__70896\,
            I => \N__70893\
        );

    \I__16972\ : Sp12to4
    port map (
            O => \N__70893\,
            I => \N__70890\
        );

    \I__16971\ : Odrv12
    port map (
            O => \N__70890\,
            I => \c0.n25_adj_4633\
        );

    \I__16970\ : InMux
    port map (
            O => \N__70887\,
            I => \N__70880\
        );

    \I__16969\ : InMux
    port map (
            O => \N__70886\,
            I => \N__70880\
        );

    \I__16968\ : InMux
    port map (
            O => \N__70885\,
            I => \N__70877\
        );

    \I__16967\ : LocalMux
    port map (
            O => \N__70880\,
            I => \N__70873\
        );

    \I__16966\ : LocalMux
    port map (
            O => \N__70877\,
            I => \N__70870\
        );

    \I__16965\ : InMux
    port map (
            O => \N__70876\,
            I => \N__70867\
        );

    \I__16964\ : Span4Mux_h
    port map (
            O => \N__70873\,
            I => \N__70864\
        );

    \I__16963\ : Span12Mux_v
    port map (
            O => \N__70870\,
            I => \N__70861\
        );

    \I__16962\ : LocalMux
    port map (
            O => \N__70867\,
            I => \c0.data_in_frame_9_3\
        );

    \I__16961\ : Odrv4
    port map (
            O => \N__70864\,
            I => \c0.data_in_frame_9_3\
        );

    \I__16960\ : Odrv12
    port map (
            O => \N__70861\,
            I => \c0.data_in_frame_9_3\
        );

    \I__16959\ : InMux
    port map (
            O => \N__70854\,
            I => \N__70851\
        );

    \I__16958\ : LocalMux
    port map (
            O => \N__70851\,
            I => \N__70844\
        );

    \I__16957\ : InMux
    port map (
            O => \N__70850\,
            I => \N__70841\
        );

    \I__16956\ : InMux
    port map (
            O => \N__70849\,
            I => \N__70838\
        );

    \I__16955\ : InMux
    port map (
            O => \N__70848\,
            I => \N__70835\
        );

    \I__16954\ : InMux
    port map (
            O => \N__70847\,
            I => \N__70832\
        );

    \I__16953\ : Span4Mux_h
    port map (
            O => \N__70844\,
            I => \N__70827\
        );

    \I__16952\ : LocalMux
    port map (
            O => \N__70841\,
            I => \N__70827\
        );

    \I__16951\ : LocalMux
    port map (
            O => \N__70838\,
            I => \c0.data_in_frame_11_2\
        );

    \I__16950\ : LocalMux
    port map (
            O => \N__70835\,
            I => \c0.data_in_frame_11_2\
        );

    \I__16949\ : LocalMux
    port map (
            O => \N__70832\,
            I => \c0.data_in_frame_11_2\
        );

    \I__16948\ : Odrv4
    port map (
            O => \N__70827\,
            I => \c0.data_in_frame_11_2\
        );

    \I__16947\ : CascadeMux
    port map (
            O => \N__70818\,
            I => \N__70815\
        );

    \I__16946\ : InMux
    port map (
            O => \N__70815\,
            I => \N__70812\
        );

    \I__16945\ : LocalMux
    port map (
            O => \N__70812\,
            I => \N__70809\
        );

    \I__16944\ : Span4Mux_v
    port map (
            O => \N__70809\,
            I => \N__70805\
        );

    \I__16943\ : CascadeMux
    port map (
            O => \N__70808\,
            I => \N__70802\
        );

    \I__16942\ : Span4Mux_h
    port map (
            O => \N__70805\,
            I => \N__70799\
        );

    \I__16941\ : InMux
    port map (
            O => \N__70802\,
            I => \N__70796\
        );

    \I__16940\ : Span4Mux_h
    port map (
            O => \N__70799\,
            I => \N__70793\
        );

    \I__16939\ : LocalMux
    port map (
            O => \N__70796\,
            I => \c0.data_in_frame_28_1\
        );

    \I__16938\ : Odrv4
    port map (
            O => \N__70793\,
            I => \c0.data_in_frame_28_1\
        );

    \I__16937\ : InMux
    port map (
            O => \N__70788\,
            I => \N__70784\
        );

    \I__16936\ : CascadeMux
    port map (
            O => \N__70787\,
            I => \N__70781\
        );

    \I__16935\ : LocalMux
    port map (
            O => \N__70784\,
            I => \N__70778\
        );

    \I__16934\ : InMux
    port map (
            O => \N__70781\,
            I => \N__70775\
        );

    \I__16933\ : Span4Mux_v
    port map (
            O => \N__70778\,
            I => \N__70771\
        );

    \I__16932\ : LocalMux
    port map (
            O => \N__70775\,
            I => \N__70768\
        );

    \I__16931\ : CascadeMux
    port map (
            O => \N__70774\,
            I => \N__70765\
        );

    \I__16930\ : Span4Mux_h
    port map (
            O => \N__70771\,
            I => \N__70760\
        );

    \I__16929\ : Span4Mux_v
    port map (
            O => \N__70768\,
            I => \N__70760\
        );

    \I__16928\ : InMux
    port map (
            O => \N__70765\,
            I => \N__70757\
        );

    \I__16927\ : Span4Mux_h
    port map (
            O => \N__70760\,
            I => \N__70754\
        );

    \I__16926\ : LocalMux
    port map (
            O => \N__70757\,
            I => \c0.data_in_frame_11_4\
        );

    \I__16925\ : Odrv4
    port map (
            O => \N__70754\,
            I => \c0.data_in_frame_11_4\
        );

    \I__16924\ : InMux
    port map (
            O => \N__70749\,
            I => \N__70746\
        );

    \I__16923\ : LocalMux
    port map (
            O => \N__70746\,
            I => \N__70743\
        );

    \I__16922\ : Span4Mux_h
    port map (
            O => \N__70743\,
            I => \N__70738\
        );

    \I__16921\ : InMux
    port map (
            O => \N__70742\,
            I => \N__70735\
        );

    \I__16920\ : CascadeMux
    port map (
            O => \N__70741\,
            I => \N__70732\
        );

    \I__16919\ : Span4Mux_v
    port map (
            O => \N__70738\,
            I => \N__70727\
        );

    \I__16918\ : LocalMux
    port map (
            O => \N__70735\,
            I => \N__70727\
        );

    \I__16917\ : InMux
    port map (
            O => \N__70732\,
            I => \N__70724\
        );

    \I__16916\ : Span4Mux_h
    port map (
            O => \N__70727\,
            I => \N__70721\
        );

    \I__16915\ : LocalMux
    port map (
            O => \N__70724\,
            I => \c0.data_in_frame_7_2\
        );

    \I__16914\ : Odrv4
    port map (
            O => \N__70721\,
            I => \c0.data_in_frame_7_2\
        );

    \I__16913\ : CascadeMux
    port map (
            O => \N__70716\,
            I => \N__70712\
        );

    \I__16912\ : InMux
    port map (
            O => \N__70715\,
            I => \N__70709\
        );

    \I__16911\ : InMux
    port map (
            O => \N__70712\,
            I => \N__70706\
        );

    \I__16910\ : LocalMux
    port map (
            O => \N__70709\,
            I => \c0.n9_adj_4220\
        );

    \I__16909\ : LocalMux
    port map (
            O => \N__70706\,
            I => \c0.n9_adj_4220\
        );

    \I__16908\ : InMux
    port map (
            O => \N__70701\,
            I => \N__70698\
        );

    \I__16907\ : LocalMux
    port map (
            O => \N__70698\,
            I => \N__70695\
        );

    \I__16906\ : Span4Mux_v
    port map (
            O => \N__70695\,
            I => \N__70691\
        );

    \I__16905\ : InMux
    port map (
            O => \N__70694\,
            I => \N__70688\
        );

    \I__16904\ : Odrv4
    port map (
            O => \N__70691\,
            I => \c0.n7_adj_4226\
        );

    \I__16903\ : LocalMux
    port map (
            O => \N__70688\,
            I => \c0.n7_adj_4226\
        );

    \I__16902\ : InMux
    port map (
            O => \N__70683\,
            I => \N__70680\
        );

    \I__16901\ : LocalMux
    port map (
            O => \N__70680\,
            I => \c0.n27_adj_4748\
        );

    \I__16900\ : CascadeMux
    port map (
            O => \N__70677\,
            I => \N__70674\
        );

    \I__16899\ : InMux
    port map (
            O => \N__70674\,
            I => \N__70669\
        );

    \I__16898\ : CascadeMux
    port map (
            O => \N__70673\,
            I => \N__70666\
        );

    \I__16897\ : InMux
    port map (
            O => \N__70672\,
            I => \N__70663\
        );

    \I__16896\ : LocalMux
    port map (
            O => \N__70669\,
            I => \N__70660\
        );

    \I__16895\ : InMux
    port map (
            O => \N__70666\,
            I => \N__70655\
        );

    \I__16894\ : LocalMux
    port map (
            O => \N__70663\,
            I => \N__70652\
        );

    \I__16893\ : Span4Mux_v
    port map (
            O => \N__70660\,
            I => \N__70649\
        );

    \I__16892\ : InMux
    port map (
            O => \N__70659\,
            I => \N__70646\
        );

    \I__16891\ : CascadeMux
    port map (
            O => \N__70658\,
            I => \N__70642\
        );

    \I__16890\ : LocalMux
    port map (
            O => \N__70655\,
            I => \N__70637\
        );

    \I__16889\ : Span4Mux_v
    port map (
            O => \N__70652\,
            I => \N__70637\
        );

    \I__16888\ : Span4Mux_h
    port map (
            O => \N__70649\,
            I => \N__70632\
        );

    \I__16887\ : LocalMux
    port map (
            O => \N__70646\,
            I => \N__70632\
        );

    \I__16886\ : InMux
    port map (
            O => \N__70645\,
            I => \N__70627\
        );

    \I__16885\ : InMux
    port map (
            O => \N__70642\,
            I => \N__70627\
        );

    \I__16884\ : Odrv4
    port map (
            O => \N__70637\,
            I => \c0.data_in_frame_11_3\
        );

    \I__16883\ : Odrv4
    port map (
            O => \N__70632\,
            I => \c0.data_in_frame_11_3\
        );

    \I__16882\ : LocalMux
    port map (
            O => \N__70627\,
            I => \c0.data_in_frame_11_3\
        );

    \I__16881\ : InMux
    port map (
            O => \N__70620\,
            I => \N__70615\
        );

    \I__16880\ : InMux
    port map (
            O => \N__70619\,
            I => \N__70612\
        );

    \I__16879\ : InMux
    port map (
            O => \N__70618\,
            I => \N__70609\
        );

    \I__16878\ : LocalMux
    port map (
            O => \N__70615\,
            I => \c0.data_in_frame_9_0\
        );

    \I__16877\ : LocalMux
    port map (
            O => \N__70612\,
            I => \c0.data_in_frame_9_0\
        );

    \I__16876\ : LocalMux
    port map (
            O => \N__70609\,
            I => \c0.data_in_frame_9_0\
        );

    \I__16875\ : InMux
    port map (
            O => \N__70602\,
            I => \N__70599\
        );

    \I__16874\ : LocalMux
    port map (
            O => \N__70599\,
            I => \N__70595\
        );

    \I__16873\ : CascadeMux
    port map (
            O => \N__70598\,
            I => \N__70592\
        );

    \I__16872\ : Span4Mux_h
    port map (
            O => \N__70595\,
            I => \N__70588\
        );

    \I__16871\ : InMux
    port map (
            O => \N__70592\,
            I => \N__70585\
        );

    \I__16870\ : InMux
    port map (
            O => \N__70591\,
            I => \N__70582\
        );

    \I__16869\ : Odrv4
    port map (
            O => \N__70588\,
            I => \c0.n4\
        );

    \I__16868\ : LocalMux
    port map (
            O => \N__70585\,
            I => \c0.n4\
        );

    \I__16867\ : LocalMux
    port map (
            O => \N__70582\,
            I => \c0.n4\
        );

    \I__16866\ : InMux
    port map (
            O => \N__70575\,
            I => \N__70572\
        );

    \I__16865\ : LocalMux
    port map (
            O => \N__70572\,
            I => \N__70568\
        );

    \I__16864\ : CascadeMux
    port map (
            O => \N__70571\,
            I => \N__70565\
        );

    \I__16863\ : Span4Mux_h
    port map (
            O => \N__70568\,
            I => \N__70562\
        );

    \I__16862\ : InMux
    port map (
            O => \N__70565\,
            I => \N__70559\
        );

    \I__16861\ : Span4Mux_v
    port map (
            O => \N__70562\,
            I => \N__70556\
        );

    \I__16860\ : LocalMux
    port map (
            O => \N__70559\,
            I => \c0.data_in_frame_28_3\
        );

    \I__16859\ : Odrv4
    port map (
            O => \N__70556\,
            I => \c0.data_in_frame_28_3\
        );

    \I__16858\ : InMux
    port map (
            O => \N__70551\,
            I => \N__70545\
        );

    \I__16857\ : CascadeMux
    port map (
            O => \N__70550\,
            I => \N__70542\
        );

    \I__16856\ : InMux
    port map (
            O => \N__70549\,
            I => \N__70537\
        );

    \I__16855\ : InMux
    port map (
            O => \N__70548\,
            I => \N__70537\
        );

    \I__16854\ : LocalMux
    port map (
            O => \N__70545\,
            I => \N__70534\
        );

    \I__16853\ : InMux
    port map (
            O => \N__70542\,
            I => \N__70531\
        );

    \I__16852\ : LocalMux
    port map (
            O => \N__70537\,
            I => \N__70528\
        );

    \I__16851\ : Span4Mux_h
    port map (
            O => \N__70534\,
            I => \N__70524\
        );

    \I__16850\ : LocalMux
    port map (
            O => \N__70531\,
            I => \N__70519\
        );

    \I__16849\ : Span4Mux_v
    port map (
            O => \N__70528\,
            I => \N__70519\
        );

    \I__16848\ : InMux
    port map (
            O => \N__70527\,
            I => \N__70516\
        );

    \I__16847\ : Span4Mux_h
    port map (
            O => \N__70524\,
            I => \N__70513\
        );

    \I__16846\ : Odrv4
    port map (
            O => \N__70519\,
            I => \c0.data_in_frame_12_3\
        );

    \I__16845\ : LocalMux
    port map (
            O => \N__70516\,
            I => \c0.data_in_frame_12_3\
        );

    \I__16844\ : Odrv4
    port map (
            O => \N__70513\,
            I => \c0.data_in_frame_12_3\
        );

    \I__16843\ : CascadeMux
    port map (
            O => \N__70506\,
            I => \N__70502\
        );

    \I__16842\ : InMux
    port map (
            O => \N__70505\,
            I => \N__70499\
        );

    \I__16841\ : InMux
    port map (
            O => \N__70502\,
            I => \N__70495\
        );

    \I__16840\ : LocalMux
    port map (
            O => \N__70499\,
            I => \N__70492\
        );

    \I__16839\ : InMux
    port map (
            O => \N__70498\,
            I => \N__70489\
        );

    \I__16838\ : LocalMux
    port map (
            O => \N__70495\,
            I => \c0.data_in_frame_15_6\
        );

    \I__16837\ : Odrv4
    port map (
            O => \N__70492\,
            I => \c0.data_in_frame_15_6\
        );

    \I__16836\ : LocalMux
    port map (
            O => \N__70489\,
            I => \c0.data_in_frame_15_6\
        );

    \I__16835\ : CascadeMux
    port map (
            O => \N__70482\,
            I => \N__70479\
        );

    \I__16834\ : InMux
    port map (
            O => \N__70479\,
            I => \N__70476\
        );

    \I__16833\ : LocalMux
    port map (
            O => \N__70476\,
            I => \N__70473\
        );

    \I__16832\ : Span4Mux_h
    port map (
            O => \N__70473\,
            I => \N__70470\
        );

    \I__16831\ : Span4Mux_h
    port map (
            O => \N__70470\,
            I => \N__70466\
        );

    \I__16830\ : InMux
    port map (
            O => \N__70469\,
            I => \N__70463\
        );

    \I__16829\ : Odrv4
    port map (
            O => \N__70466\,
            I => \c0.n22379\
        );

    \I__16828\ : LocalMux
    port map (
            O => \N__70463\,
            I => \c0.n22379\
        );

    \I__16827\ : CascadeMux
    port map (
            O => \N__70458\,
            I => \N__70455\
        );

    \I__16826\ : InMux
    port map (
            O => \N__70455\,
            I => \N__70452\
        );

    \I__16825\ : LocalMux
    port map (
            O => \N__70452\,
            I => \c0.n6_adj_4559\
        );

    \I__16824\ : CascadeMux
    port map (
            O => \N__70449\,
            I => \N__70446\
        );

    \I__16823\ : InMux
    port map (
            O => \N__70446\,
            I => \N__70440\
        );

    \I__16822\ : InMux
    port map (
            O => \N__70445\,
            I => \N__70432\
        );

    \I__16821\ : InMux
    port map (
            O => \N__70444\,
            I => \N__70432\
        );

    \I__16820\ : InMux
    port map (
            O => \N__70443\,
            I => \N__70432\
        );

    \I__16819\ : LocalMux
    port map (
            O => \N__70440\,
            I => \N__70429\
        );

    \I__16818\ : InMux
    port map (
            O => \N__70439\,
            I => \N__70426\
        );

    \I__16817\ : LocalMux
    port map (
            O => \N__70432\,
            I => \N__70422\
        );

    \I__16816\ : Span4Mux_v
    port map (
            O => \N__70429\,
            I => \N__70417\
        );

    \I__16815\ : LocalMux
    port map (
            O => \N__70426\,
            I => \N__70417\
        );

    \I__16814\ : InMux
    port map (
            O => \N__70425\,
            I => \N__70414\
        );

    \I__16813\ : Span4Mux_h
    port map (
            O => \N__70422\,
            I => \N__70411\
        );

    \I__16812\ : Span4Mux_h
    port map (
            O => \N__70417\,
            I => \N__70408\
        );

    \I__16811\ : LocalMux
    port map (
            O => \N__70414\,
            I => \c0.data_in_frame_9_5\
        );

    \I__16810\ : Odrv4
    port map (
            O => \N__70411\,
            I => \c0.data_in_frame_9_5\
        );

    \I__16809\ : Odrv4
    port map (
            O => \N__70408\,
            I => \c0.data_in_frame_9_5\
        );

    \I__16808\ : InMux
    port map (
            O => \N__70401\,
            I => \N__70397\
        );

    \I__16807\ : InMux
    port map (
            O => \N__70400\,
            I => \N__70394\
        );

    \I__16806\ : LocalMux
    port map (
            O => \N__70397\,
            I => \N__70391\
        );

    \I__16805\ : LocalMux
    port map (
            O => \N__70394\,
            I => \N__70388\
        );

    \I__16804\ : Span4Mux_v
    port map (
            O => \N__70391\,
            I => \N__70384\
        );

    \I__16803\ : Span12Mux_h
    port map (
            O => \N__70388\,
            I => \N__70381\
        );

    \I__16802\ : InMux
    port map (
            O => \N__70387\,
            I => \N__70378\
        );

    \I__16801\ : Sp12to4
    port map (
            O => \N__70384\,
            I => \N__70373\
        );

    \I__16800\ : Span12Mux_v
    port map (
            O => \N__70381\,
            I => \N__70373\
        );

    \I__16799\ : LocalMux
    port map (
            O => \N__70378\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__16798\ : Odrv12
    port map (
            O => \N__70373\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__16797\ : SRMux
    port map (
            O => \N__70368\,
            I => \N__70365\
        );

    \I__16796\ : LocalMux
    port map (
            O => \N__70365\,
            I => \N__70362\
        );

    \I__16795\ : Span4Mux_v
    port map (
            O => \N__70362\,
            I => \N__70359\
        );

    \I__16794\ : Span4Mux_h
    port map (
            O => \N__70359\,
            I => \N__70356\
        );

    \I__16793\ : Odrv4
    port map (
            O => \N__70356\,
            I => \c0.n3_adj_4410\
        );

    \I__16792\ : InMux
    port map (
            O => \N__70353\,
            I => \N__70349\
        );

    \I__16791\ : InMux
    port map (
            O => \N__70352\,
            I => \N__70344\
        );

    \I__16790\ : LocalMux
    port map (
            O => \N__70349\,
            I => \N__70341\
        );

    \I__16789\ : InMux
    port map (
            O => \N__70348\,
            I => \N__70338\
        );

    \I__16788\ : CascadeMux
    port map (
            O => \N__70347\,
            I => \N__70335\
        );

    \I__16787\ : LocalMux
    port map (
            O => \N__70344\,
            I => \N__70332\
        );

    \I__16786\ : Span4Mux_h
    port map (
            O => \N__70341\,
            I => \N__70329\
        );

    \I__16785\ : LocalMux
    port map (
            O => \N__70338\,
            I => \N__70325\
        );

    \I__16784\ : InMux
    port map (
            O => \N__70335\,
            I => \N__70322\
        );

    \I__16783\ : Span4Mux_h
    port map (
            O => \N__70332\,
            I => \N__70319\
        );

    \I__16782\ : Span4Mux_h
    port map (
            O => \N__70329\,
            I => \N__70316\
        );

    \I__16781\ : InMux
    port map (
            O => \N__70328\,
            I => \N__70313\
        );

    \I__16780\ : Span4Mux_h
    port map (
            O => \N__70325\,
            I => \N__70310\
        );

    \I__16779\ : LocalMux
    port map (
            O => \N__70322\,
            I => \c0.data_in_frame_7_4\
        );

    \I__16778\ : Odrv4
    port map (
            O => \N__70319\,
            I => \c0.data_in_frame_7_4\
        );

    \I__16777\ : Odrv4
    port map (
            O => \N__70316\,
            I => \c0.data_in_frame_7_4\
        );

    \I__16776\ : LocalMux
    port map (
            O => \N__70313\,
            I => \c0.data_in_frame_7_4\
        );

    \I__16775\ : Odrv4
    port map (
            O => \N__70310\,
            I => \c0.data_in_frame_7_4\
        );

    \I__16774\ : InMux
    port map (
            O => \N__70299\,
            I => \N__70294\
        );

    \I__16773\ : InMux
    port map (
            O => \N__70298\,
            I => \N__70291\
        );

    \I__16772\ : InMux
    port map (
            O => \N__70297\,
            I => \N__70288\
        );

    \I__16771\ : LocalMux
    port map (
            O => \N__70294\,
            I => \N__70285\
        );

    \I__16770\ : LocalMux
    port map (
            O => \N__70291\,
            I => \N__70281\
        );

    \I__16769\ : LocalMux
    port map (
            O => \N__70288\,
            I => \N__70278\
        );

    \I__16768\ : Span4Mux_v
    port map (
            O => \N__70285\,
            I => \N__70274\
        );

    \I__16767\ : InMux
    port map (
            O => \N__70284\,
            I => \N__70271\
        );

    \I__16766\ : Span4Mux_v
    port map (
            O => \N__70281\,
            I => \N__70268\
        );

    \I__16765\ : Span4Mux_v
    port map (
            O => \N__70278\,
            I => \N__70265\
        );

    \I__16764\ : CascadeMux
    port map (
            O => \N__70277\,
            I => \N__70261\
        );

    \I__16763\ : Span4Mux_h
    port map (
            O => \N__70274\,
            I => \N__70258\
        );

    \I__16762\ : LocalMux
    port map (
            O => \N__70271\,
            I => \N__70253\
        );

    \I__16761\ : Span4Mux_h
    port map (
            O => \N__70268\,
            I => \N__70253\
        );

    \I__16760\ : Span4Mux_h
    port map (
            O => \N__70265\,
            I => \N__70250\
        );

    \I__16759\ : InMux
    port map (
            O => \N__70264\,
            I => \N__70247\
        );

    \I__16758\ : InMux
    port map (
            O => \N__70261\,
            I => \N__70244\
        );

    \I__16757\ : Odrv4
    port map (
            O => \N__70258\,
            I => data_in_frame_5_1
        );

    \I__16756\ : Odrv4
    port map (
            O => \N__70253\,
            I => data_in_frame_5_1
        );

    \I__16755\ : Odrv4
    port map (
            O => \N__70250\,
            I => data_in_frame_5_1
        );

    \I__16754\ : LocalMux
    port map (
            O => \N__70247\,
            I => data_in_frame_5_1
        );

    \I__16753\ : LocalMux
    port map (
            O => \N__70244\,
            I => data_in_frame_5_1
        );

    \I__16752\ : InMux
    port map (
            O => \N__70233\,
            I => \N__70230\
        );

    \I__16751\ : LocalMux
    port map (
            O => \N__70230\,
            I => \N__70226\
        );

    \I__16750\ : InMux
    port map (
            O => \N__70229\,
            I => \N__70222\
        );

    \I__16749\ : Span4Mux_h
    port map (
            O => \N__70226\,
            I => \N__70219\
        );

    \I__16748\ : InMux
    port map (
            O => \N__70225\,
            I => \N__70216\
        );

    \I__16747\ : LocalMux
    port map (
            O => \N__70222\,
            I => \N__70212\
        );

    \I__16746\ : Span4Mux_h
    port map (
            O => \N__70219\,
            I => \N__70209\
        );

    \I__16745\ : LocalMux
    port map (
            O => \N__70216\,
            I => \N__70206\
        );

    \I__16744\ : InMux
    port map (
            O => \N__70215\,
            I => \N__70203\
        );

    \I__16743\ : Odrv12
    port map (
            O => \N__70212\,
            I => \c0.n40_adj_4288\
        );

    \I__16742\ : Odrv4
    port map (
            O => \N__70209\,
            I => \c0.n40_adj_4288\
        );

    \I__16741\ : Odrv4
    port map (
            O => \N__70206\,
            I => \c0.n40_adj_4288\
        );

    \I__16740\ : LocalMux
    port map (
            O => \N__70203\,
            I => \c0.n40_adj_4288\
        );

    \I__16739\ : InMux
    port map (
            O => \N__70194\,
            I => \N__70188\
        );

    \I__16738\ : InMux
    port map (
            O => \N__70193\,
            I => \N__70188\
        );

    \I__16737\ : LocalMux
    port map (
            O => \N__70188\,
            I => \N__70183\
        );

    \I__16736\ : InMux
    port map (
            O => \N__70187\,
            I => \N__70180\
        );

    \I__16735\ : CascadeMux
    port map (
            O => \N__70186\,
            I => \N__70175\
        );

    \I__16734\ : Span4Mux_v
    port map (
            O => \N__70183\,
            I => \N__70159\
        );

    \I__16733\ : LocalMux
    port map (
            O => \N__70180\,
            I => \N__70159\
        );

    \I__16732\ : InMux
    port map (
            O => \N__70179\,
            I => \N__70156\
        );

    \I__16731\ : InMux
    port map (
            O => \N__70178\,
            I => \N__70131\
        );

    \I__16730\ : InMux
    port map (
            O => \N__70175\,
            I => \N__70131\
        );

    \I__16729\ : InMux
    port map (
            O => \N__70174\,
            I => \N__70131\
        );

    \I__16728\ : InMux
    port map (
            O => \N__70173\,
            I => \N__70128\
        );

    \I__16727\ : InMux
    port map (
            O => \N__70172\,
            I => \N__70121\
        );

    \I__16726\ : InMux
    port map (
            O => \N__70171\,
            I => \N__70121\
        );

    \I__16725\ : InMux
    port map (
            O => \N__70170\,
            I => \N__70121\
        );

    \I__16724\ : InMux
    port map (
            O => \N__70169\,
            I => \N__70116\
        );

    \I__16723\ : InMux
    port map (
            O => \N__70168\,
            I => \N__70116\
        );

    \I__16722\ : InMux
    port map (
            O => \N__70167\,
            I => \N__70107\
        );

    \I__16721\ : InMux
    port map (
            O => \N__70166\,
            I => \N__70107\
        );

    \I__16720\ : InMux
    port map (
            O => \N__70165\,
            I => \N__70107\
        );

    \I__16719\ : InMux
    port map (
            O => \N__70164\,
            I => \N__70107\
        );

    \I__16718\ : Span4Mux_h
    port map (
            O => \N__70159\,
            I => \N__70102\
        );

    \I__16717\ : LocalMux
    port map (
            O => \N__70156\,
            I => \N__70102\
        );

    \I__16716\ : InMux
    port map (
            O => \N__70155\,
            I => \N__70097\
        );

    \I__16715\ : InMux
    port map (
            O => \N__70154\,
            I => \N__70097\
        );

    \I__16714\ : InMux
    port map (
            O => \N__70153\,
            I => \N__70094\
        );

    \I__16713\ : InMux
    port map (
            O => \N__70152\,
            I => \N__70091\
        );

    \I__16712\ : InMux
    port map (
            O => \N__70151\,
            I => \N__70088\
        );

    \I__16711\ : CascadeMux
    port map (
            O => \N__70150\,
            I => \N__70084\
        );

    \I__16710\ : InMux
    port map (
            O => \N__70149\,
            I => \N__70075\
        );

    \I__16709\ : InMux
    port map (
            O => \N__70148\,
            I => \N__70070\
        );

    \I__16708\ : InMux
    port map (
            O => \N__70147\,
            I => \N__70070\
        );

    \I__16707\ : InMux
    port map (
            O => \N__70146\,
            I => \N__70063\
        );

    \I__16706\ : InMux
    port map (
            O => \N__70145\,
            I => \N__70063\
        );

    \I__16705\ : InMux
    port map (
            O => \N__70144\,
            I => \N__70063\
        );

    \I__16704\ : InMux
    port map (
            O => \N__70143\,
            I => \N__70058\
        );

    \I__16703\ : InMux
    port map (
            O => \N__70142\,
            I => \N__70058\
        );

    \I__16702\ : InMux
    port map (
            O => \N__70141\,
            I => \N__70055\
        );

    \I__16701\ : InMux
    port map (
            O => \N__70140\,
            I => \N__70048\
        );

    \I__16700\ : InMux
    port map (
            O => \N__70139\,
            I => \N__70048\
        );

    \I__16699\ : InMux
    port map (
            O => \N__70138\,
            I => \N__70048\
        );

    \I__16698\ : LocalMux
    port map (
            O => \N__70131\,
            I => \N__70045\
        );

    \I__16697\ : LocalMux
    port map (
            O => \N__70128\,
            I => \N__70038\
        );

    \I__16696\ : LocalMux
    port map (
            O => \N__70121\,
            I => \N__70038\
        );

    \I__16695\ : LocalMux
    port map (
            O => \N__70116\,
            I => \N__70038\
        );

    \I__16694\ : LocalMux
    port map (
            O => \N__70107\,
            I => \N__70031\
        );

    \I__16693\ : Span4Mux_h
    port map (
            O => \N__70102\,
            I => \N__70031\
        );

    \I__16692\ : LocalMux
    port map (
            O => \N__70097\,
            I => \N__70031\
        );

    \I__16691\ : LocalMux
    port map (
            O => \N__70094\,
            I => \N__70024\
        );

    \I__16690\ : LocalMux
    port map (
            O => \N__70091\,
            I => \N__70024\
        );

    \I__16689\ : LocalMux
    port map (
            O => \N__70088\,
            I => \N__70024\
        );

    \I__16688\ : CascadeMux
    port map (
            O => \N__70087\,
            I => \N__70019\
        );

    \I__16687\ : InMux
    port map (
            O => \N__70084\,
            I => \N__70005\
        );

    \I__16686\ : InMux
    port map (
            O => \N__70083\,
            I => \N__70005\
        );

    \I__16685\ : InMux
    port map (
            O => \N__70082\,
            I => \N__70005\
        );

    \I__16684\ : InMux
    port map (
            O => \N__70081\,
            I => \N__70005\
        );

    \I__16683\ : InMux
    port map (
            O => \N__70080\,
            I => \N__69998\
        );

    \I__16682\ : InMux
    port map (
            O => \N__70079\,
            I => \N__69998\
        );

    \I__16681\ : InMux
    port map (
            O => \N__70078\,
            I => \N__69998\
        );

    \I__16680\ : LocalMux
    port map (
            O => \N__70075\,
            I => \N__69993\
        );

    \I__16679\ : LocalMux
    port map (
            O => \N__70070\,
            I => \N__69993\
        );

    \I__16678\ : LocalMux
    port map (
            O => \N__70063\,
            I => \N__69988\
        );

    \I__16677\ : LocalMux
    port map (
            O => \N__70058\,
            I => \N__69988\
        );

    \I__16676\ : LocalMux
    port map (
            O => \N__70055\,
            I => \N__69979\
        );

    \I__16675\ : LocalMux
    port map (
            O => \N__70048\,
            I => \N__69979\
        );

    \I__16674\ : Span4Mux_h
    port map (
            O => \N__70045\,
            I => \N__69979\
        );

    \I__16673\ : Span4Mux_v
    port map (
            O => \N__70038\,
            I => \N__69979\
        );

    \I__16672\ : Span4Mux_v
    port map (
            O => \N__70031\,
            I => \N__69974\
        );

    \I__16671\ : Span4Mux_v
    port map (
            O => \N__70024\,
            I => \N__69974\
        );

    \I__16670\ : InMux
    port map (
            O => \N__70023\,
            I => \N__69969\
        );

    \I__16669\ : InMux
    port map (
            O => \N__70022\,
            I => \N__69969\
        );

    \I__16668\ : InMux
    port map (
            O => \N__70019\,
            I => \N__69966\
        );

    \I__16667\ : InMux
    port map (
            O => \N__70018\,
            I => \N__69963\
        );

    \I__16666\ : InMux
    port map (
            O => \N__70017\,
            I => \N__69954\
        );

    \I__16665\ : InMux
    port map (
            O => \N__70016\,
            I => \N__69954\
        );

    \I__16664\ : InMux
    port map (
            O => \N__70015\,
            I => \N__69954\
        );

    \I__16663\ : InMux
    port map (
            O => \N__70014\,
            I => \N__69954\
        );

    \I__16662\ : LocalMux
    port map (
            O => \N__70005\,
            I => \N__69951\
        );

    \I__16661\ : LocalMux
    port map (
            O => \N__69998\,
            I => \N__69946\
        );

    \I__16660\ : Span4Mux_v
    port map (
            O => \N__69993\,
            I => \N__69946\
        );

    \I__16659\ : Span4Mux_h
    port map (
            O => \N__69988\,
            I => \N__69941\
        );

    \I__16658\ : Span4Mux_h
    port map (
            O => \N__69979\,
            I => \N__69941\
        );

    \I__16657\ : Sp12to4
    port map (
            O => \N__69974\,
            I => \N__69938\
        );

    \I__16656\ : LocalMux
    port map (
            O => \N__69969\,
            I => \N__69935\
        );

    \I__16655\ : LocalMux
    port map (
            O => \N__69966\,
            I => \N__69928\
        );

    \I__16654\ : LocalMux
    port map (
            O => \N__69963\,
            I => \N__69928\
        );

    \I__16653\ : LocalMux
    port map (
            O => \N__69954\,
            I => \N__69928\
        );

    \I__16652\ : Span4Mux_v
    port map (
            O => \N__69951\,
            I => \N__69925\
        );

    \I__16651\ : Span4Mux_h
    port map (
            O => \N__69946\,
            I => \N__69920\
        );

    \I__16650\ : Span4Mux_v
    port map (
            O => \N__69941\,
            I => \N__69920\
        );

    \I__16649\ : Span12Mux_h
    port map (
            O => \N__69938\,
            I => \N__69917\
        );

    \I__16648\ : Span4Mux_v
    port map (
            O => \N__69935\,
            I => \N__69912\
        );

    \I__16647\ : Span4Mux_h
    port map (
            O => \N__69928\,
            I => \N__69912\
        );

    \I__16646\ : Odrv4
    port map (
            O => \N__69925\,
            I => \c0.n22120\
        );

    \I__16645\ : Odrv4
    port map (
            O => \N__69920\,
            I => \c0.n22120\
        );

    \I__16644\ : Odrv12
    port map (
            O => \N__69917\,
            I => \c0.n22120\
        );

    \I__16643\ : Odrv4
    port map (
            O => \N__69912\,
            I => \c0.n22120\
        );

    \I__16642\ : InMux
    port map (
            O => \N__69903\,
            I => \N__69899\
        );

    \I__16641\ : CascadeMux
    port map (
            O => \N__69902\,
            I => \N__69895\
        );

    \I__16640\ : LocalMux
    port map (
            O => \N__69899\,
            I => \N__69891\
        );

    \I__16639\ : InMux
    port map (
            O => \N__69898\,
            I => \N__69888\
        );

    \I__16638\ : InMux
    port map (
            O => \N__69895\,
            I => \N__69885\
        );

    \I__16637\ : InMux
    port map (
            O => \N__69894\,
            I => \N__69881\
        );

    \I__16636\ : Span4Mux_h
    port map (
            O => \N__69891\,
            I => \N__69878\
        );

    \I__16635\ : LocalMux
    port map (
            O => \N__69888\,
            I => \N__69873\
        );

    \I__16634\ : LocalMux
    port map (
            O => \N__69885\,
            I => \N__69873\
        );

    \I__16633\ : CascadeMux
    port map (
            O => \N__69884\,
            I => \N__69870\
        );

    \I__16632\ : LocalMux
    port map (
            O => \N__69881\,
            I => \N__69867\
        );

    \I__16631\ : Span4Mux_v
    port map (
            O => \N__69878\,
            I => \N__69862\
        );

    \I__16630\ : Span4Mux_v
    port map (
            O => \N__69873\,
            I => \N__69862\
        );

    \I__16629\ : InMux
    port map (
            O => \N__69870\,
            I => \N__69857\
        );

    \I__16628\ : Span4Mux_v
    port map (
            O => \N__69867\,
            I => \N__69852\
        );

    \I__16627\ : Span4Mux_h
    port map (
            O => \N__69862\,
            I => \N__69852\
        );

    \I__16626\ : InMux
    port map (
            O => \N__69861\,
            I => \N__69847\
        );

    \I__16625\ : InMux
    port map (
            O => \N__69860\,
            I => \N__69847\
        );

    \I__16624\ : LocalMux
    port map (
            O => \N__69857\,
            I => \N__69844\
        );

    \I__16623\ : Odrv4
    port map (
            O => \N__69852\,
            I => \c0.data_in_frame_7_3\
        );

    \I__16622\ : LocalMux
    port map (
            O => \N__69847\,
            I => \c0.data_in_frame_7_3\
        );

    \I__16621\ : Odrv4
    port map (
            O => \N__69844\,
            I => \c0.data_in_frame_7_3\
        );

    \I__16620\ : InMux
    port map (
            O => \N__69837\,
            I => \N__69834\
        );

    \I__16619\ : LocalMux
    port map (
            O => \N__69834\,
            I => \N__69829\
        );

    \I__16618\ : CascadeMux
    port map (
            O => \N__69833\,
            I => \N__69826\
        );

    \I__16617\ : CascadeMux
    port map (
            O => \N__69832\,
            I => \N__69822\
        );

    \I__16616\ : Span4Mux_h
    port map (
            O => \N__69829\,
            I => \N__69819\
        );

    \I__16615\ : InMux
    port map (
            O => \N__69826\,
            I => \N__69814\
        );

    \I__16614\ : InMux
    port map (
            O => \N__69825\,
            I => \N__69814\
        );

    \I__16613\ : InMux
    port map (
            O => \N__69822\,
            I => \N__69811\
        );

    \I__16612\ : Odrv4
    port map (
            O => \N__69819\,
            I => \c0.data_in_frame_12_0\
        );

    \I__16611\ : LocalMux
    port map (
            O => \N__69814\,
            I => \c0.data_in_frame_12_0\
        );

    \I__16610\ : LocalMux
    port map (
            O => \N__69811\,
            I => \c0.data_in_frame_12_0\
        );

    \I__16609\ : InMux
    port map (
            O => \N__69804\,
            I => \N__69801\
        );

    \I__16608\ : LocalMux
    port map (
            O => \N__69801\,
            I => \N__69797\
        );

    \I__16607\ : InMux
    port map (
            O => \N__69800\,
            I => \N__69794\
        );

    \I__16606\ : Span4Mux_v
    port map (
            O => \N__69797\,
            I => \N__69789\
        );

    \I__16605\ : LocalMux
    port map (
            O => \N__69794\,
            I => \N__69785\
        );

    \I__16604\ : InMux
    port map (
            O => \N__69793\,
            I => \N__69780\
        );

    \I__16603\ : InMux
    port map (
            O => \N__69792\,
            I => \N__69780\
        );

    \I__16602\ : Span4Mux_h
    port map (
            O => \N__69789\,
            I => \N__69777\
        );

    \I__16601\ : InMux
    port map (
            O => \N__69788\,
            I => \N__69774\
        );

    \I__16600\ : Odrv12
    port map (
            O => \N__69785\,
            I => \c0.data_in_frame_12_1\
        );

    \I__16599\ : LocalMux
    port map (
            O => \N__69780\,
            I => \c0.data_in_frame_12_1\
        );

    \I__16598\ : Odrv4
    port map (
            O => \N__69777\,
            I => \c0.data_in_frame_12_1\
        );

    \I__16597\ : LocalMux
    port map (
            O => \N__69774\,
            I => \c0.data_in_frame_12_1\
        );

    \I__16596\ : InMux
    port map (
            O => \N__69765\,
            I => \N__69762\
        );

    \I__16595\ : LocalMux
    port map (
            O => \N__69762\,
            I => \N__69755\
        );

    \I__16594\ : InMux
    port map (
            O => \N__69761\,
            I => \N__69752\
        );

    \I__16593\ : InMux
    port map (
            O => \N__69760\,
            I => \N__69747\
        );

    \I__16592\ : InMux
    port map (
            O => \N__69759\,
            I => \N__69747\
        );

    \I__16591\ : InMux
    port map (
            O => \N__69758\,
            I => \N__69744\
        );

    \I__16590\ : Span4Mux_h
    port map (
            O => \N__69755\,
            I => \N__69741\
        );

    \I__16589\ : LocalMux
    port map (
            O => \N__69752\,
            I => \N__69738\
        );

    \I__16588\ : LocalMux
    port map (
            O => \N__69747\,
            I => \N__69735\
        );

    \I__16587\ : LocalMux
    port map (
            O => \N__69744\,
            I => \N__69732\
        );

    \I__16586\ : Span4Mux_h
    port map (
            O => \N__69741\,
            I => \N__69729\
        );

    \I__16585\ : Span4Mux_v
    port map (
            O => \N__69738\,
            I => \N__69725\
        );

    \I__16584\ : Span4Mux_v
    port map (
            O => \N__69735\,
            I => \N__69720\
        );

    \I__16583\ : Span4Mux_h
    port map (
            O => \N__69732\,
            I => \N__69720\
        );

    \I__16582\ : Span4Mux_v
    port map (
            O => \N__69729\,
            I => \N__69717\
        );

    \I__16581\ : InMux
    port map (
            O => \N__69728\,
            I => \N__69714\
        );

    \I__16580\ : Span4Mux_h
    port map (
            O => \N__69725\,
            I => \N__69709\
        );

    \I__16579\ : Span4Mux_v
    port map (
            O => \N__69720\,
            I => \N__69709\
        );

    \I__16578\ : Odrv4
    port map (
            O => \N__69717\,
            I => \c0.n39\
        );

    \I__16577\ : LocalMux
    port map (
            O => \N__69714\,
            I => \c0.n39\
        );

    \I__16576\ : Odrv4
    port map (
            O => \N__69709\,
            I => \c0.n39\
        );

    \I__16575\ : InMux
    port map (
            O => \N__69702\,
            I => \N__69697\
        );

    \I__16574\ : InMux
    port map (
            O => \N__69701\,
            I => \N__69694\
        );

    \I__16573\ : InMux
    port map (
            O => \N__69700\,
            I => \N__69690\
        );

    \I__16572\ : LocalMux
    port map (
            O => \N__69697\,
            I => \N__69687\
        );

    \I__16571\ : LocalMux
    port map (
            O => \N__69694\,
            I => \N__69684\
        );

    \I__16570\ : InMux
    port map (
            O => \N__69693\,
            I => \N__69681\
        );

    \I__16569\ : LocalMux
    port map (
            O => \N__69690\,
            I => \N__69672\
        );

    \I__16568\ : Span4Mux_h
    port map (
            O => \N__69687\,
            I => \N__69672\
        );

    \I__16567\ : Span4Mux_v
    port map (
            O => \N__69684\,
            I => \N__69672\
        );

    \I__16566\ : LocalMux
    port map (
            O => \N__69681\,
            I => \N__69672\
        );

    \I__16565\ : Odrv4
    port map (
            O => \N__69672\,
            I => \c0.n61\
        );

    \I__16564\ : CascadeMux
    port map (
            O => \N__69669\,
            I => \N__69666\
        );

    \I__16563\ : InMux
    port map (
            O => \N__69666\,
            I => \N__69663\
        );

    \I__16562\ : LocalMux
    port map (
            O => \N__69663\,
            I => \N__69660\
        );

    \I__16561\ : Span4Mux_v
    port map (
            O => \N__69660\,
            I => \N__69657\
        );

    \I__16560\ : Span4Mux_h
    port map (
            O => \N__69657\,
            I => \N__69654\
        );

    \I__16559\ : Span4Mux_h
    port map (
            O => \N__69654\,
            I => \N__69651\
        );

    \I__16558\ : Odrv4
    port map (
            O => \N__69651\,
            I => \c0.n13253\
        );

    \I__16557\ : CascadeMux
    port map (
            O => \N__69648\,
            I => \c0.n13253_cascade_\
        );

    \I__16556\ : CascadeMux
    port map (
            O => \N__69645\,
            I => \N__69641\
        );

    \I__16555\ : InMux
    port map (
            O => \N__69644\,
            I => \N__69637\
        );

    \I__16554\ : InMux
    port map (
            O => \N__69641\,
            I => \N__69634\
        );

    \I__16553\ : CascadeMux
    port map (
            O => \N__69640\,
            I => \N__69631\
        );

    \I__16552\ : LocalMux
    port map (
            O => \N__69637\,
            I => \N__69627\
        );

    \I__16551\ : LocalMux
    port map (
            O => \N__69634\,
            I => \N__69624\
        );

    \I__16550\ : InMux
    port map (
            O => \N__69631\,
            I => \N__69619\
        );

    \I__16549\ : InMux
    port map (
            O => \N__69630\,
            I => \N__69619\
        );

    \I__16548\ : Span4Mux_h
    port map (
            O => \N__69627\,
            I => \N__69616\
        );

    \I__16547\ : Odrv4
    port map (
            O => \N__69624\,
            I => \c0.n22518\
        );

    \I__16546\ : LocalMux
    port map (
            O => \N__69619\,
            I => \c0.n22518\
        );

    \I__16545\ : Odrv4
    port map (
            O => \N__69616\,
            I => \c0.n22518\
        );

    \I__16544\ : InMux
    port map (
            O => \N__69609\,
            I => \N__69605\
        );

    \I__16543\ : InMux
    port map (
            O => \N__69608\,
            I => \N__69602\
        );

    \I__16542\ : LocalMux
    port map (
            O => \N__69605\,
            I => \N__69599\
        );

    \I__16541\ : LocalMux
    port map (
            O => \N__69602\,
            I => \N__69596\
        );

    \I__16540\ : Span4Mux_v
    port map (
            O => \N__69599\,
            I => \N__69593\
        );

    \I__16539\ : Sp12to4
    port map (
            O => \N__69596\,
            I => \N__69590\
        );

    \I__16538\ : Odrv4
    port map (
            O => \N__69593\,
            I => \c0.n22828\
        );

    \I__16537\ : Odrv12
    port map (
            O => \N__69590\,
            I => \c0.n22828\
        );

    \I__16536\ : InMux
    port map (
            O => \N__69585\,
            I => \N__69577\
        );

    \I__16535\ : InMux
    port map (
            O => \N__69584\,
            I => \N__69574\
        );

    \I__16534\ : InMux
    port map (
            O => \N__69583\,
            I => \N__69567\
        );

    \I__16533\ : InMux
    port map (
            O => \N__69582\,
            I => \N__69567\
        );

    \I__16532\ : InMux
    port map (
            O => \N__69581\,
            I => \N__69567\
        );

    \I__16531\ : InMux
    port map (
            O => \N__69580\,
            I => \N__69564\
        );

    \I__16530\ : LocalMux
    port map (
            O => \N__69577\,
            I => \N__69561\
        );

    \I__16529\ : LocalMux
    port map (
            O => \N__69574\,
            I => \N__69558\
        );

    \I__16528\ : LocalMux
    port map (
            O => \N__69567\,
            I => \N__69554\
        );

    \I__16527\ : LocalMux
    port map (
            O => \N__69564\,
            I => \N__69551\
        );

    \I__16526\ : Span4Mux_h
    port map (
            O => \N__69561\,
            I => \N__69543\
        );

    \I__16525\ : Span4Mux_h
    port map (
            O => \N__69558\,
            I => \N__69540\
        );

    \I__16524\ : InMux
    port map (
            O => \N__69557\,
            I => \N__69537\
        );

    \I__16523\ : Span4Mux_v
    port map (
            O => \N__69554\,
            I => \N__69532\
        );

    \I__16522\ : Span4Mux_h
    port map (
            O => \N__69551\,
            I => \N__69532\
        );

    \I__16521\ : InMux
    port map (
            O => \N__69550\,
            I => \N__69525\
        );

    \I__16520\ : InMux
    port map (
            O => \N__69549\,
            I => \N__69525\
        );

    \I__16519\ : InMux
    port map (
            O => \N__69548\,
            I => \N__69525\
        );

    \I__16518\ : InMux
    port map (
            O => \N__69547\,
            I => \N__69522\
        );

    \I__16517\ : InMux
    port map (
            O => \N__69546\,
            I => \N__69519\
        );

    \I__16516\ : Odrv4
    port map (
            O => \N__69543\,
            I => \c0.data_in_frame_0_0\
        );

    \I__16515\ : Odrv4
    port map (
            O => \N__69540\,
            I => \c0.data_in_frame_0_0\
        );

    \I__16514\ : LocalMux
    port map (
            O => \N__69537\,
            I => \c0.data_in_frame_0_0\
        );

    \I__16513\ : Odrv4
    port map (
            O => \N__69532\,
            I => \c0.data_in_frame_0_0\
        );

    \I__16512\ : LocalMux
    port map (
            O => \N__69525\,
            I => \c0.data_in_frame_0_0\
        );

    \I__16511\ : LocalMux
    port map (
            O => \N__69522\,
            I => \c0.data_in_frame_0_0\
        );

    \I__16510\ : LocalMux
    port map (
            O => \N__69519\,
            I => \c0.data_in_frame_0_0\
        );

    \I__16509\ : CascadeMux
    port map (
            O => \N__69504\,
            I => \N__69501\
        );

    \I__16508\ : InMux
    port map (
            O => \N__69501\,
            I => \N__69495\
        );

    \I__16507\ : InMux
    port map (
            O => \N__69500\,
            I => \N__69495\
        );

    \I__16506\ : LocalMux
    port map (
            O => \N__69495\,
            I => \c0.n22701\
        );

    \I__16505\ : InMux
    port map (
            O => \N__69492\,
            I => \N__69488\
        );

    \I__16504\ : InMux
    port map (
            O => \N__69491\,
            I => \N__69485\
        );

    \I__16503\ : LocalMux
    port map (
            O => \N__69488\,
            I => \N__69482\
        );

    \I__16502\ : LocalMux
    port map (
            O => \N__69485\,
            I => \N__69475\
        );

    \I__16501\ : Span4Mux_h
    port map (
            O => \N__69482\,
            I => \N__69475\
        );

    \I__16500\ : InMux
    port map (
            O => \N__69481\,
            I => \N__69472\
        );

    \I__16499\ : InMux
    port map (
            O => \N__69480\,
            I => \N__69469\
        );

    \I__16498\ : Odrv4
    port map (
            O => \N__69475\,
            I => \c0.n5_adj_4323\
        );

    \I__16497\ : LocalMux
    port map (
            O => \N__69472\,
            I => \c0.n5_adj_4323\
        );

    \I__16496\ : LocalMux
    port map (
            O => \N__69469\,
            I => \c0.n5_adj_4323\
        );

    \I__16495\ : InMux
    port map (
            O => \N__69462\,
            I => \N__69454\
        );

    \I__16494\ : InMux
    port map (
            O => \N__69461\,
            I => \N__69454\
        );

    \I__16493\ : InMux
    port map (
            O => \N__69460\,
            I => \N__69451\
        );

    \I__16492\ : InMux
    port map (
            O => \N__69459\,
            I => \N__69447\
        );

    \I__16491\ : LocalMux
    port map (
            O => \N__69454\,
            I => \N__69444\
        );

    \I__16490\ : LocalMux
    port map (
            O => \N__69451\,
            I => \N__69441\
        );

    \I__16489\ : InMux
    port map (
            O => \N__69450\,
            I => \N__69438\
        );

    \I__16488\ : LocalMux
    port map (
            O => \N__69447\,
            I => \N__69434\
        );

    \I__16487\ : Span4Mux_h
    port map (
            O => \N__69444\,
            I => \N__69431\
        );

    \I__16486\ : Span4Mux_v
    port map (
            O => \N__69441\,
            I => \N__69426\
        );

    \I__16485\ : LocalMux
    port map (
            O => \N__69438\,
            I => \N__69426\
        );

    \I__16484\ : InMux
    port map (
            O => \N__69437\,
            I => \N__69423\
        );

    \I__16483\ : Span4Mux_h
    port map (
            O => \N__69434\,
            I => \N__69420\
        );

    \I__16482\ : Span4Mux_v
    port map (
            O => \N__69431\,
            I => \N__69415\
        );

    \I__16481\ : Span4Mux_h
    port map (
            O => \N__69426\,
            I => \N__69415\
        );

    \I__16480\ : LocalMux
    port map (
            O => \N__69423\,
            I => \N__69412\
        );

    \I__16479\ : Span4Mux_v
    port map (
            O => \N__69420\,
            I => \N__69407\
        );

    \I__16478\ : Span4Mux_h
    port map (
            O => \N__69415\,
            I => \N__69402\
        );

    \I__16477\ : Span4Mux_v
    port map (
            O => \N__69412\,
            I => \N__69402\
        );

    \I__16476\ : InMux
    port map (
            O => \N__69411\,
            I => \N__69399\
        );

    \I__16475\ : InMux
    port map (
            O => \N__69410\,
            I => \N__69396\
        );

    \I__16474\ : Odrv4
    port map (
            O => \N__69407\,
            I => n22101
        );

    \I__16473\ : Odrv4
    port map (
            O => \N__69402\,
            I => n22101
        );

    \I__16472\ : LocalMux
    port map (
            O => \N__69399\,
            I => n22101
        );

    \I__16471\ : LocalMux
    port map (
            O => \N__69396\,
            I => n22101
        );

    \I__16470\ : CascadeMux
    port map (
            O => \N__69387\,
            I => \c0.n9_cascade_\
        );

    \I__16469\ : CascadeMux
    port map (
            O => \N__69384\,
            I => \N__69381\
        );

    \I__16468\ : InMux
    port map (
            O => \N__69381\,
            I => \N__69377\
        );

    \I__16467\ : InMux
    port map (
            O => \N__69380\,
            I => \N__69373\
        );

    \I__16466\ : LocalMux
    port map (
            O => \N__69377\,
            I => \N__69370\
        );

    \I__16465\ : InMux
    port map (
            O => \N__69376\,
            I => \N__69367\
        );

    \I__16464\ : LocalMux
    port map (
            O => \N__69373\,
            I => \N__69364\
        );

    \I__16463\ : Span4Mux_v
    port map (
            O => \N__69370\,
            I => \N__69355\
        );

    \I__16462\ : LocalMux
    port map (
            O => \N__69367\,
            I => \N__69355\
        );

    \I__16461\ : Span4Mux_v
    port map (
            O => \N__69364\,
            I => \N__69355\
        );

    \I__16460\ : CascadeMux
    port map (
            O => \N__69363\,
            I => \N__69351\
        );

    \I__16459\ : CascadeMux
    port map (
            O => \N__69362\,
            I => \N__69348\
        );

    \I__16458\ : Span4Mux_v
    port map (
            O => \N__69355\,
            I => \N__69345\
        );

    \I__16457\ : InMux
    port map (
            O => \N__69354\,
            I => \N__69342\
        );

    \I__16456\ : InMux
    port map (
            O => \N__69351\,
            I => \N__69337\
        );

    \I__16455\ : InMux
    port map (
            O => \N__69348\,
            I => \N__69337\
        );

    \I__16454\ : Odrv4
    port map (
            O => \N__69345\,
            I => \c0.data_in_frame_9_1\
        );

    \I__16453\ : LocalMux
    port map (
            O => \N__69342\,
            I => \c0.data_in_frame_9_1\
        );

    \I__16452\ : LocalMux
    port map (
            O => \N__69337\,
            I => \c0.data_in_frame_9_1\
        );

    \I__16451\ : InMux
    port map (
            O => \N__69330\,
            I => \N__69326\
        );

    \I__16450\ : InMux
    port map (
            O => \N__69329\,
            I => \N__69322\
        );

    \I__16449\ : LocalMux
    port map (
            O => \N__69326\,
            I => \N__69317\
        );

    \I__16448\ : CascadeMux
    port map (
            O => \N__69325\,
            I => \N__69314\
        );

    \I__16447\ : LocalMux
    port map (
            O => \N__69322\,
            I => \N__69310\
        );

    \I__16446\ : InMux
    port map (
            O => \N__69321\,
            I => \N__69305\
        );

    \I__16445\ : InMux
    port map (
            O => \N__69320\,
            I => \N__69305\
        );

    \I__16444\ : Span4Mux_h
    port map (
            O => \N__69317\,
            I => \N__69302\
        );

    \I__16443\ : InMux
    port map (
            O => \N__69314\,
            I => \N__69298\
        );

    \I__16442\ : InMux
    port map (
            O => \N__69313\,
            I => \N__69295\
        );

    \I__16441\ : Span4Mux_h
    port map (
            O => \N__69310\,
            I => \N__69288\
        );

    \I__16440\ : LocalMux
    port map (
            O => \N__69305\,
            I => \N__69288\
        );

    \I__16439\ : Span4Mux_v
    port map (
            O => \N__69302\,
            I => \N__69288\
        );

    \I__16438\ : InMux
    port map (
            O => \N__69301\,
            I => \N__69285\
        );

    \I__16437\ : LocalMux
    port map (
            O => \N__69298\,
            I => \c0.data_in_frame_8_6\
        );

    \I__16436\ : LocalMux
    port map (
            O => \N__69295\,
            I => \c0.data_in_frame_8_6\
        );

    \I__16435\ : Odrv4
    port map (
            O => \N__69288\,
            I => \c0.data_in_frame_8_6\
        );

    \I__16434\ : LocalMux
    port map (
            O => \N__69285\,
            I => \c0.data_in_frame_8_6\
        );

    \I__16433\ : CascadeMux
    port map (
            O => \N__69276\,
            I => \N__69272\
        );

    \I__16432\ : InMux
    port map (
            O => \N__69275\,
            I => \N__69267\
        );

    \I__16431\ : InMux
    port map (
            O => \N__69272\,
            I => \N__69267\
        );

    \I__16430\ : LocalMux
    port map (
            O => \N__69267\,
            I => \c0.data_in_frame_18_0\
        );

    \I__16429\ : InMux
    port map (
            O => \N__69264\,
            I => \N__69255\
        );

    \I__16428\ : InMux
    port map (
            O => \N__69263\,
            I => \N__69255\
        );

    \I__16427\ : InMux
    port map (
            O => \N__69262\,
            I => \N__69255\
        );

    \I__16426\ : LocalMux
    port map (
            O => \N__69255\,
            I => data_in_frame_6_5
        );

    \I__16425\ : CascadeMux
    port map (
            O => \N__69252\,
            I => \N__69249\
        );

    \I__16424\ : InMux
    port map (
            O => \N__69249\,
            I => \N__69246\
        );

    \I__16423\ : LocalMux
    port map (
            O => \N__69246\,
            I => \N__69243\
        );

    \I__16422\ : Span4Mux_h
    port map (
            O => \N__69243\,
            I => \N__69240\
        );

    \I__16421\ : Odrv4
    port map (
            O => \N__69240\,
            I => \c0.n19_adj_4620\
        );

    \I__16420\ : InMux
    port map (
            O => \N__69237\,
            I => \N__69228\
        );

    \I__16419\ : InMux
    port map (
            O => \N__69236\,
            I => \N__69228\
        );

    \I__16418\ : InMux
    port map (
            O => \N__69235\,
            I => \N__69228\
        );

    \I__16417\ : LocalMux
    port map (
            O => \N__69228\,
            I => \N__69220\
        );

    \I__16416\ : InMux
    port map (
            O => \N__69227\,
            I => \N__69215\
        );

    \I__16415\ : InMux
    port map (
            O => \N__69226\,
            I => \N__69215\
        );

    \I__16414\ : CascadeMux
    port map (
            O => \N__69225\,
            I => \N__69212\
        );

    \I__16413\ : InMux
    port map (
            O => \N__69224\,
            I => \N__69205\
        );

    \I__16412\ : InMux
    port map (
            O => \N__69223\,
            I => \N__69205\
        );

    \I__16411\ : Span4Mux_v
    port map (
            O => \N__69220\,
            I => \N__69201\
        );

    \I__16410\ : LocalMux
    port map (
            O => \N__69215\,
            I => \N__69196\
        );

    \I__16409\ : InMux
    port map (
            O => \N__69212\,
            I => \N__69191\
        );

    \I__16408\ : InMux
    port map (
            O => \N__69211\,
            I => \N__69186\
        );

    \I__16407\ : InMux
    port map (
            O => \N__69210\,
            I => \N__69186\
        );

    \I__16406\ : LocalMux
    port map (
            O => \N__69205\,
            I => \N__69177\
        );

    \I__16405\ : InMux
    port map (
            O => \N__69204\,
            I => \N__69174\
        );

    \I__16404\ : Span4Mux_v
    port map (
            O => \N__69201\,
            I => \N__69171\
        );

    \I__16403\ : CascadeMux
    port map (
            O => \N__69200\,
            I => \N__69167\
        );

    \I__16402\ : CascadeMux
    port map (
            O => \N__69199\,
            I => \N__69163\
        );

    \I__16401\ : Span4Mux_v
    port map (
            O => \N__69196\,
            I => \N__69158\
        );

    \I__16400\ : InMux
    port map (
            O => \N__69195\,
            I => \N__69151\
        );

    \I__16399\ : InMux
    port map (
            O => \N__69194\,
            I => \N__69151\
        );

    \I__16398\ : LocalMux
    port map (
            O => \N__69191\,
            I => \N__69147\
        );

    \I__16397\ : LocalMux
    port map (
            O => \N__69186\,
            I => \N__69144\
        );

    \I__16396\ : InMux
    port map (
            O => \N__69185\,
            I => \N__69141\
        );

    \I__16395\ : InMux
    port map (
            O => \N__69184\,
            I => \N__69136\
        );

    \I__16394\ : InMux
    port map (
            O => \N__69183\,
            I => \N__69136\
        );

    \I__16393\ : InMux
    port map (
            O => \N__69182\,
            I => \N__69129\
        );

    \I__16392\ : InMux
    port map (
            O => \N__69181\,
            I => \N__69129\
        );

    \I__16391\ : InMux
    port map (
            O => \N__69180\,
            I => \N__69129\
        );

    \I__16390\ : Span4Mux_h
    port map (
            O => \N__69177\,
            I => \N__69124\
        );

    \I__16389\ : LocalMux
    port map (
            O => \N__69174\,
            I => \N__69124\
        );

    \I__16388\ : Span4Mux_h
    port map (
            O => \N__69171\,
            I => \N__69121\
        );

    \I__16387\ : CascadeMux
    port map (
            O => \N__69170\,
            I => \N__69118\
        );

    \I__16386\ : InMux
    port map (
            O => \N__69167\,
            I => \N__69112\
        );

    \I__16385\ : InMux
    port map (
            O => \N__69166\,
            I => \N__69112\
        );

    \I__16384\ : InMux
    port map (
            O => \N__69163\,
            I => \N__69109\
        );

    \I__16383\ : InMux
    port map (
            O => \N__69162\,
            I => \N__69104\
        );

    \I__16382\ : InMux
    port map (
            O => \N__69161\,
            I => \N__69104\
        );

    \I__16381\ : Sp12to4
    port map (
            O => \N__69158\,
            I => \N__69101\
        );

    \I__16380\ : InMux
    port map (
            O => \N__69157\,
            I => \N__69098\
        );

    \I__16379\ : InMux
    port map (
            O => \N__69156\,
            I => \N__69095\
        );

    \I__16378\ : LocalMux
    port map (
            O => \N__69151\,
            I => \N__69092\
        );

    \I__16377\ : InMux
    port map (
            O => \N__69150\,
            I => \N__69088\
        );

    \I__16376\ : Span4Mux_v
    port map (
            O => \N__69147\,
            I => \N__69085\
        );

    \I__16375\ : Span4Mux_v
    port map (
            O => \N__69144\,
            I => \N__69078\
        );

    \I__16374\ : LocalMux
    port map (
            O => \N__69141\,
            I => \N__69078\
        );

    \I__16373\ : LocalMux
    port map (
            O => \N__69136\,
            I => \N__69078\
        );

    \I__16372\ : LocalMux
    port map (
            O => \N__69129\,
            I => \N__69075\
        );

    \I__16371\ : Span4Mux_h
    port map (
            O => \N__69124\,
            I => \N__69072\
        );

    \I__16370\ : Sp12to4
    port map (
            O => \N__69121\,
            I => \N__69069\
        );

    \I__16369\ : InMux
    port map (
            O => \N__69118\,
            I => \N__69065\
        );

    \I__16368\ : InMux
    port map (
            O => \N__69117\,
            I => \N__69062\
        );

    \I__16367\ : LocalMux
    port map (
            O => \N__69112\,
            I => \N__69059\
        );

    \I__16366\ : LocalMux
    port map (
            O => \N__69109\,
            I => \N__69050\
        );

    \I__16365\ : LocalMux
    port map (
            O => \N__69104\,
            I => \N__69050\
        );

    \I__16364\ : Span12Mux_s9_v
    port map (
            O => \N__69101\,
            I => \N__69050\
        );

    \I__16363\ : LocalMux
    port map (
            O => \N__69098\,
            I => \N__69050\
        );

    \I__16362\ : LocalMux
    port map (
            O => \N__69095\,
            I => \N__69047\
        );

    \I__16361\ : Span4Mux_h
    port map (
            O => \N__69092\,
            I => \N__69044\
        );

    \I__16360\ : InMux
    port map (
            O => \N__69091\,
            I => \N__69041\
        );

    \I__16359\ : LocalMux
    port map (
            O => \N__69088\,
            I => \N__69038\
        );

    \I__16358\ : Span4Mux_h
    port map (
            O => \N__69085\,
            I => \N__69035\
        );

    \I__16357\ : Span4Mux_h
    port map (
            O => \N__69078\,
            I => \N__69032\
        );

    \I__16356\ : Sp12to4
    port map (
            O => \N__69075\,
            I => \N__69025\
        );

    \I__16355\ : Sp12to4
    port map (
            O => \N__69072\,
            I => \N__69025\
        );

    \I__16354\ : Span12Mux_h
    port map (
            O => \N__69069\,
            I => \N__69025\
        );

    \I__16353\ : InMux
    port map (
            O => \N__69068\,
            I => \N__69022\
        );

    \I__16352\ : LocalMux
    port map (
            O => \N__69065\,
            I => \N__69019\
        );

    \I__16351\ : LocalMux
    port map (
            O => \N__69062\,
            I => \N__69012\
        );

    \I__16350\ : Span12Mux_s10_v
    port map (
            O => \N__69059\,
            I => \N__69012\
        );

    \I__16349\ : Span12Mux_v
    port map (
            O => \N__69050\,
            I => \N__69012\
        );

    \I__16348\ : Span4Mux_h
    port map (
            O => \N__69047\,
            I => \N__69007\
        );

    \I__16347\ : Span4Mux_v
    port map (
            O => \N__69044\,
            I => \N__69007\
        );

    \I__16346\ : LocalMux
    port map (
            O => \N__69041\,
            I => \N__69000\
        );

    \I__16345\ : Span4Mux_v
    port map (
            O => \N__69038\,
            I => \N__69000\
        );

    \I__16344\ : Span4Mux_v
    port map (
            O => \N__69035\,
            I => \N__69000\
        );

    \I__16343\ : Sp12to4
    port map (
            O => \N__69032\,
            I => \N__68995\
        );

    \I__16342\ : Span12Mux_v
    port map (
            O => \N__69025\,
            I => \N__68995\
        );

    \I__16341\ : LocalMux
    port map (
            O => \N__69022\,
            I => \c0.n9\
        );

    \I__16340\ : Odrv4
    port map (
            O => \N__69019\,
            I => \c0.n9\
        );

    \I__16339\ : Odrv12
    port map (
            O => \N__69012\,
            I => \c0.n9\
        );

    \I__16338\ : Odrv4
    port map (
            O => \N__69007\,
            I => \c0.n9\
        );

    \I__16337\ : Odrv4
    port map (
            O => \N__69000\,
            I => \c0.n9\
        );

    \I__16336\ : Odrv12
    port map (
            O => \N__68995\,
            I => \c0.n9\
        );

    \I__16335\ : InMux
    port map (
            O => \N__68982\,
            I => \N__68979\
        );

    \I__16334\ : LocalMux
    port map (
            O => \N__68979\,
            I => \N__68976\
        );

    \I__16333\ : Span4Mux_v
    port map (
            O => \N__68976\,
            I => \N__68973\
        );

    \I__16332\ : Odrv4
    port map (
            O => \N__68973\,
            I => \c0.n22392\
        );

    \I__16331\ : InMux
    port map (
            O => \N__68970\,
            I => \N__68966\
        );

    \I__16330\ : CascadeMux
    port map (
            O => \N__68969\,
            I => \N__68963\
        );

    \I__16329\ : LocalMux
    port map (
            O => \N__68966\,
            I => \N__68960\
        );

    \I__16328\ : InMux
    port map (
            O => \N__68963\,
            I => \N__68954\
        );

    \I__16327\ : Span4Mux_h
    port map (
            O => \N__68960\,
            I => \N__68951\
        );

    \I__16326\ : InMux
    port map (
            O => \N__68959\,
            I => \N__68948\
        );

    \I__16325\ : InMux
    port map (
            O => \N__68958\,
            I => \N__68945\
        );

    \I__16324\ : InMux
    port map (
            O => \N__68957\,
            I => \N__68942\
        );

    \I__16323\ : LocalMux
    port map (
            O => \N__68954\,
            I => \c0.data_in_frame_4_3\
        );

    \I__16322\ : Odrv4
    port map (
            O => \N__68951\,
            I => \c0.data_in_frame_4_3\
        );

    \I__16321\ : LocalMux
    port map (
            O => \N__68948\,
            I => \c0.data_in_frame_4_3\
        );

    \I__16320\ : LocalMux
    port map (
            O => \N__68945\,
            I => \c0.data_in_frame_4_3\
        );

    \I__16319\ : LocalMux
    port map (
            O => \N__68942\,
            I => \c0.data_in_frame_4_3\
        );

    \I__16318\ : CascadeMux
    port map (
            O => \N__68931\,
            I => \c0.n6_adj_4687_cascade_\
        );

    \I__16317\ : InMux
    port map (
            O => \N__68928\,
            I => \N__68924\
        );

    \I__16316\ : CascadeMux
    port map (
            O => \N__68927\,
            I => \N__68920\
        );

    \I__16315\ : LocalMux
    port map (
            O => \N__68924\,
            I => \N__68917\
        );

    \I__16314\ : InMux
    port map (
            O => \N__68923\,
            I => \N__68914\
        );

    \I__16313\ : InMux
    port map (
            O => \N__68920\,
            I => \N__68911\
        );

    \I__16312\ : Span4Mux_v
    port map (
            O => \N__68917\,
            I => \N__68908\
        );

    \I__16311\ : LocalMux
    port map (
            O => \N__68914\,
            I => \c0.n23274\
        );

    \I__16310\ : LocalMux
    port map (
            O => \N__68911\,
            I => \c0.n23274\
        );

    \I__16309\ : Odrv4
    port map (
            O => \N__68908\,
            I => \c0.n23274\
        );

    \I__16308\ : InMux
    port map (
            O => \N__68901\,
            I => \N__68895\
        );

    \I__16307\ : InMux
    port map (
            O => \N__68900\,
            I => \N__68895\
        );

    \I__16306\ : LocalMux
    port map (
            O => \N__68895\,
            I => \c0.n23282\
        );

    \I__16305\ : CascadeMux
    port map (
            O => \N__68892\,
            I => \c0.n23274_cascade_\
        );

    \I__16304\ : InMux
    port map (
            O => \N__68889\,
            I => \N__68886\
        );

    \I__16303\ : LocalMux
    port map (
            O => \N__68886\,
            I => \c0.n20_adj_4316\
        );

    \I__16302\ : InMux
    port map (
            O => \N__68883\,
            I => \N__68880\
        );

    \I__16301\ : LocalMux
    port map (
            O => \N__68880\,
            I => \N__68876\
        );

    \I__16300\ : CascadeMux
    port map (
            O => \N__68879\,
            I => \N__68873\
        );

    \I__16299\ : Span4Mux_v
    port map (
            O => \N__68876\,
            I => \N__68870\
        );

    \I__16298\ : InMux
    port map (
            O => \N__68873\,
            I => \N__68867\
        );

    \I__16297\ : Span4Mux_h
    port map (
            O => \N__68870\,
            I => \N__68864\
        );

    \I__16296\ : LocalMux
    port map (
            O => \N__68867\,
            I => \N__68861\
        );

    \I__16295\ : Span4Mux_v
    port map (
            O => \N__68864\,
            I => \N__68858\
        );

    \I__16294\ : Span12Mux_h
    port map (
            O => \N__68861\,
            I => \N__68855\
        );

    \I__16293\ : Odrv4
    port map (
            O => \N__68858\,
            I => \c0.n29_adj_4287\
        );

    \I__16292\ : Odrv12
    port map (
            O => \N__68855\,
            I => \c0.n29_adj_4287\
        );

    \I__16291\ : InMux
    port map (
            O => \N__68850\,
            I => \N__68837\
        );

    \I__16290\ : InMux
    port map (
            O => \N__68849\,
            I => \N__68832\
        );

    \I__16289\ : InMux
    port map (
            O => \N__68848\,
            I => \N__68832\
        );

    \I__16288\ : InMux
    port map (
            O => \N__68847\,
            I => \N__68829\
        );

    \I__16287\ : InMux
    port map (
            O => \N__68846\,
            I => \N__68826\
        );

    \I__16286\ : InMux
    port map (
            O => \N__68845\,
            I => \N__68821\
        );

    \I__16285\ : InMux
    port map (
            O => \N__68844\,
            I => \N__68821\
        );

    \I__16284\ : InMux
    port map (
            O => \N__68843\,
            I => \N__68814\
        );

    \I__16283\ : InMux
    port map (
            O => \N__68842\,
            I => \N__68814\
        );

    \I__16282\ : InMux
    port map (
            O => \N__68841\,
            I => \N__68814\
        );

    \I__16281\ : InMux
    port map (
            O => \N__68840\,
            I => \N__68811\
        );

    \I__16280\ : LocalMux
    port map (
            O => \N__68837\,
            I => \c0.data_in_frame_0_2\
        );

    \I__16279\ : LocalMux
    port map (
            O => \N__68832\,
            I => \c0.data_in_frame_0_2\
        );

    \I__16278\ : LocalMux
    port map (
            O => \N__68829\,
            I => \c0.data_in_frame_0_2\
        );

    \I__16277\ : LocalMux
    port map (
            O => \N__68826\,
            I => \c0.data_in_frame_0_2\
        );

    \I__16276\ : LocalMux
    port map (
            O => \N__68821\,
            I => \c0.data_in_frame_0_2\
        );

    \I__16275\ : LocalMux
    port map (
            O => \N__68814\,
            I => \c0.data_in_frame_0_2\
        );

    \I__16274\ : LocalMux
    port map (
            O => \N__68811\,
            I => \c0.data_in_frame_0_2\
        );

    \I__16273\ : CascadeMux
    port map (
            O => \N__68796\,
            I => \N__68790\
        );

    \I__16272\ : InMux
    port map (
            O => \N__68795\,
            I => \N__68787\
        );

    \I__16271\ : InMux
    port map (
            O => \N__68794\,
            I => \N__68782\
        );

    \I__16270\ : InMux
    port map (
            O => \N__68793\,
            I => \N__68782\
        );

    \I__16269\ : InMux
    port map (
            O => \N__68790\,
            I => \N__68777\
        );

    \I__16268\ : LocalMux
    port map (
            O => \N__68787\,
            I => \N__68774\
        );

    \I__16267\ : LocalMux
    port map (
            O => \N__68782\,
            I => \N__68771\
        );

    \I__16266\ : InMux
    port map (
            O => \N__68781\,
            I => \N__68766\
        );

    \I__16265\ : InMux
    port map (
            O => \N__68780\,
            I => \N__68766\
        );

    \I__16264\ : LocalMux
    port map (
            O => \N__68777\,
            I => \c0.data_in_frame_2_3\
        );

    \I__16263\ : Odrv4
    port map (
            O => \N__68774\,
            I => \c0.data_in_frame_2_3\
        );

    \I__16262\ : Odrv4
    port map (
            O => \N__68771\,
            I => \c0.data_in_frame_2_3\
        );

    \I__16261\ : LocalMux
    port map (
            O => \N__68766\,
            I => \c0.data_in_frame_2_3\
        );

    \I__16260\ : InMux
    port map (
            O => \N__68757\,
            I => \N__68753\
        );

    \I__16259\ : CascadeMux
    port map (
            O => \N__68756\,
            I => \N__68746\
        );

    \I__16258\ : LocalMux
    port map (
            O => \N__68753\,
            I => \N__68743\
        );

    \I__16257\ : InMux
    port map (
            O => \N__68752\,
            I => \N__68740\
        );

    \I__16256\ : InMux
    port map (
            O => \N__68751\,
            I => \N__68737\
        );

    \I__16255\ : InMux
    port map (
            O => \N__68750\,
            I => \N__68734\
        );

    \I__16254\ : CascadeMux
    port map (
            O => \N__68749\,
            I => \N__68729\
        );

    \I__16253\ : InMux
    port map (
            O => \N__68746\,
            I => \N__68723\
        );

    \I__16252\ : Span4Mux_h
    port map (
            O => \N__68743\,
            I => \N__68716\
        );

    \I__16251\ : LocalMux
    port map (
            O => \N__68740\,
            I => \N__68716\
        );

    \I__16250\ : LocalMux
    port map (
            O => \N__68737\,
            I => \N__68716\
        );

    \I__16249\ : LocalMux
    port map (
            O => \N__68734\,
            I => \N__68713\
        );

    \I__16248\ : InMux
    port map (
            O => \N__68733\,
            I => \N__68710\
        );

    \I__16247\ : InMux
    port map (
            O => \N__68732\,
            I => \N__68707\
        );

    \I__16246\ : InMux
    port map (
            O => \N__68729\,
            I => \N__68702\
        );

    \I__16245\ : InMux
    port map (
            O => \N__68728\,
            I => \N__68702\
        );

    \I__16244\ : InMux
    port map (
            O => \N__68727\,
            I => \N__68699\
        );

    \I__16243\ : InMux
    port map (
            O => \N__68726\,
            I => \N__68696\
        );

    \I__16242\ : LocalMux
    port map (
            O => \N__68723\,
            I => \c0.data_in_frame_0_1\
        );

    \I__16241\ : Odrv4
    port map (
            O => \N__68716\,
            I => \c0.data_in_frame_0_1\
        );

    \I__16240\ : Odrv4
    port map (
            O => \N__68713\,
            I => \c0.data_in_frame_0_1\
        );

    \I__16239\ : LocalMux
    port map (
            O => \N__68710\,
            I => \c0.data_in_frame_0_1\
        );

    \I__16238\ : LocalMux
    port map (
            O => \N__68707\,
            I => \c0.data_in_frame_0_1\
        );

    \I__16237\ : LocalMux
    port map (
            O => \N__68702\,
            I => \c0.data_in_frame_0_1\
        );

    \I__16236\ : LocalMux
    port map (
            O => \N__68699\,
            I => \c0.data_in_frame_0_1\
        );

    \I__16235\ : LocalMux
    port map (
            O => \N__68696\,
            I => \c0.data_in_frame_0_1\
        );

    \I__16234\ : InMux
    port map (
            O => \N__68679\,
            I => \N__68672\
        );

    \I__16233\ : InMux
    port map (
            O => \N__68678\,
            I => \N__68672\
        );

    \I__16232\ : InMux
    port map (
            O => \N__68677\,
            I => \N__68666\
        );

    \I__16231\ : LocalMux
    port map (
            O => \N__68672\,
            I => \N__68663\
        );

    \I__16230\ : InMux
    port map (
            O => \N__68671\,
            I => \N__68660\
        );

    \I__16229\ : InMux
    port map (
            O => \N__68670\,
            I => \N__68655\
        );

    \I__16228\ : InMux
    port map (
            O => \N__68669\,
            I => \N__68655\
        );

    \I__16227\ : LocalMux
    port map (
            O => \N__68666\,
            I => \c0.data_in_frame_4_4\
        );

    \I__16226\ : Odrv12
    port map (
            O => \N__68663\,
            I => \c0.data_in_frame_4_4\
        );

    \I__16225\ : LocalMux
    port map (
            O => \N__68660\,
            I => \c0.data_in_frame_4_4\
        );

    \I__16224\ : LocalMux
    port map (
            O => \N__68655\,
            I => \c0.data_in_frame_4_4\
        );

    \I__16223\ : InMux
    port map (
            O => \N__68646\,
            I => \N__68642\
        );

    \I__16222\ : InMux
    port map (
            O => \N__68645\,
            I => \N__68639\
        );

    \I__16221\ : LocalMux
    port map (
            O => \N__68642\,
            I => \c0.n23276\
        );

    \I__16220\ : LocalMux
    port map (
            O => \N__68639\,
            I => \c0.n23276\
        );

    \I__16219\ : InMux
    port map (
            O => \N__68634\,
            I => \N__68628\
        );

    \I__16218\ : InMux
    port map (
            O => \N__68633\,
            I => \N__68628\
        );

    \I__16217\ : LocalMux
    port map (
            O => \N__68628\,
            I => \N__68625\
        );

    \I__16216\ : Span4Mux_v
    port map (
            O => \N__68625\,
            I => \N__68619\
        );

    \I__16215\ : InMux
    port map (
            O => \N__68624\,
            I => \N__68612\
        );

    \I__16214\ : InMux
    port map (
            O => \N__68623\,
            I => \N__68612\
        );

    \I__16213\ : InMux
    port map (
            O => \N__68622\,
            I => \N__68612\
        );

    \I__16212\ : Odrv4
    port map (
            O => \N__68619\,
            I => \c0.n22322\
        );

    \I__16211\ : LocalMux
    port map (
            O => \N__68612\,
            I => \c0.n22322\
        );

    \I__16210\ : CascadeMux
    port map (
            O => \N__68607\,
            I => \c0.n23276_cascade_\
        );

    \I__16209\ : InMux
    port map (
            O => \N__68604\,
            I => \N__68601\
        );

    \I__16208\ : LocalMux
    port map (
            O => \N__68601\,
            I => \N__68597\
        );

    \I__16207\ : InMux
    port map (
            O => \N__68600\,
            I => \N__68594\
        );

    \I__16206\ : Span4Mux_v
    port map (
            O => \N__68597\,
            I => \N__68588\
        );

    \I__16205\ : LocalMux
    port map (
            O => \N__68594\,
            I => \N__68588\
        );

    \I__16204\ : InMux
    port map (
            O => \N__68593\,
            I => \N__68585\
        );

    \I__16203\ : Span4Mux_h
    port map (
            O => \N__68588\,
            I => \N__68582\
        );

    \I__16202\ : LocalMux
    port map (
            O => \N__68585\,
            I => \N__68579\
        );

    \I__16201\ : Span4Mux_h
    port map (
            O => \N__68582\,
            I => \N__68576\
        );

    \I__16200\ : Odrv4
    port map (
            O => \N__68579\,
            I => \c0.n25\
        );

    \I__16199\ : Odrv4
    port map (
            O => \N__68576\,
            I => \c0.n25\
        );

    \I__16198\ : InMux
    port map (
            O => \N__68571\,
            I => \N__68567\
        );

    \I__16197\ : InMux
    port map (
            O => \N__68570\,
            I => \N__68564\
        );

    \I__16196\ : LocalMux
    port map (
            O => \N__68567\,
            I => \c0.n24_adj_4213\
        );

    \I__16195\ : LocalMux
    port map (
            O => \N__68564\,
            I => \c0.n24_adj_4213\
        );

    \I__16194\ : CascadeMux
    port map (
            O => \N__68559\,
            I => \c0.n8_cascade_\
        );

    \I__16193\ : InMux
    port map (
            O => \N__68556\,
            I => \N__68552\
        );

    \I__16192\ : CascadeMux
    port map (
            O => \N__68555\,
            I => \N__68549\
        );

    \I__16191\ : LocalMux
    port map (
            O => \N__68552\,
            I => \N__68546\
        );

    \I__16190\ : InMux
    port map (
            O => \N__68549\,
            I => \N__68539\
        );

    \I__16189\ : Span4Mux_h
    port map (
            O => \N__68546\,
            I => \N__68536\
        );

    \I__16188\ : InMux
    port map (
            O => \N__68545\,
            I => \N__68533\
        );

    \I__16187\ : InMux
    port map (
            O => \N__68544\,
            I => \N__68528\
        );

    \I__16186\ : CascadeMux
    port map (
            O => \N__68543\,
            I => \N__68524\
        );

    \I__16185\ : CascadeMux
    port map (
            O => \N__68542\,
            I => \N__68521\
        );

    \I__16184\ : LocalMux
    port map (
            O => \N__68539\,
            I => \N__68518\
        );

    \I__16183\ : Span4Mux_v
    port map (
            O => \N__68536\,
            I => \N__68513\
        );

    \I__16182\ : LocalMux
    port map (
            O => \N__68533\,
            I => \N__68513\
        );

    \I__16181\ : InMux
    port map (
            O => \N__68532\,
            I => \N__68507\
        );

    \I__16180\ : InMux
    port map (
            O => \N__68531\,
            I => \N__68504\
        );

    \I__16179\ : LocalMux
    port map (
            O => \N__68528\,
            I => \N__68501\
        );

    \I__16178\ : InMux
    port map (
            O => \N__68527\,
            I => \N__68498\
        );

    \I__16177\ : InMux
    port map (
            O => \N__68524\,
            I => \N__68490\
        );

    \I__16176\ : InMux
    port map (
            O => \N__68521\,
            I => \N__68490\
        );

    \I__16175\ : Span4Mux_v
    port map (
            O => \N__68518\,
            I => \N__68485\
        );

    \I__16174\ : Span4Mux_v
    port map (
            O => \N__68513\,
            I => \N__68485\
        );

    \I__16173\ : InMux
    port map (
            O => \N__68512\,
            I => \N__68482\
        );

    \I__16172\ : InMux
    port map (
            O => \N__68511\,
            I => \N__68477\
        );

    \I__16171\ : InMux
    port map (
            O => \N__68510\,
            I => \N__68477\
        );

    \I__16170\ : LocalMux
    port map (
            O => \N__68507\,
            I => \N__68472\
        );

    \I__16169\ : LocalMux
    port map (
            O => \N__68504\,
            I => \N__68472\
        );

    \I__16168\ : Span4Mux_v
    port map (
            O => \N__68501\,
            I => \N__68467\
        );

    \I__16167\ : LocalMux
    port map (
            O => \N__68498\,
            I => \N__68467\
        );

    \I__16166\ : InMux
    port map (
            O => \N__68497\,
            I => \N__68464\
        );

    \I__16165\ : InMux
    port map (
            O => \N__68496\,
            I => \N__68459\
        );

    \I__16164\ : InMux
    port map (
            O => \N__68495\,
            I => \N__68459\
        );

    \I__16163\ : LocalMux
    port map (
            O => \N__68490\,
            I => \c0.data_in_frame_0_4\
        );

    \I__16162\ : Odrv4
    port map (
            O => \N__68485\,
            I => \c0.data_in_frame_0_4\
        );

    \I__16161\ : LocalMux
    port map (
            O => \N__68482\,
            I => \c0.data_in_frame_0_4\
        );

    \I__16160\ : LocalMux
    port map (
            O => \N__68477\,
            I => \c0.data_in_frame_0_4\
        );

    \I__16159\ : Odrv4
    port map (
            O => \N__68472\,
            I => \c0.data_in_frame_0_4\
        );

    \I__16158\ : Odrv4
    port map (
            O => \N__68467\,
            I => \c0.data_in_frame_0_4\
        );

    \I__16157\ : LocalMux
    port map (
            O => \N__68464\,
            I => \c0.data_in_frame_0_4\
        );

    \I__16156\ : LocalMux
    port map (
            O => \N__68459\,
            I => \c0.data_in_frame_0_4\
        );

    \I__16155\ : InMux
    port map (
            O => \N__68442\,
            I => \N__68438\
        );

    \I__16154\ : InMux
    port map (
            O => \N__68441\,
            I => \N__68434\
        );

    \I__16153\ : LocalMux
    port map (
            O => \N__68438\,
            I => \N__68429\
        );

    \I__16152\ : InMux
    port map (
            O => \N__68437\,
            I => \N__68426\
        );

    \I__16151\ : LocalMux
    port map (
            O => \N__68434\,
            I => \N__68423\
        );

    \I__16150\ : InMux
    port map (
            O => \N__68433\,
            I => \N__68419\
        );

    \I__16149\ : InMux
    port map (
            O => \N__68432\,
            I => \N__68416\
        );

    \I__16148\ : Span4Mux_h
    port map (
            O => \N__68429\,
            I => \N__68411\
        );

    \I__16147\ : LocalMux
    port map (
            O => \N__68426\,
            I => \N__68411\
        );

    \I__16146\ : Span4Mux_v
    port map (
            O => \N__68423\,
            I => \N__68408\
        );

    \I__16145\ : InMux
    port map (
            O => \N__68422\,
            I => \N__68405\
        );

    \I__16144\ : LocalMux
    port map (
            O => \N__68419\,
            I => \N__68402\
        );

    \I__16143\ : LocalMux
    port map (
            O => \N__68416\,
            I => \N__68399\
        );

    \I__16142\ : Span4Mux_h
    port map (
            O => \N__68411\,
            I => \N__68396\
        );

    \I__16141\ : Sp12to4
    port map (
            O => \N__68408\,
            I => \N__68390\
        );

    \I__16140\ : LocalMux
    port map (
            O => \N__68405\,
            I => \N__68390\
        );

    \I__16139\ : Span12Mux_h
    port map (
            O => \N__68402\,
            I => \N__68387\
        );

    \I__16138\ : Span4Mux_h
    port map (
            O => \N__68399\,
            I => \N__68382\
        );

    \I__16137\ : Span4Mux_h
    port map (
            O => \N__68396\,
            I => \N__68382\
        );

    \I__16136\ : InMux
    port map (
            O => \N__68395\,
            I => \N__68379\
        );

    \I__16135\ : Odrv12
    port map (
            O => \N__68390\,
            I => n22121
        );

    \I__16134\ : Odrv12
    port map (
            O => \N__68387\,
            I => n22121
        );

    \I__16133\ : Odrv4
    port map (
            O => \N__68382\,
            I => n22121
        );

    \I__16132\ : LocalMux
    port map (
            O => \N__68379\,
            I => n22121
        );

    \I__16131\ : InMux
    port map (
            O => \N__68370\,
            I => \N__68367\
        );

    \I__16130\ : LocalMux
    port map (
            O => \N__68367\,
            I => \N__68362\
        );

    \I__16129\ : InMux
    port map (
            O => \N__68366\,
            I => \N__68359\
        );

    \I__16128\ : InMux
    port map (
            O => \N__68365\,
            I => \N__68356\
        );

    \I__16127\ : Span4Mux_v
    port map (
            O => \N__68362\,
            I => \N__68353\
        );

    \I__16126\ : LocalMux
    port map (
            O => \N__68359\,
            I => \N__68350\
        );

    \I__16125\ : LocalMux
    port map (
            O => \N__68356\,
            I => \N__68346\
        );

    \I__16124\ : Span4Mux_h
    port map (
            O => \N__68353\,
            I => \N__68343\
        );

    \I__16123\ : Span4Mux_v
    port map (
            O => \N__68350\,
            I => \N__68340\
        );

    \I__16122\ : InMux
    port map (
            O => \N__68349\,
            I => \N__68337\
        );

    \I__16121\ : Span12Mux_h
    port map (
            O => \N__68346\,
            I => \N__68334\
        );

    \I__16120\ : Span4Mux_h
    port map (
            O => \N__68343\,
            I => \N__68331\
        );

    \I__16119\ : Span4Mux_h
    port map (
            O => \N__68340\,
            I => \N__68328\
        );

    \I__16118\ : LocalMux
    port map (
            O => \N__68337\,
            I => \c0.data_in_frame_26_3\
        );

    \I__16117\ : Odrv12
    port map (
            O => \N__68334\,
            I => \c0.data_in_frame_26_3\
        );

    \I__16116\ : Odrv4
    port map (
            O => \N__68331\,
            I => \c0.data_in_frame_26_3\
        );

    \I__16115\ : Odrv4
    port map (
            O => \N__68328\,
            I => \c0.data_in_frame_26_3\
        );

    \I__16114\ : CascadeMux
    port map (
            O => \N__68319\,
            I => \c0.n22362_cascade_\
        );

    \I__16113\ : InMux
    port map (
            O => \N__68316\,
            I => \N__68313\
        );

    \I__16112\ : LocalMux
    port map (
            O => \N__68313\,
            I => \N__68308\
        );

    \I__16111\ : InMux
    port map (
            O => \N__68312\,
            I => \N__68305\
        );

    \I__16110\ : InMux
    port map (
            O => \N__68311\,
            I => \N__68302\
        );

    \I__16109\ : Odrv4
    port map (
            O => \N__68308\,
            I => \c0.n12559\
        );

    \I__16108\ : LocalMux
    port map (
            O => \N__68305\,
            I => \c0.n12559\
        );

    \I__16107\ : LocalMux
    port map (
            O => \N__68302\,
            I => \c0.n12559\
        );

    \I__16106\ : CascadeMux
    port map (
            O => \N__68295\,
            I => \N__68292\
        );

    \I__16105\ : InMux
    port map (
            O => \N__68292\,
            I => \N__68289\
        );

    \I__16104\ : LocalMux
    port map (
            O => \N__68289\,
            I => \N__68286\
        );

    \I__16103\ : Span4Mux_h
    port map (
            O => \N__68286\,
            I => \N__68283\
        );

    \I__16102\ : Odrv4
    port map (
            O => \N__68283\,
            I => \c0.n13_adj_4527\
        );

    \I__16101\ : InMux
    port map (
            O => \N__68280\,
            I => \N__68275\
        );

    \I__16100\ : InMux
    port map (
            O => \N__68279\,
            I => \N__68270\
        );

    \I__16099\ : InMux
    port map (
            O => \N__68278\,
            I => \N__68270\
        );

    \I__16098\ : LocalMux
    port map (
            O => \N__68275\,
            I => \N__68267\
        );

    \I__16097\ : LocalMux
    port map (
            O => \N__68270\,
            I => \c0.n20802\
        );

    \I__16096\ : Odrv4
    port map (
            O => \N__68267\,
            I => \c0.n20802\
        );

    \I__16095\ : InMux
    port map (
            O => \N__68262\,
            I => \N__68258\
        );

    \I__16094\ : InMux
    port map (
            O => \N__68261\,
            I => \N__68255\
        );

    \I__16093\ : LocalMux
    port map (
            O => \N__68258\,
            I => \N__68252\
        );

    \I__16092\ : LocalMux
    port map (
            O => \N__68255\,
            I => \c0.n20358\
        );

    \I__16091\ : Odrv12
    port map (
            O => \N__68252\,
            I => \c0.n20358\
        );

    \I__16090\ : InMux
    port map (
            O => \N__68247\,
            I => \N__68244\
        );

    \I__16089\ : LocalMux
    port map (
            O => \N__68244\,
            I => \c0.n12_adj_4491\
        );

    \I__16088\ : CascadeMux
    port map (
            O => \N__68241\,
            I => \N__68237\
        );

    \I__16087\ : InMux
    port map (
            O => \N__68240\,
            I => \N__68232\
        );

    \I__16086\ : InMux
    port map (
            O => \N__68237\,
            I => \N__68232\
        );

    \I__16085\ : LocalMux
    port map (
            O => \N__68232\,
            I => \c0.data_in_frame_28_6\
        );

    \I__16084\ : InMux
    port map (
            O => \N__68229\,
            I => \N__68223\
        );

    \I__16083\ : InMux
    port map (
            O => \N__68228\,
            I => \N__68223\
        );

    \I__16082\ : LocalMux
    port map (
            O => \N__68223\,
            I => \N__68220\
        );

    \I__16081\ : Odrv4
    port map (
            O => \N__68220\,
            I => \c0.data_in_frame_28_4\
        );

    \I__16080\ : InMux
    port map (
            O => \N__68217\,
            I => \N__68212\
        );

    \I__16079\ : CascadeMux
    port map (
            O => \N__68216\,
            I => \N__68209\
        );

    \I__16078\ : InMux
    port map (
            O => \N__68215\,
            I => \N__68206\
        );

    \I__16077\ : LocalMux
    port map (
            O => \N__68212\,
            I => \N__68203\
        );

    \I__16076\ : InMux
    port map (
            O => \N__68209\,
            I => \N__68200\
        );

    \I__16075\ : LocalMux
    port map (
            O => \N__68206\,
            I => \N__68197\
        );

    \I__16074\ : Odrv12
    port map (
            O => \N__68203\,
            I => \c0.n13904\
        );

    \I__16073\ : LocalMux
    port map (
            O => \N__68200\,
            I => \c0.n13904\
        );

    \I__16072\ : Odrv4
    port map (
            O => \N__68197\,
            I => \c0.n13904\
        );

    \I__16071\ : InMux
    port map (
            O => \N__68190\,
            I => \N__68186\
        );

    \I__16070\ : InMux
    port map (
            O => \N__68189\,
            I => \N__68183\
        );

    \I__16069\ : LocalMux
    port map (
            O => \N__68186\,
            I => \N__68180\
        );

    \I__16068\ : LocalMux
    port map (
            O => \N__68183\,
            I => \N__68177\
        );

    \I__16067\ : Span4Mux_h
    port map (
            O => \N__68180\,
            I => \N__68174\
        );

    \I__16066\ : Sp12to4
    port map (
            O => \N__68177\,
            I => \N__68171\
        );

    \I__16065\ : Span4Mux_v
    port map (
            O => \N__68174\,
            I => \N__68168\
        );

    \I__16064\ : Odrv12
    port map (
            O => \N__68171\,
            I => \c0.n28_adj_4286\
        );

    \I__16063\ : Odrv4
    port map (
            O => \N__68168\,
            I => \c0.n28_adj_4286\
        );

    \I__16062\ : InMux
    port map (
            O => \N__68163\,
            I => \N__68157\
        );

    \I__16061\ : InMux
    port map (
            O => \N__68162\,
            I => \N__68150\
        );

    \I__16060\ : InMux
    port map (
            O => \N__68161\,
            I => \N__68150\
        );

    \I__16059\ : InMux
    port map (
            O => \N__68160\,
            I => \N__68150\
        );

    \I__16058\ : LocalMux
    port map (
            O => \N__68157\,
            I => data_in_frame_5_0
        );

    \I__16057\ : LocalMux
    port map (
            O => \N__68150\,
            I => data_in_frame_5_0
        );

    \I__16056\ : InMux
    port map (
            O => \N__68145\,
            I => \N__68142\
        );

    \I__16055\ : LocalMux
    port map (
            O => \N__68142\,
            I => \N__68137\
        );

    \I__16054\ : InMux
    port map (
            O => \N__68141\,
            I => \N__68132\
        );

    \I__16053\ : InMux
    port map (
            O => \N__68140\,
            I => \N__68132\
        );

    \I__16052\ : Odrv4
    port map (
            O => \N__68137\,
            I => \c0.n23302\
        );

    \I__16051\ : LocalMux
    port map (
            O => \N__68132\,
            I => \c0.n23302\
        );

    \I__16050\ : InMux
    port map (
            O => \N__68127\,
            I => \N__68123\
        );

    \I__16049\ : InMux
    port map (
            O => \N__68126\,
            I => \N__68117\
        );

    \I__16048\ : LocalMux
    port map (
            O => \N__68123\,
            I => \N__68114\
        );

    \I__16047\ : InMux
    port map (
            O => \N__68122\,
            I => \N__68111\
        );

    \I__16046\ : CascadeMux
    port map (
            O => \N__68121\,
            I => \N__68105\
        );

    \I__16045\ : InMux
    port map (
            O => \N__68120\,
            I => \N__68102\
        );

    \I__16044\ : LocalMux
    port map (
            O => \N__68117\,
            I => \N__68097\
        );

    \I__16043\ : Span4Mux_v
    port map (
            O => \N__68114\,
            I => \N__68097\
        );

    \I__16042\ : LocalMux
    port map (
            O => \N__68111\,
            I => \N__68090\
        );

    \I__16041\ : InMux
    port map (
            O => \N__68110\,
            I => \N__68083\
        );

    \I__16040\ : InMux
    port map (
            O => \N__68109\,
            I => \N__68083\
        );

    \I__16039\ : InMux
    port map (
            O => \N__68108\,
            I => \N__68083\
        );

    \I__16038\ : InMux
    port map (
            O => \N__68105\,
            I => \N__68078\
        );

    \I__16037\ : LocalMux
    port map (
            O => \N__68102\,
            I => \N__68073\
        );

    \I__16036\ : Span4Mux_h
    port map (
            O => \N__68097\,
            I => \N__68073\
        );

    \I__16035\ : InMux
    port map (
            O => \N__68096\,
            I => \N__68068\
        );

    \I__16034\ : InMux
    port map (
            O => \N__68095\,
            I => \N__68068\
        );

    \I__16033\ : InMux
    port map (
            O => \N__68094\,
            I => \N__68063\
        );

    \I__16032\ : InMux
    port map (
            O => \N__68093\,
            I => \N__68063\
        );

    \I__16031\ : Span4Mux_h
    port map (
            O => \N__68090\,
            I => \N__68058\
        );

    \I__16030\ : LocalMux
    port map (
            O => \N__68083\,
            I => \N__68058\
        );

    \I__16029\ : InMux
    port map (
            O => \N__68082\,
            I => \N__68053\
        );

    \I__16028\ : InMux
    port map (
            O => \N__68081\,
            I => \N__68053\
        );

    \I__16027\ : LocalMux
    port map (
            O => \N__68078\,
            I => \c0.data_in_frame_0_3\
        );

    \I__16026\ : Odrv4
    port map (
            O => \N__68073\,
            I => \c0.data_in_frame_0_3\
        );

    \I__16025\ : LocalMux
    port map (
            O => \N__68068\,
            I => \c0.data_in_frame_0_3\
        );

    \I__16024\ : LocalMux
    port map (
            O => \N__68063\,
            I => \c0.data_in_frame_0_3\
        );

    \I__16023\ : Odrv4
    port map (
            O => \N__68058\,
            I => \c0.data_in_frame_0_3\
        );

    \I__16022\ : LocalMux
    port map (
            O => \N__68053\,
            I => \c0.data_in_frame_0_3\
        );

    \I__16021\ : CascadeMux
    port map (
            O => \N__68040\,
            I => \N__68035\
        );

    \I__16020\ : CascadeMux
    port map (
            O => \N__68039\,
            I => \N__68031\
        );

    \I__16019\ : InMux
    port map (
            O => \N__68038\,
            I => \N__68025\
        );

    \I__16018\ : InMux
    port map (
            O => \N__68035\,
            I => \N__68022\
        );

    \I__16017\ : InMux
    port map (
            O => \N__68034\,
            I => \N__68019\
        );

    \I__16016\ : InMux
    port map (
            O => \N__68031\,
            I => \N__68014\
        );

    \I__16015\ : InMux
    port map (
            O => \N__68030\,
            I => \N__68014\
        );

    \I__16014\ : InMux
    port map (
            O => \N__68029\,
            I => \N__68009\
        );

    \I__16013\ : InMux
    port map (
            O => \N__68028\,
            I => \N__68009\
        );

    \I__16012\ : LocalMux
    port map (
            O => \N__68025\,
            I => \c0.data_in_frame_2_4\
        );

    \I__16011\ : LocalMux
    port map (
            O => \N__68022\,
            I => \c0.data_in_frame_2_4\
        );

    \I__16010\ : LocalMux
    port map (
            O => \N__68019\,
            I => \c0.data_in_frame_2_4\
        );

    \I__16009\ : LocalMux
    port map (
            O => \N__68014\,
            I => \c0.data_in_frame_2_4\
        );

    \I__16008\ : LocalMux
    port map (
            O => \N__68009\,
            I => \c0.data_in_frame_2_4\
        );

    \I__16007\ : InMux
    port map (
            O => \N__67998\,
            I => \N__67995\
        );

    \I__16006\ : LocalMux
    port map (
            O => \N__67995\,
            I => \N__67992\
        );

    \I__16005\ : Span12Mux_h
    port map (
            O => \N__67992\,
            I => \N__67989\
        );

    \I__16004\ : Odrv12
    port map (
            O => \N__67989\,
            I => \c0.n42_adj_4746\
        );

    \I__16003\ : InMux
    port map (
            O => \N__67986\,
            I => \N__67981\
        );

    \I__16002\ : InMux
    port map (
            O => \N__67985\,
            I => \N__67978\
        );

    \I__16001\ : CascadeMux
    port map (
            O => \N__67984\,
            I => \N__67975\
        );

    \I__16000\ : LocalMux
    port map (
            O => \N__67981\,
            I => \N__67972\
        );

    \I__15999\ : LocalMux
    port map (
            O => \N__67978\,
            I => \N__67969\
        );

    \I__15998\ : InMux
    port map (
            O => \N__67975\,
            I => \N__67964\
        );

    \I__15997\ : Span4Mux_v
    port map (
            O => \N__67972\,
            I => \N__67959\
        );

    \I__15996\ : Span4Mux_h
    port map (
            O => \N__67969\,
            I => \N__67959\
        );

    \I__15995\ : InMux
    port map (
            O => \N__67968\,
            I => \N__67956\
        );

    \I__15994\ : InMux
    port map (
            O => \N__67967\,
            I => \N__67953\
        );

    \I__15993\ : LocalMux
    port map (
            O => \N__67964\,
            I => \c0.data_in_frame_7_1\
        );

    \I__15992\ : Odrv4
    port map (
            O => \N__67959\,
            I => \c0.data_in_frame_7_1\
        );

    \I__15991\ : LocalMux
    port map (
            O => \N__67956\,
            I => \c0.data_in_frame_7_1\
        );

    \I__15990\ : LocalMux
    port map (
            O => \N__67953\,
            I => \c0.data_in_frame_7_1\
        );

    \I__15989\ : CascadeMux
    port map (
            O => \N__67944\,
            I => \N__67938\
        );

    \I__15988\ : CascadeMux
    port map (
            O => \N__67943\,
            I => \N__67935\
        );

    \I__15987\ : InMux
    port map (
            O => \N__67942\,
            I => \N__67931\
        );

    \I__15986\ : InMux
    port map (
            O => \N__67941\,
            I => \N__67928\
        );

    \I__15985\ : InMux
    port map (
            O => \N__67938\,
            I => \N__67925\
        );

    \I__15984\ : InMux
    port map (
            O => \N__67935\,
            I => \N__67922\
        );

    \I__15983\ : InMux
    port map (
            O => \N__67934\,
            I => \N__67919\
        );

    \I__15982\ : LocalMux
    port map (
            O => \N__67931\,
            I => \N__67916\
        );

    \I__15981\ : LocalMux
    port map (
            O => \N__67928\,
            I => \N__67911\
        );

    \I__15980\ : LocalMux
    port map (
            O => \N__67925\,
            I => \N__67908\
        );

    \I__15979\ : LocalMux
    port map (
            O => \N__67922\,
            I => \N__67903\
        );

    \I__15978\ : LocalMux
    port map (
            O => \N__67919\,
            I => \N__67903\
        );

    \I__15977\ : Span4Mux_h
    port map (
            O => \N__67916\,
            I => \N__67900\
        );

    \I__15976\ : InMux
    port map (
            O => \N__67915\,
            I => \N__67895\
        );

    \I__15975\ : InMux
    port map (
            O => \N__67914\,
            I => \N__67895\
        );

    \I__15974\ : Odrv4
    port map (
            O => \N__67911\,
            I => \c0.data_in_frame_2_5\
        );

    \I__15973\ : Odrv4
    port map (
            O => \N__67908\,
            I => \c0.data_in_frame_2_5\
        );

    \I__15972\ : Odrv4
    port map (
            O => \N__67903\,
            I => \c0.data_in_frame_2_5\
        );

    \I__15971\ : Odrv4
    port map (
            O => \N__67900\,
            I => \c0.data_in_frame_2_5\
        );

    \I__15970\ : LocalMux
    port map (
            O => \N__67895\,
            I => \c0.data_in_frame_2_5\
        );

    \I__15969\ : InMux
    port map (
            O => \N__67884\,
            I => \N__67880\
        );

    \I__15968\ : InMux
    port map (
            O => \N__67883\,
            I => \N__67877\
        );

    \I__15967\ : LocalMux
    port map (
            O => \N__67880\,
            I => \N__67874\
        );

    \I__15966\ : LocalMux
    port map (
            O => \N__67877\,
            I => \N__67870\
        );

    \I__15965\ : Span4Mux_v
    port map (
            O => \N__67874\,
            I => \N__67867\
        );

    \I__15964\ : CascadeMux
    port map (
            O => \N__67873\,
            I => \N__67864\
        );

    \I__15963\ : Span4Mux_v
    port map (
            O => \N__67870\,
            I => \N__67859\
        );

    \I__15962\ : Sp12to4
    port map (
            O => \N__67867\,
            I => \N__67856\
        );

    \I__15961\ : InMux
    port map (
            O => \N__67864\,
            I => \N__67853\
        );

    \I__15960\ : CascadeMux
    port map (
            O => \N__67863\,
            I => \N__67850\
        );

    \I__15959\ : InMux
    port map (
            O => \N__67862\,
            I => \N__67847\
        );

    \I__15958\ : Span4Mux_h
    port map (
            O => \N__67859\,
            I => \N__67844\
        );

    \I__15957\ : Span12Mux_h
    port map (
            O => \N__67856\,
            I => \N__67841\
        );

    \I__15956\ : LocalMux
    port map (
            O => \N__67853\,
            I => \N__67838\
        );

    \I__15955\ : InMux
    port map (
            O => \N__67850\,
            I => \N__67835\
        );

    \I__15954\ : LocalMux
    port map (
            O => \N__67847\,
            I => \c0.data_in_frame_27_2\
        );

    \I__15953\ : Odrv4
    port map (
            O => \N__67844\,
            I => \c0.data_in_frame_27_2\
        );

    \I__15952\ : Odrv12
    port map (
            O => \N__67841\,
            I => \c0.data_in_frame_27_2\
        );

    \I__15951\ : Odrv12
    port map (
            O => \N__67838\,
            I => \c0.data_in_frame_27_2\
        );

    \I__15950\ : LocalMux
    port map (
            O => \N__67835\,
            I => \c0.data_in_frame_27_2\
        );

    \I__15949\ : InMux
    port map (
            O => \N__67824\,
            I => \N__67821\
        );

    \I__15948\ : LocalMux
    port map (
            O => \N__67821\,
            I => \N__67816\
        );

    \I__15947\ : InMux
    port map (
            O => \N__67820\,
            I => \N__67813\
        );

    \I__15946\ : InMux
    port map (
            O => \N__67819\,
            I => \N__67810\
        );

    \I__15945\ : Span4Mux_v
    port map (
            O => \N__67816\,
            I => \N__67805\
        );

    \I__15944\ : LocalMux
    port map (
            O => \N__67813\,
            I => \N__67805\
        );

    \I__15943\ : LocalMux
    port map (
            O => \N__67810\,
            I => \N__67802\
        );

    \I__15942\ : Odrv4
    port map (
            O => \N__67805\,
            I => \c0.n25_adj_4469\
        );

    \I__15941\ : Odrv4
    port map (
            O => \N__67802\,
            I => \c0.n25_adj_4469\
        );

    \I__15940\ : InMux
    port map (
            O => \N__67797\,
            I => \N__67794\
        );

    \I__15939\ : LocalMux
    port map (
            O => \N__67794\,
            I => \N__67789\
        );

    \I__15938\ : InMux
    port map (
            O => \N__67793\,
            I => \N__67786\
        );

    \I__15937\ : InMux
    port map (
            O => \N__67792\,
            I => \N__67783\
        );

    \I__15936\ : Span4Mux_h
    port map (
            O => \N__67789\,
            I => \N__67780\
        );

    \I__15935\ : LocalMux
    port map (
            O => \N__67786\,
            I => \c0.n26_adj_4470\
        );

    \I__15934\ : LocalMux
    port map (
            O => \N__67783\,
            I => \c0.n26_adj_4470\
        );

    \I__15933\ : Odrv4
    port map (
            O => \N__67780\,
            I => \c0.n26_adj_4470\
        );

    \I__15932\ : InMux
    port map (
            O => \N__67773\,
            I => \N__67770\
        );

    \I__15931\ : LocalMux
    port map (
            O => \N__67770\,
            I => \c0.n39_adj_4467\
        );

    \I__15930\ : InMux
    port map (
            O => \N__67767\,
            I => \N__67764\
        );

    \I__15929\ : LocalMux
    port map (
            O => \N__67764\,
            I => \c0.n38_adj_4468\
        );

    \I__15928\ : InMux
    port map (
            O => \N__67761\,
            I => \N__67758\
        );

    \I__15927\ : LocalMux
    port map (
            O => \N__67758\,
            I => \N__67755\
        );

    \I__15926\ : Odrv4
    port map (
            O => \N__67755\,
            I => \c0.n37_adj_4473\
        );

    \I__15925\ : CascadeMux
    port map (
            O => \N__67752\,
            I => \c0.n44_adj_4471_cascade_\
        );

    \I__15924\ : InMux
    port map (
            O => \N__67749\,
            I => \N__67745\
        );

    \I__15923\ : InMux
    port map (
            O => \N__67748\,
            I => \N__67742\
        );

    \I__15922\ : LocalMux
    port map (
            O => \N__67745\,
            I => \N__67739\
        );

    \I__15921\ : LocalMux
    port map (
            O => \N__67742\,
            I => \N__67736\
        );

    \I__15920\ : Span4Mux_v
    port map (
            O => \N__67739\,
            I => \N__67733\
        );

    \I__15919\ : Span4Mux_v
    port map (
            O => \N__67736\,
            I => \N__67730\
        );

    \I__15918\ : Odrv4
    port map (
            O => \N__67733\,
            I => \c0.n45_adj_4476\
        );

    \I__15917\ : Odrv4
    port map (
            O => \N__67730\,
            I => \c0.n45_adj_4476\
        );

    \I__15916\ : InMux
    port map (
            O => \N__67725\,
            I => \N__67722\
        );

    \I__15915\ : LocalMux
    port map (
            O => \N__67722\,
            I => \N__67719\
        );

    \I__15914\ : Odrv12
    port map (
            O => \N__67719\,
            I => \c0.n14_adj_4529\
        );

    \I__15913\ : InMux
    port map (
            O => \N__67716\,
            I => \N__67713\
        );

    \I__15912\ : LocalMux
    port map (
            O => \N__67713\,
            I => \N__67710\
        );

    \I__15911\ : Span4Mux_h
    port map (
            O => \N__67710\,
            I => \N__67707\
        );

    \I__15910\ : Span4Mux_v
    port map (
            O => \N__67707\,
            I => \N__67703\
        );

    \I__15909\ : InMux
    port map (
            O => \N__67706\,
            I => \N__67700\
        );

    \I__15908\ : Odrv4
    port map (
            O => \N__67703\,
            I => \c0.n15_adj_4508\
        );

    \I__15907\ : LocalMux
    port map (
            O => \N__67700\,
            I => \c0.n15_adj_4508\
        );

    \I__15906\ : CascadeMux
    port map (
            O => \N__67695\,
            I => \c0.n24362_cascade_\
        );

    \I__15905\ : InMux
    port map (
            O => \N__67692\,
            I => \N__67689\
        );

    \I__15904\ : LocalMux
    port map (
            O => \N__67689\,
            I => \N__67686\
        );

    \I__15903\ : Span4Mux_h
    port map (
            O => \N__67686\,
            I => \N__67683\
        );

    \I__15902\ : Odrv4
    port map (
            O => \N__67683\,
            I => \c0.n18_adj_4475\
        );

    \I__15901\ : InMux
    port map (
            O => \N__67680\,
            I => \N__67677\
        );

    \I__15900\ : LocalMux
    port map (
            O => \N__67677\,
            I => \N__67674\
        );

    \I__15899\ : Span4Mux_v
    port map (
            O => \N__67674\,
            I => \N__67671\
        );

    \I__15898\ : Span4Mux_h
    port map (
            O => \N__67671\,
            I => \N__67668\
        );

    \I__15897\ : Odrv4
    port map (
            O => \N__67668\,
            I => \c0.n26_adj_4530\
        );

    \I__15896\ : InMux
    port map (
            O => \N__67665\,
            I => \N__67661\
        );

    \I__15895\ : InMux
    port map (
            O => \N__67664\,
            I => \N__67658\
        );

    \I__15894\ : LocalMux
    port map (
            O => \N__67661\,
            I => \N__67652\
        );

    \I__15893\ : LocalMux
    port map (
            O => \N__67658\,
            I => \N__67652\
        );

    \I__15892\ : InMux
    port map (
            O => \N__67657\,
            I => \N__67649\
        );

    \I__15891\ : Span4Mux_v
    port map (
            O => \N__67652\,
            I => \N__67645\
        );

    \I__15890\ : LocalMux
    port map (
            O => \N__67649\,
            I => \N__67641\
        );

    \I__15889\ : InMux
    port map (
            O => \N__67648\,
            I => \N__67637\
        );

    \I__15888\ : Span4Mux_h
    port map (
            O => \N__67645\,
            I => \N__67634\
        );

    \I__15887\ : InMux
    port map (
            O => \N__67644\,
            I => \N__67631\
        );

    \I__15886\ : Span4Mux_h
    port map (
            O => \N__67641\,
            I => \N__67628\
        );

    \I__15885\ : InMux
    port map (
            O => \N__67640\,
            I => \N__67625\
        );

    \I__15884\ : LocalMux
    port map (
            O => \N__67637\,
            I => \N__67622\
        );

    \I__15883\ : Span4Mux_v
    port map (
            O => \N__67634\,
            I => \N__67617\
        );

    \I__15882\ : LocalMux
    port map (
            O => \N__67631\,
            I => \N__67614\
        );

    \I__15881\ : Span4Mux_h
    port map (
            O => \N__67628\,
            I => \N__67607\
        );

    \I__15880\ : LocalMux
    port map (
            O => \N__67625\,
            I => \N__67607\
        );

    \I__15879\ : Span4Mux_h
    port map (
            O => \N__67622\,
            I => \N__67607\
        );

    \I__15878\ : InMux
    port map (
            O => \N__67621\,
            I => \N__67602\
        );

    \I__15877\ : InMux
    port map (
            O => \N__67620\,
            I => \N__67602\
        );

    \I__15876\ : Odrv4
    port map (
            O => \N__67617\,
            I => n22103
        );

    \I__15875\ : Odrv4
    port map (
            O => \N__67614\,
            I => n22103
        );

    \I__15874\ : Odrv4
    port map (
            O => \N__67607\,
            I => n22103
        );

    \I__15873\ : LocalMux
    port map (
            O => \N__67602\,
            I => n22103
        );

    \I__15872\ : InMux
    port map (
            O => \N__67593\,
            I => \N__67588\
        );

    \I__15871\ : InMux
    port map (
            O => \N__67592\,
            I => \N__67585\
        );

    \I__15870\ : InMux
    port map (
            O => \N__67591\,
            I => \N__67582\
        );

    \I__15869\ : LocalMux
    port map (
            O => \N__67588\,
            I => \N__67577\
        );

    \I__15868\ : LocalMux
    port map (
            O => \N__67585\,
            I => \N__67577\
        );

    \I__15867\ : LocalMux
    port map (
            O => \N__67582\,
            I => \N__67574\
        );

    \I__15866\ : Span4Mux_v
    port map (
            O => \N__67577\,
            I => \N__67571\
        );

    \I__15865\ : Odrv4
    port map (
            O => \N__67574\,
            I => \c0.n22632\
        );

    \I__15864\ : Odrv4
    port map (
            O => \N__67571\,
            I => \c0.n22632\
        );

    \I__15863\ : CascadeMux
    port map (
            O => \N__67566\,
            I => \c0.n22632_cascade_\
        );

    \I__15862\ : InMux
    port map (
            O => \N__67563\,
            I => \N__67560\
        );

    \I__15861\ : LocalMux
    port map (
            O => \N__67560\,
            I => \N__67556\
        );

    \I__15860\ : InMux
    port map (
            O => \N__67559\,
            I => \N__67553\
        );

    \I__15859\ : Span4Mux_v
    port map (
            O => \N__67556\,
            I => \N__67544\
        );

    \I__15858\ : LocalMux
    port map (
            O => \N__67553\,
            I => \N__67544\
        );

    \I__15857\ : InMux
    port map (
            O => \N__67552\,
            I => \N__67539\
        );

    \I__15856\ : InMux
    port map (
            O => \N__67551\,
            I => \N__67539\
        );

    \I__15855\ : InMux
    port map (
            O => \N__67550\,
            I => \N__67536\
        );

    \I__15854\ : InMux
    port map (
            O => \N__67549\,
            I => \N__67533\
        );

    \I__15853\ : Span4Mux_h
    port map (
            O => \N__67544\,
            I => \N__67529\
        );

    \I__15852\ : LocalMux
    port map (
            O => \N__67539\,
            I => \N__67522\
        );

    \I__15851\ : LocalMux
    port map (
            O => \N__67536\,
            I => \N__67522\
        );

    \I__15850\ : LocalMux
    port map (
            O => \N__67533\,
            I => \N__67522\
        );

    \I__15849\ : InMux
    port map (
            O => \N__67532\,
            I => \N__67519\
        );

    \I__15848\ : Span4Mux_h
    port map (
            O => \N__67529\,
            I => \N__67516\
        );

    \I__15847\ : Span12Mux_h
    port map (
            O => \N__67522\,
            I => \N__67513\
        );

    \I__15846\ : LocalMux
    port map (
            O => \N__67519\,
            I => \c0.data_in_frame_24_2\
        );

    \I__15845\ : Odrv4
    port map (
            O => \N__67516\,
            I => \c0.data_in_frame_24_2\
        );

    \I__15844\ : Odrv12
    port map (
            O => \N__67513\,
            I => \c0.data_in_frame_24_2\
        );

    \I__15843\ : InMux
    port map (
            O => \N__67506\,
            I => \N__67502\
        );

    \I__15842\ : InMux
    port map (
            O => \N__67505\,
            I => \N__67496\
        );

    \I__15841\ : LocalMux
    port map (
            O => \N__67502\,
            I => \N__67493\
        );

    \I__15840\ : InMux
    port map (
            O => \N__67501\,
            I => \N__67488\
        );

    \I__15839\ : InMux
    port map (
            O => \N__67500\,
            I => \N__67483\
        );

    \I__15838\ : InMux
    port map (
            O => \N__67499\,
            I => \N__67483\
        );

    \I__15837\ : LocalMux
    port map (
            O => \N__67496\,
            I => \N__67480\
        );

    \I__15836\ : Span4Mux_h
    port map (
            O => \N__67493\,
            I => \N__67477\
        );

    \I__15835\ : InMux
    port map (
            O => \N__67492\,
            I => \N__67472\
        );

    \I__15834\ : InMux
    port map (
            O => \N__67491\,
            I => \N__67472\
        );

    \I__15833\ : LocalMux
    port map (
            O => \N__67488\,
            I => \c0.n21316\
        );

    \I__15832\ : LocalMux
    port map (
            O => \N__67483\,
            I => \c0.n21316\
        );

    \I__15831\ : Odrv12
    port map (
            O => \N__67480\,
            I => \c0.n21316\
        );

    \I__15830\ : Odrv4
    port map (
            O => \N__67477\,
            I => \c0.n21316\
        );

    \I__15829\ : LocalMux
    port map (
            O => \N__67472\,
            I => \c0.n21316\
        );

    \I__15828\ : InMux
    port map (
            O => \N__67461\,
            I => \N__67458\
        );

    \I__15827\ : LocalMux
    port map (
            O => \N__67458\,
            I => \c0.n39_adj_4487\
        );

    \I__15826\ : CascadeMux
    port map (
            O => \N__67455\,
            I => \c0.n30_adj_4489_cascade_\
        );

    \I__15825\ : InMux
    port map (
            O => \N__67452\,
            I => \N__67449\
        );

    \I__15824\ : LocalMux
    port map (
            O => \N__67449\,
            I => \c0.n23209\
        );

    \I__15823\ : CascadeMux
    port map (
            O => \N__67446\,
            I => \c0.n45_adj_4490_cascade_\
        );

    \I__15822\ : InMux
    port map (
            O => \N__67443\,
            I => \N__67440\
        );

    \I__15821\ : LocalMux
    port map (
            O => \N__67440\,
            I => \N__67437\
        );

    \I__15820\ : Odrv4
    port map (
            O => \N__67437\,
            I => \c0.n44_adj_4501\
        );

    \I__15819\ : InMux
    port map (
            O => \N__67434\,
            I => \N__67431\
        );

    \I__15818\ : LocalMux
    port map (
            O => \N__67431\,
            I => \N__67428\
        );

    \I__15817\ : Span4Mux_h
    port map (
            O => \N__67428\,
            I => \N__67425\
        );

    \I__15816\ : Odrv4
    port map (
            O => \N__67425\,
            I => \c0.n11_adj_4505\
        );

    \I__15815\ : CascadeMux
    port map (
            O => \N__67422\,
            I => \c0.n48_adj_4503_cascade_\
        );

    \I__15814\ : InMux
    port map (
            O => \N__67419\,
            I => \N__67416\
        );

    \I__15813\ : LocalMux
    port map (
            O => \N__67416\,
            I => \N__67412\
        );

    \I__15812\ : CascadeMux
    port map (
            O => \N__67415\,
            I => \N__67409\
        );

    \I__15811\ : Span4Mux_h
    port map (
            O => \N__67412\,
            I => \N__67406\
        );

    \I__15810\ : InMux
    port map (
            O => \N__67409\,
            I => \N__67403\
        );

    \I__15809\ : Odrv4
    port map (
            O => \N__67406\,
            I => \c0.n28_adj_4504\
        );

    \I__15808\ : LocalMux
    port map (
            O => \N__67403\,
            I => \c0.n28_adj_4504\
        );

    \I__15807\ : InMux
    port map (
            O => \N__67398\,
            I => \N__67395\
        );

    \I__15806\ : LocalMux
    port map (
            O => \N__67395\,
            I => \N__67392\
        );

    \I__15805\ : Span4Mux_v
    port map (
            O => \N__67392\,
            I => \N__67389\
        );

    \I__15804\ : Odrv4
    port map (
            O => \N__67389\,
            I => \c0.n24573\
        );

    \I__15803\ : InMux
    port map (
            O => \N__67386\,
            I => \N__67383\
        );

    \I__15802\ : LocalMux
    port map (
            O => \N__67383\,
            I => \c0.n41_adj_4488\
        );

    \I__15801\ : InMux
    port map (
            O => \N__67380\,
            I => \N__67377\
        );

    \I__15800\ : LocalMux
    port map (
            O => \N__67377\,
            I => \N__67373\
        );

    \I__15799\ : InMux
    port map (
            O => \N__67376\,
            I => \N__67370\
        );

    \I__15798\ : Span4Mux_v
    port map (
            O => \N__67373\,
            I => \N__67365\
        );

    \I__15797\ : LocalMux
    port map (
            O => \N__67370\,
            I => \N__67365\
        );

    \I__15796\ : Odrv4
    port map (
            O => \N__67365\,
            I => \c0.n17_adj_4354\
        );

    \I__15795\ : InMux
    port map (
            O => \N__67362\,
            I => \N__67358\
        );

    \I__15794\ : InMux
    port map (
            O => \N__67361\,
            I => \N__67355\
        );

    \I__15793\ : LocalMux
    port map (
            O => \N__67358\,
            I => \N__67352\
        );

    \I__15792\ : LocalMux
    port map (
            O => \N__67355\,
            I => \N__67348\
        );

    \I__15791\ : Span4Mux_h
    port map (
            O => \N__67352\,
            I => \N__67345\
        );

    \I__15790\ : InMux
    port map (
            O => \N__67351\,
            I => \N__67342\
        );

    \I__15789\ : Odrv4
    port map (
            O => \N__67348\,
            I => \c0.n28_adj_4343\
        );

    \I__15788\ : Odrv4
    port map (
            O => \N__67345\,
            I => \c0.n28_adj_4343\
        );

    \I__15787\ : LocalMux
    port map (
            O => \N__67342\,
            I => \c0.n28_adj_4343\
        );

    \I__15786\ : InMux
    port map (
            O => \N__67335\,
            I => \N__67332\
        );

    \I__15785\ : LocalMux
    port map (
            O => \N__67332\,
            I => \c0.n27_adj_4502\
        );

    \I__15784\ : CascadeMux
    port map (
            O => \N__67329\,
            I => \N__67324\
        );

    \I__15783\ : InMux
    port map (
            O => \N__67328\,
            I => \N__67321\
        );

    \I__15782\ : CascadeMux
    port map (
            O => \N__67327\,
            I => \N__67318\
        );

    \I__15781\ : InMux
    port map (
            O => \N__67324\,
            I => \N__67315\
        );

    \I__15780\ : LocalMux
    port map (
            O => \N__67321\,
            I => \N__67310\
        );

    \I__15779\ : InMux
    port map (
            O => \N__67318\,
            I => \N__67307\
        );

    \I__15778\ : LocalMux
    port map (
            O => \N__67315\,
            I => \N__67304\
        );

    \I__15777\ : InMux
    port map (
            O => \N__67314\,
            I => \N__67301\
        );

    \I__15776\ : InMux
    port map (
            O => \N__67313\,
            I => \N__67298\
        );

    \I__15775\ : Span4Mux_h
    port map (
            O => \N__67310\,
            I => \N__67287\
        );

    \I__15774\ : LocalMux
    port map (
            O => \N__67307\,
            I => \N__67287\
        );

    \I__15773\ : Span4Mux_h
    port map (
            O => \N__67304\,
            I => \N__67287\
        );

    \I__15772\ : LocalMux
    port map (
            O => \N__67301\,
            I => \N__67287\
        );

    \I__15771\ : LocalMux
    port map (
            O => \N__67298\,
            I => \N__67284\
        );

    \I__15770\ : InMux
    port map (
            O => \N__67297\,
            I => \N__67281\
        );

    \I__15769\ : InMux
    port map (
            O => \N__67296\,
            I => \N__67278\
        );

    \I__15768\ : Span4Mux_h
    port map (
            O => \N__67287\,
            I => \N__67275\
        );

    \I__15767\ : Span12Mux_h
    port map (
            O => \N__67284\,
            I => \N__67272\
        );

    \I__15766\ : LocalMux
    port map (
            O => \N__67281\,
            I => \N__67269\
        );

    \I__15765\ : LocalMux
    port map (
            O => \N__67278\,
            I => \c0.data_in_frame_26_7\
        );

    \I__15764\ : Odrv4
    port map (
            O => \N__67275\,
            I => \c0.data_in_frame_26_7\
        );

    \I__15763\ : Odrv12
    port map (
            O => \N__67272\,
            I => \c0.data_in_frame_26_7\
        );

    \I__15762\ : Odrv12
    port map (
            O => \N__67269\,
            I => \c0.data_in_frame_26_7\
        );

    \I__15761\ : InMux
    port map (
            O => \N__67260\,
            I => \N__67257\
        );

    \I__15760\ : LocalMux
    port map (
            O => \N__67257\,
            I => \N__67252\
        );

    \I__15759\ : InMux
    port map (
            O => \N__67256\,
            I => \N__67243\
        );

    \I__15758\ : InMux
    port map (
            O => \N__67255\,
            I => \N__67243\
        );

    \I__15757\ : Span4Mux_v
    port map (
            O => \N__67252\,
            I => \N__67240\
        );

    \I__15756\ : InMux
    port map (
            O => \N__67251\,
            I => \N__67235\
        );

    \I__15755\ : InMux
    port map (
            O => \N__67250\,
            I => \N__67235\
        );

    \I__15754\ : InMux
    port map (
            O => \N__67249\,
            I => \N__67230\
        );

    \I__15753\ : InMux
    port map (
            O => \N__67248\,
            I => \N__67230\
        );

    \I__15752\ : LocalMux
    port map (
            O => \N__67243\,
            I => \N__67223\
        );

    \I__15751\ : Sp12to4
    port map (
            O => \N__67240\,
            I => \N__67223\
        );

    \I__15750\ : LocalMux
    port map (
            O => \N__67235\,
            I => \N__67223\
        );

    \I__15749\ : LocalMux
    port map (
            O => \N__67230\,
            I => \c0.data_in_frame_24_4\
        );

    \I__15748\ : Odrv12
    port map (
            O => \N__67223\,
            I => \c0.data_in_frame_24_4\
        );

    \I__15747\ : CascadeMux
    port map (
            O => \N__67218\,
            I => \N__67215\
        );

    \I__15746\ : InMux
    port map (
            O => \N__67215\,
            I => \N__67209\
        );

    \I__15745\ : InMux
    port map (
            O => \N__67214\,
            I => \N__67204\
        );

    \I__15744\ : InMux
    port map (
            O => \N__67213\,
            I => \N__67204\
        );

    \I__15743\ : InMux
    port map (
            O => \N__67212\,
            I => \N__67201\
        );

    \I__15742\ : LocalMux
    port map (
            O => \N__67209\,
            I => data_in_frame_21_6
        );

    \I__15741\ : LocalMux
    port map (
            O => \N__67204\,
            I => data_in_frame_21_6
        );

    \I__15740\ : LocalMux
    port map (
            O => \N__67201\,
            I => data_in_frame_21_6
        );

    \I__15739\ : InMux
    port map (
            O => \N__67194\,
            I => \N__67190\
        );

    \I__15738\ : InMux
    port map (
            O => \N__67193\,
            I => \N__67187\
        );

    \I__15737\ : LocalMux
    port map (
            O => \N__67190\,
            I => \N__67184\
        );

    \I__15736\ : LocalMux
    port map (
            O => \N__67187\,
            I => \N__67181\
        );

    \I__15735\ : Span4Mux_v
    port map (
            O => \N__67184\,
            I => \N__67177\
        );

    \I__15734\ : Span4Mux_v
    port map (
            O => \N__67181\,
            I => \N__67174\
        );

    \I__15733\ : InMux
    port map (
            O => \N__67180\,
            I => \N__67171\
        );

    \I__15732\ : Odrv4
    port map (
            O => \N__67177\,
            I => \c0.n21301\
        );

    \I__15731\ : Odrv4
    port map (
            O => \N__67174\,
            I => \c0.n21301\
        );

    \I__15730\ : LocalMux
    port map (
            O => \N__67171\,
            I => \c0.n21301\
        );

    \I__15729\ : InMux
    port map (
            O => \N__67164\,
            I => \N__67160\
        );

    \I__15728\ : InMux
    port map (
            O => \N__67163\,
            I => \N__67157\
        );

    \I__15727\ : LocalMux
    port map (
            O => \N__67160\,
            I => \c0.n23_adj_4582\
        );

    \I__15726\ : LocalMux
    port map (
            O => \N__67157\,
            I => \c0.n23_adj_4582\
        );

    \I__15725\ : CascadeMux
    port map (
            O => \N__67152\,
            I => \N__67144\
        );

    \I__15724\ : InMux
    port map (
            O => \N__67151\,
            I => \N__67141\
        );

    \I__15723\ : CascadeMux
    port map (
            O => \N__67150\,
            I => \N__67137\
        );

    \I__15722\ : InMux
    port map (
            O => \N__67149\,
            I => \N__67128\
        );

    \I__15721\ : InMux
    port map (
            O => \N__67148\,
            I => \N__67128\
        );

    \I__15720\ : InMux
    port map (
            O => \N__67147\,
            I => \N__67128\
        );

    \I__15719\ : InMux
    port map (
            O => \N__67144\,
            I => \N__67128\
        );

    \I__15718\ : LocalMux
    port map (
            O => \N__67141\,
            I => \N__67125\
        );

    \I__15717\ : InMux
    port map (
            O => \N__67140\,
            I => \N__67122\
        );

    \I__15716\ : InMux
    port map (
            O => \N__67137\,
            I => \N__67118\
        );

    \I__15715\ : LocalMux
    port map (
            O => \N__67128\,
            I => \N__67115\
        );

    \I__15714\ : Span4Mux_v
    port map (
            O => \N__67125\,
            I => \N__67112\
        );

    \I__15713\ : LocalMux
    port map (
            O => \N__67122\,
            I => \N__67109\
        );

    \I__15712\ : InMux
    port map (
            O => \N__67121\,
            I => \N__67106\
        );

    \I__15711\ : LocalMux
    port map (
            O => \N__67118\,
            I => \N__67099\
        );

    \I__15710\ : Span4Mux_v
    port map (
            O => \N__67115\,
            I => \N__67099\
        );

    \I__15709\ : Span4Mux_h
    port map (
            O => \N__67112\,
            I => \N__67099\
        );

    \I__15708\ : Span4Mux_v
    port map (
            O => \N__67109\,
            I => \N__67096\
        );

    \I__15707\ : LocalMux
    port map (
            O => \N__67106\,
            I => \c0.data_in_frame_24_6\
        );

    \I__15706\ : Odrv4
    port map (
            O => \N__67099\,
            I => \c0.data_in_frame_24_6\
        );

    \I__15705\ : Odrv4
    port map (
            O => \N__67096\,
            I => \c0.data_in_frame_24_6\
        );

    \I__15704\ : InMux
    port map (
            O => \N__67089\,
            I => \N__67086\
        );

    \I__15703\ : LocalMux
    port map (
            O => \N__67086\,
            I => \N__67083\
        );

    \I__15702\ : Span4Mux_h
    port map (
            O => \N__67083\,
            I => \N__67079\
        );

    \I__15701\ : InMux
    port map (
            O => \N__67082\,
            I => \N__67076\
        );

    \I__15700\ : Odrv4
    port map (
            O => \N__67079\,
            I => \c0.n22495\
        );

    \I__15699\ : LocalMux
    port map (
            O => \N__67076\,
            I => \c0.n22495\
        );

    \I__15698\ : CascadeMux
    port map (
            O => \N__67071\,
            I => \N__67067\
        );

    \I__15697\ : InMux
    port map (
            O => \N__67070\,
            I => \N__67064\
        );

    \I__15696\ : InMux
    port map (
            O => \N__67067\,
            I => \N__67061\
        );

    \I__15695\ : LocalMux
    port map (
            O => \N__67064\,
            I => \c0.data_in_frame_20_1\
        );

    \I__15694\ : LocalMux
    port map (
            O => \N__67061\,
            I => \c0.data_in_frame_20_1\
        );

    \I__15693\ : InMux
    port map (
            O => \N__67056\,
            I => \N__67052\
        );

    \I__15692\ : InMux
    port map (
            O => \N__67055\,
            I => \N__67049\
        );

    \I__15691\ : LocalMux
    port map (
            O => \N__67052\,
            I => \N__67046\
        );

    \I__15690\ : LocalMux
    port map (
            O => \N__67049\,
            I => \N__67043\
        );

    \I__15689\ : Odrv4
    port map (
            O => \N__67046\,
            I => \c0.n58_adj_4355\
        );

    \I__15688\ : Odrv4
    port map (
            O => \N__67043\,
            I => \c0.n58_adj_4355\
        );

    \I__15687\ : InMux
    port map (
            O => \N__67038\,
            I => \N__67034\
        );

    \I__15686\ : InMux
    port map (
            O => \N__67037\,
            I => \N__67030\
        );

    \I__15685\ : LocalMux
    port map (
            O => \N__67034\,
            I => \N__67027\
        );

    \I__15684\ : InMux
    port map (
            O => \N__67033\,
            I => \N__67024\
        );

    \I__15683\ : LocalMux
    port map (
            O => \N__67030\,
            I => \N__67021\
        );

    \I__15682\ : Span4Mux_h
    port map (
            O => \N__67027\,
            I => \N__67018\
        );

    \I__15681\ : LocalMux
    port map (
            O => \N__67024\,
            I => \N__67015\
        );

    \I__15680\ : Span4Mux_v
    port map (
            O => \N__67021\,
            I => \N__67012\
        );

    \I__15679\ : Odrv4
    port map (
            O => \N__67018\,
            I => \c0.n59_adj_4351\
        );

    \I__15678\ : Odrv12
    port map (
            O => \N__67015\,
            I => \c0.n59_adj_4351\
        );

    \I__15677\ : Odrv4
    port map (
            O => \N__67012\,
            I => \c0.n59_adj_4351\
        );

    \I__15676\ : InMux
    port map (
            O => \N__67005\,
            I => \N__67002\
        );

    \I__15675\ : LocalMux
    port map (
            O => \N__67002\,
            I => \N__66999\
        );

    \I__15674\ : Span4Mux_v
    port map (
            O => \N__66999\,
            I => \N__66995\
        );

    \I__15673\ : InMux
    port map (
            O => \N__66998\,
            I => \N__66992\
        );

    \I__15672\ : Odrv4
    port map (
            O => \N__66995\,
            I => \c0.n28_adj_4363\
        );

    \I__15671\ : LocalMux
    port map (
            O => \N__66992\,
            I => \c0.n28_adj_4363\
        );

    \I__15670\ : InMux
    port map (
            O => \N__66987\,
            I => \N__66979\
        );

    \I__15669\ : InMux
    port map (
            O => \N__66986\,
            I => \N__66979\
        );

    \I__15668\ : InMux
    port map (
            O => \N__66985\,
            I => \N__66976\
        );

    \I__15667\ : InMux
    port map (
            O => \N__66984\,
            I => \N__66973\
        );

    \I__15666\ : LocalMux
    port map (
            O => \N__66979\,
            I => \N__66970\
        );

    \I__15665\ : LocalMux
    port map (
            O => \N__66976\,
            I => \N__66965\
        );

    \I__15664\ : LocalMux
    port map (
            O => \N__66973\,
            I => \N__66965\
        );

    \I__15663\ : Span4Mux_v
    port map (
            O => \N__66970\,
            I => \N__66962\
        );

    \I__15662\ : Odrv4
    port map (
            O => \N__66965\,
            I => \c0.n23691\
        );

    \I__15661\ : Odrv4
    port map (
            O => \N__66962\,
            I => \c0.n23691\
        );

    \I__15660\ : CascadeMux
    port map (
            O => \N__66957\,
            I => \N__66954\
        );

    \I__15659\ : InMux
    port map (
            O => \N__66954\,
            I => \N__66951\
        );

    \I__15658\ : LocalMux
    port map (
            O => \N__66951\,
            I => \N__66947\
        );

    \I__15657\ : InMux
    port map (
            O => \N__66950\,
            I => \N__66944\
        );

    \I__15656\ : Span4Mux_h
    port map (
            O => \N__66947\,
            I => \N__66939\
        );

    \I__15655\ : LocalMux
    port map (
            O => \N__66944\,
            I => \N__66939\
        );

    \I__15654\ : Span4Mux_h
    port map (
            O => \N__66939\,
            I => \N__66936\
        );

    \I__15653\ : Span4Mux_h
    port map (
            O => \N__66936\,
            I => \N__66933\
        );

    \I__15652\ : Odrv4
    port map (
            O => \N__66933\,
            I => \c0.n22577\
        );

    \I__15651\ : InMux
    port map (
            O => \N__66930\,
            I => \N__66926\
        );

    \I__15650\ : InMux
    port map (
            O => \N__66929\,
            I => \N__66923\
        );

    \I__15649\ : LocalMux
    port map (
            O => \N__66926\,
            I => \N__66920\
        );

    \I__15648\ : LocalMux
    port map (
            O => \N__66923\,
            I => \N__66916\
        );

    \I__15647\ : Span4Mux_h
    port map (
            O => \N__66920\,
            I => \N__66913\
        );

    \I__15646\ : InMux
    port map (
            O => \N__66919\,
            I => \N__66910\
        );

    \I__15645\ : Odrv12
    port map (
            O => \N__66916\,
            I => \c0.n21414\
        );

    \I__15644\ : Odrv4
    port map (
            O => \N__66913\,
            I => \c0.n21414\
        );

    \I__15643\ : LocalMux
    port map (
            O => \N__66910\,
            I => \c0.n21414\
        );

    \I__15642\ : CascadeMux
    port map (
            O => \N__66903\,
            I => \c0.n10_adj_4524_cascade_\
        );

    \I__15641\ : CascadeMux
    port map (
            O => \N__66900\,
            I => \N__66894\
        );

    \I__15640\ : InMux
    port map (
            O => \N__66899\,
            I => \N__66890\
        );

    \I__15639\ : InMux
    port map (
            O => \N__66898\,
            I => \N__66887\
        );

    \I__15638\ : InMux
    port map (
            O => \N__66897\,
            I => \N__66884\
        );

    \I__15637\ : InMux
    port map (
            O => \N__66894\,
            I => \N__66881\
        );

    \I__15636\ : InMux
    port map (
            O => \N__66893\,
            I => \N__66878\
        );

    \I__15635\ : LocalMux
    port map (
            O => \N__66890\,
            I => \N__66875\
        );

    \I__15634\ : LocalMux
    port map (
            O => \N__66887\,
            I => \N__66872\
        );

    \I__15633\ : LocalMux
    port map (
            O => \N__66884\,
            I => \N__66864\
        );

    \I__15632\ : LocalMux
    port map (
            O => \N__66881\,
            I => \N__66864\
        );

    \I__15631\ : LocalMux
    port map (
            O => \N__66878\,
            I => \N__66864\
        );

    \I__15630\ : Span4Mux_v
    port map (
            O => \N__66875\,
            I => \N__66858\
        );

    \I__15629\ : Span4Mux_h
    port map (
            O => \N__66872\,
            I => \N__66858\
        );

    \I__15628\ : InMux
    port map (
            O => \N__66871\,
            I => \N__66855\
        );

    \I__15627\ : Span4Mux_v
    port map (
            O => \N__66864\,
            I => \N__66852\
        );

    \I__15626\ : InMux
    port map (
            O => \N__66863\,
            I => \N__66849\
        );

    \I__15625\ : Span4Mux_v
    port map (
            O => \N__66858\,
            I => \N__66846\
        );

    \I__15624\ : LocalMux
    port map (
            O => \N__66855\,
            I => \N__66841\
        );

    \I__15623\ : Span4Mux_h
    port map (
            O => \N__66852\,
            I => \N__66841\
        );

    \I__15622\ : LocalMux
    port map (
            O => \N__66849\,
            I => \N__66838\
        );

    \I__15621\ : Odrv4
    port map (
            O => \N__66846\,
            I => \c0.n13797\
        );

    \I__15620\ : Odrv4
    port map (
            O => \N__66841\,
            I => \c0.n13797\
        );

    \I__15619\ : Odrv4
    port map (
            O => \N__66838\,
            I => \c0.n13797\
        );

    \I__15618\ : InMux
    port map (
            O => \N__66831\,
            I => \N__66828\
        );

    \I__15617\ : LocalMux
    port map (
            O => \N__66828\,
            I => \N__66824\
        );

    \I__15616\ : InMux
    port map (
            O => \N__66827\,
            I => \N__66821\
        );

    \I__15615\ : Span4Mux_v
    port map (
            O => \N__66824\,
            I => \N__66818\
        );

    \I__15614\ : LocalMux
    port map (
            O => \N__66821\,
            I => \c0.n24576\
        );

    \I__15613\ : Odrv4
    port map (
            O => \N__66818\,
            I => \c0.n24576\
        );

    \I__15612\ : InMux
    port map (
            O => \N__66813\,
            I => \N__66808\
        );

    \I__15611\ : InMux
    port map (
            O => \N__66812\,
            I => \N__66802\
        );

    \I__15610\ : InMux
    port map (
            O => \N__66811\,
            I => \N__66802\
        );

    \I__15609\ : LocalMux
    port map (
            O => \N__66808\,
            I => \N__66799\
        );

    \I__15608\ : CascadeMux
    port map (
            O => \N__66807\,
            I => \N__66796\
        );

    \I__15607\ : LocalMux
    port map (
            O => \N__66802\,
            I => \N__66793\
        );

    \I__15606\ : Span4Mux_h
    port map (
            O => \N__66799\,
            I => \N__66790\
        );

    \I__15605\ : InMux
    port map (
            O => \N__66796\,
            I => \N__66787\
        );

    \I__15604\ : Span4Mux_h
    port map (
            O => \N__66793\,
            I => \N__66784\
        );

    \I__15603\ : Span4Mux_h
    port map (
            O => \N__66790\,
            I => \N__66781\
        );

    \I__15602\ : LocalMux
    port map (
            O => \N__66787\,
            I => \N__66776\
        );

    \I__15601\ : Span4Mux_h
    port map (
            O => \N__66784\,
            I => \N__66776\
        );

    \I__15600\ : Odrv4
    port map (
            O => \N__66781\,
            I => \c0.data_in_frame_26_2\
        );

    \I__15599\ : Odrv4
    port map (
            O => \N__66776\,
            I => \c0.data_in_frame_26_2\
        );

    \I__15598\ : CascadeMux
    port map (
            O => \N__66771\,
            I => \c0.n24576_cascade_\
        );

    \I__15597\ : InMux
    port map (
            O => \N__66768\,
            I => \N__66765\
        );

    \I__15596\ : LocalMux
    port map (
            O => \N__66765\,
            I => \N__66762\
        );

    \I__15595\ : Span4Mux_v
    port map (
            O => \N__66762\,
            I => \N__66759\
        );

    \I__15594\ : Odrv4
    port map (
            O => \N__66759\,
            I => \c0.n14_adj_4519\
        );

    \I__15593\ : InMux
    port map (
            O => \N__66756\,
            I => \N__66753\
        );

    \I__15592\ : LocalMux
    port map (
            O => \N__66753\,
            I => \N__66747\
        );

    \I__15591\ : InMux
    port map (
            O => \N__66752\,
            I => \N__66743\
        );

    \I__15590\ : InMux
    port map (
            O => \N__66751\,
            I => \N__66740\
        );

    \I__15589\ : InMux
    port map (
            O => \N__66750\,
            I => \N__66737\
        );

    \I__15588\ : Span4Mux_h
    port map (
            O => \N__66747\,
            I => \N__66734\
        );

    \I__15587\ : InMux
    port map (
            O => \N__66746\,
            I => \N__66731\
        );

    \I__15586\ : LocalMux
    port map (
            O => \N__66743\,
            I => \N__66724\
        );

    \I__15585\ : LocalMux
    port map (
            O => \N__66740\,
            I => \N__66724\
        );

    \I__15584\ : LocalMux
    port map (
            O => \N__66737\,
            I => \N__66724\
        );

    \I__15583\ : Span4Mux_h
    port map (
            O => \N__66734\,
            I => \N__66721\
        );

    \I__15582\ : LocalMux
    port map (
            O => \N__66731\,
            I => data_in_frame_21_4
        );

    \I__15581\ : Odrv12
    port map (
            O => \N__66724\,
            I => data_in_frame_21_4
        );

    \I__15580\ : Odrv4
    port map (
            O => \N__66721\,
            I => data_in_frame_21_4
        );

    \I__15579\ : InMux
    port map (
            O => \N__66714\,
            I => \N__66711\
        );

    \I__15578\ : LocalMux
    port map (
            O => \N__66711\,
            I => \N__66706\
        );

    \I__15577\ : InMux
    port map (
            O => \N__66710\,
            I => \N__66703\
        );

    \I__15576\ : InMux
    port map (
            O => \N__66709\,
            I => \N__66700\
        );

    \I__15575\ : Span4Mux_h
    port map (
            O => \N__66706\,
            I => \N__66697\
        );

    \I__15574\ : LocalMux
    port map (
            O => \N__66703\,
            I => \N__66694\
        );

    \I__15573\ : LocalMux
    port map (
            O => \N__66700\,
            I => \c0.n23733\
        );

    \I__15572\ : Odrv4
    port map (
            O => \N__66697\,
            I => \c0.n23733\
        );

    \I__15571\ : Odrv4
    port map (
            O => \N__66694\,
            I => \c0.n23733\
        );

    \I__15570\ : InMux
    port map (
            O => \N__66687\,
            I => \N__66684\
        );

    \I__15569\ : LocalMux
    port map (
            O => \N__66684\,
            I => \c0.n22686\
        );

    \I__15568\ : InMux
    port map (
            O => \N__66681\,
            I => \N__66678\
        );

    \I__15567\ : LocalMux
    port map (
            O => \N__66678\,
            I => \N__66675\
        );

    \I__15566\ : Span4Mux_v
    port map (
            O => \N__66675\,
            I => \N__66672\
        );

    \I__15565\ : Odrv4
    port map (
            O => \N__66672\,
            I => \c0.n5_adj_4472\
        );

    \I__15564\ : CascadeMux
    port map (
            O => \N__66669\,
            I => \c0.n22686_cascade_\
        );

    \I__15563\ : InMux
    port map (
            O => \N__66666\,
            I => \N__66663\
        );

    \I__15562\ : LocalMux
    port map (
            O => \N__66663\,
            I => \N__66658\
        );

    \I__15561\ : InMux
    port map (
            O => \N__66662\,
            I => \N__66655\
        );

    \I__15560\ : InMux
    port map (
            O => \N__66661\,
            I => \N__66651\
        );

    \I__15559\ : Span4Mux_v
    port map (
            O => \N__66658\,
            I => \N__66647\
        );

    \I__15558\ : LocalMux
    port map (
            O => \N__66655\,
            I => \N__66644\
        );

    \I__15557\ : InMux
    port map (
            O => \N__66654\,
            I => \N__66641\
        );

    \I__15556\ : LocalMux
    port map (
            O => \N__66651\,
            I => \N__66638\
        );

    \I__15555\ : InMux
    port map (
            O => \N__66650\,
            I => \N__66634\
        );

    \I__15554\ : Span4Mux_h
    port map (
            O => \N__66647\,
            I => \N__66629\
        );

    \I__15553\ : Span4Mux_v
    port map (
            O => \N__66644\,
            I => \N__66629\
        );

    \I__15552\ : LocalMux
    port map (
            O => \N__66641\,
            I => \N__66624\
        );

    \I__15551\ : Span4Mux_h
    port map (
            O => \N__66638\,
            I => \N__66624\
        );

    \I__15550\ : InMux
    port map (
            O => \N__66637\,
            I => \N__66621\
        );

    \I__15549\ : LocalMux
    port map (
            O => \N__66634\,
            I => \c0.data_in_frame_18_3\
        );

    \I__15548\ : Odrv4
    port map (
            O => \N__66629\,
            I => \c0.data_in_frame_18_3\
        );

    \I__15547\ : Odrv4
    port map (
            O => \N__66624\,
            I => \c0.data_in_frame_18_3\
        );

    \I__15546\ : LocalMux
    port map (
            O => \N__66621\,
            I => \c0.data_in_frame_18_3\
        );

    \I__15545\ : InMux
    port map (
            O => \N__66612\,
            I => \N__66609\
        );

    \I__15544\ : LocalMux
    port map (
            O => \N__66609\,
            I => \N__66605\
        );

    \I__15543\ : InMux
    port map (
            O => \N__66608\,
            I => \N__66602\
        );

    \I__15542\ : Odrv4
    port map (
            O => \N__66605\,
            I => \c0.n5_adj_4335\
        );

    \I__15541\ : LocalMux
    port map (
            O => \N__66602\,
            I => \c0.n5_adj_4335\
        );

    \I__15540\ : InMux
    port map (
            O => \N__66597\,
            I => \N__66594\
        );

    \I__15539\ : LocalMux
    port map (
            O => \N__66594\,
            I => \N__66590\
        );

    \I__15538\ : InMux
    port map (
            O => \N__66593\,
            I => \N__66587\
        );

    \I__15537\ : Span4Mux_h
    port map (
            O => \N__66590\,
            I => \N__66584\
        );

    \I__15536\ : LocalMux
    port map (
            O => \N__66587\,
            I => \c0.n4_adj_4568\
        );

    \I__15535\ : Odrv4
    port map (
            O => \N__66584\,
            I => \c0.n4_adj_4568\
        );

    \I__15534\ : InMux
    port map (
            O => \N__66579\,
            I => \N__66576\
        );

    \I__15533\ : LocalMux
    port map (
            O => \N__66576\,
            I => \N__66573\
        );

    \I__15532\ : Odrv12
    port map (
            O => \N__66573\,
            I => \c0.n15_adj_4569\
        );

    \I__15531\ : InMux
    port map (
            O => \N__66570\,
            I => \N__66566\
        );

    \I__15530\ : InMux
    port map (
            O => \N__66569\,
            I => \N__66562\
        );

    \I__15529\ : LocalMux
    port map (
            O => \N__66566\,
            I => \N__66559\
        );

    \I__15528\ : InMux
    port map (
            O => \N__66565\,
            I => \N__66556\
        );

    \I__15527\ : LocalMux
    port map (
            O => \N__66562\,
            I => \N__66553\
        );

    \I__15526\ : Span4Mux_h
    port map (
            O => \N__66559\,
            I => \N__66549\
        );

    \I__15525\ : LocalMux
    port map (
            O => \N__66556\,
            I => \N__66546\
        );

    \I__15524\ : Span4Mux_v
    port map (
            O => \N__66553\,
            I => \N__66543\
        );

    \I__15523\ : InMux
    port map (
            O => \N__66552\,
            I => \N__66540\
        );

    \I__15522\ : Span4Mux_h
    port map (
            O => \N__66549\,
            I => \N__66537\
        );

    \I__15521\ : Span4Mux_v
    port map (
            O => \N__66546\,
            I => \N__66532\
        );

    \I__15520\ : Span4Mux_h
    port map (
            O => \N__66543\,
            I => \N__66532\
        );

    \I__15519\ : LocalMux
    port map (
            O => \N__66540\,
            I => \c0.data_in_frame_18_7\
        );

    \I__15518\ : Odrv4
    port map (
            O => \N__66537\,
            I => \c0.data_in_frame_18_7\
        );

    \I__15517\ : Odrv4
    port map (
            O => \N__66532\,
            I => \c0.data_in_frame_18_7\
        );

    \I__15516\ : InMux
    port map (
            O => \N__66525\,
            I => \N__66522\
        );

    \I__15515\ : LocalMux
    port map (
            O => \N__66522\,
            I => \N__66518\
        );

    \I__15514\ : CascadeMux
    port map (
            O => \N__66521\,
            I => \N__66514\
        );

    \I__15513\ : Span12Mux_v
    port map (
            O => \N__66518\,
            I => \N__66511\
        );

    \I__15512\ : InMux
    port map (
            O => \N__66517\,
            I => \N__66506\
        );

    \I__15511\ : InMux
    port map (
            O => \N__66514\,
            I => \N__66506\
        );

    \I__15510\ : Odrv12
    port map (
            O => \N__66511\,
            I => data_in_frame_22_5
        );

    \I__15509\ : LocalMux
    port map (
            O => \N__66506\,
            I => data_in_frame_22_5
        );

    \I__15508\ : CascadeMux
    port map (
            O => \N__66501\,
            I => \N__66497\
        );

    \I__15507\ : CascadeMux
    port map (
            O => \N__66500\,
            I => \N__66492\
        );

    \I__15506\ : InMux
    port map (
            O => \N__66497\,
            I => \N__66487\
        );

    \I__15505\ : InMux
    port map (
            O => \N__66496\,
            I => \N__66487\
        );

    \I__15504\ : InMux
    port map (
            O => \N__66495\,
            I => \N__66484\
        );

    \I__15503\ : InMux
    port map (
            O => \N__66492\,
            I => \N__66481\
        );

    \I__15502\ : LocalMux
    port map (
            O => \N__66487\,
            I => \N__66478\
        );

    \I__15501\ : LocalMux
    port map (
            O => \N__66484\,
            I => \N__66475\
        );

    \I__15500\ : LocalMux
    port map (
            O => \N__66481\,
            I => \N__66470\
        );

    \I__15499\ : Span4Mux_h
    port map (
            O => \N__66478\,
            I => \N__66470\
        );

    \I__15498\ : Odrv4
    port map (
            O => \N__66475\,
            I => \c0.data_in_frame_17_5\
        );

    \I__15497\ : Odrv4
    port map (
            O => \N__66470\,
            I => \c0.data_in_frame_17_5\
        );

    \I__15496\ : InMux
    port map (
            O => \N__66465\,
            I => \N__66461\
        );

    \I__15495\ : InMux
    port map (
            O => \N__66464\,
            I => \N__66458\
        );

    \I__15494\ : LocalMux
    port map (
            O => \N__66461\,
            I => \N__66455\
        );

    \I__15493\ : LocalMux
    port map (
            O => \N__66458\,
            I => \N__66452\
        );

    \I__15492\ : Span4Mux_v
    port map (
            O => \N__66455\,
            I => \N__66447\
        );

    \I__15491\ : Span4Mux_h
    port map (
            O => \N__66452\,
            I => \N__66447\
        );

    \I__15490\ : Odrv4
    port map (
            O => \N__66447\,
            I => \c0.n22748\
        );

    \I__15489\ : CascadeMux
    port map (
            O => \N__66444\,
            I => \c0.n14_adj_4623_cascade_\
        );

    \I__15488\ : InMux
    port map (
            O => \N__66441\,
            I => \N__66438\
        );

    \I__15487\ : LocalMux
    port map (
            O => \N__66438\,
            I => \c0.n15_adj_4624\
        );

    \I__15486\ : InMux
    port map (
            O => \N__66435\,
            I => \N__66432\
        );

    \I__15485\ : LocalMux
    port map (
            O => \N__66432\,
            I => \N__66427\
        );

    \I__15484\ : InMux
    port map (
            O => \N__66431\,
            I => \N__66422\
        );

    \I__15483\ : InMux
    port map (
            O => \N__66430\,
            I => \N__66419\
        );

    \I__15482\ : Span4Mux_h
    port map (
            O => \N__66427\,
            I => \N__66416\
        );

    \I__15481\ : InMux
    port map (
            O => \N__66426\,
            I => \N__66411\
        );

    \I__15480\ : InMux
    port map (
            O => \N__66425\,
            I => \N__66411\
        );

    \I__15479\ : LocalMux
    port map (
            O => \N__66422\,
            I => \N__66408\
        );

    \I__15478\ : LocalMux
    port map (
            O => \N__66419\,
            I => \N__66403\
        );

    \I__15477\ : Span4Mux_h
    port map (
            O => \N__66416\,
            I => \N__66403\
        );

    \I__15476\ : LocalMux
    port map (
            O => \N__66411\,
            I => data_in_frame_21_1
        );

    \I__15475\ : Odrv4
    port map (
            O => \N__66408\,
            I => data_in_frame_21_1
        );

    \I__15474\ : Odrv4
    port map (
            O => \N__66403\,
            I => data_in_frame_21_1
        );

    \I__15473\ : CascadeMux
    port map (
            O => \N__66396\,
            I => \c0.n13963_cascade_\
        );

    \I__15472\ : InMux
    port map (
            O => \N__66393\,
            I => \N__66389\
        );

    \I__15471\ : InMux
    port map (
            O => \N__66392\,
            I => \N__66386\
        );

    \I__15470\ : LocalMux
    port map (
            O => \N__66389\,
            I => \N__66381\
        );

    \I__15469\ : LocalMux
    port map (
            O => \N__66386\,
            I => \N__66381\
        );

    \I__15468\ : Span4Mux_v
    port map (
            O => \N__66381\,
            I => \N__66378\
        );

    \I__15467\ : Odrv4
    port map (
            O => \N__66378\,
            I => \c0.n22508\
        );

    \I__15466\ : InMux
    port map (
            O => \N__66375\,
            I => \N__66372\
        );

    \I__15465\ : LocalMux
    port map (
            O => \N__66372\,
            I => \c0.n40_adj_4342\
        );

    \I__15464\ : InMux
    port map (
            O => \N__66369\,
            I => \N__66366\
        );

    \I__15463\ : LocalMux
    port map (
            O => \N__66366\,
            I => \N__66361\
        );

    \I__15462\ : InMux
    port map (
            O => \N__66365\,
            I => \N__66356\
        );

    \I__15461\ : InMux
    port map (
            O => \N__66364\,
            I => \N__66356\
        );

    \I__15460\ : Span12Mux_h
    port map (
            O => \N__66361\,
            I => \N__66352\
        );

    \I__15459\ : LocalMux
    port map (
            O => \N__66356\,
            I => \N__66349\
        );

    \I__15458\ : InMux
    port map (
            O => \N__66355\,
            I => \N__66346\
        );

    \I__15457\ : Odrv12
    port map (
            O => \N__66352\,
            I => \c0.n13604\
        );

    \I__15456\ : Odrv4
    port map (
            O => \N__66349\,
            I => \c0.n13604\
        );

    \I__15455\ : LocalMux
    port map (
            O => \N__66346\,
            I => \c0.n13604\
        );

    \I__15454\ : CascadeMux
    port map (
            O => \N__66339\,
            I => \c0.n7_adj_4251_cascade_\
        );

    \I__15453\ : InMux
    port map (
            O => \N__66336\,
            I => \N__66330\
        );

    \I__15452\ : InMux
    port map (
            O => \N__66335\,
            I => \N__66327\
        );

    \I__15451\ : InMux
    port map (
            O => \N__66334\,
            I => \N__66322\
        );

    \I__15450\ : InMux
    port map (
            O => \N__66333\,
            I => \N__66322\
        );

    \I__15449\ : LocalMux
    port map (
            O => \N__66330\,
            I => \c0.n23224\
        );

    \I__15448\ : LocalMux
    port map (
            O => \N__66327\,
            I => \c0.n23224\
        );

    \I__15447\ : LocalMux
    port map (
            O => \N__66322\,
            I => \c0.n23224\
        );

    \I__15446\ : InMux
    port map (
            O => \N__66315\,
            I => \N__66312\
        );

    \I__15445\ : LocalMux
    port map (
            O => \N__66312\,
            I => \c0.n7_adj_4251\
        );

    \I__15444\ : InMux
    port map (
            O => \N__66309\,
            I => \N__66306\
        );

    \I__15443\ : LocalMux
    port map (
            O => \N__66306\,
            I => \N__66303\
        );

    \I__15442\ : Span4Mux_h
    port map (
            O => \N__66303\,
            I => \N__66299\
        );

    \I__15441\ : InMux
    port map (
            O => \N__66302\,
            I => \N__66296\
        );

    \I__15440\ : Span4Mux_h
    port map (
            O => \N__66299\,
            I => \N__66293\
        );

    \I__15439\ : LocalMux
    port map (
            O => \N__66296\,
            I => data_in_frame_22_7
        );

    \I__15438\ : Odrv4
    port map (
            O => \N__66293\,
            I => data_in_frame_22_7
        );

    \I__15437\ : InMux
    port map (
            O => \N__66288\,
            I => \N__66285\
        );

    \I__15436\ : LocalMux
    port map (
            O => \N__66285\,
            I => \N__66282\
        );

    \I__15435\ : Span4Mux_v
    port map (
            O => \N__66282\,
            I => \N__66279\
        );

    \I__15434\ : Sp12to4
    port map (
            O => \N__66279\,
            I => \N__66276\
        );

    \I__15433\ : Odrv12
    port map (
            O => \N__66276\,
            I => \c0.n22825\
        );

    \I__15432\ : CascadeMux
    port map (
            O => \N__66273\,
            I => \N__66268\
        );

    \I__15431\ : InMux
    port map (
            O => \N__66272\,
            I => \N__66265\
        );

    \I__15430\ : InMux
    port map (
            O => \N__66271\,
            I => \N__66262\
        );

    \I__15429\ : InMux
    port map (
            O => \N__66268\,
            I => \N__66259\
        );

    \I__15428\ : LocalMux
    port map (
            O => \N__66265\,
            I => \N__66256\
        );

    \I__15427\ : LocalMux
    port map (
            O => \N__66262\,
            I => \N__66253\
        );

    \I__15426\ : LocalMux
    port map (
            O => \N__66259\,
            I => \c0.data_in_frame_15_4\
        );

    \I__15425\ : Odrv12
    port map (
            O => \N__66256\,
            I => \c0.data_in_frame_15_4\
        );

    \I__15424\ : Odrv4
    port map (
            O => \N__66253\,
            I => \c0.data_in_frame_15_4\
        );

    \I__15423\ : InMux
    port map (
            O => \N__66246\,
            I => \N__66243\
        );

    \I__15422\ : LocalMux
    port map (
            O => \N__66243\,
            I => \N__66239\
        );

    \I__15421\ : InMux
    port map (
            O => \N__66242\,
            I => \N__66236\
        );

    \I__15420\ : Span4Mux_v
    port map (
            O => \N__66239\,
            I => \N__66233\
        );

    \I__15419\ : LocalMux
    port map (
            O => \N__66236\,
            I => \c0.data_in_frame_18_2\
        );

    \I__15418\ : Odrv4
    port map (
            O => \N__66233\,
            I => \c0.data_in_frame_18_2\
        );

    \I__15417\ : InMux
    port map (
            O => \N__66228\,
            I => \N__66224\
        );

    \I__15416\ : InMux
    port map (
            O => \N__66227\,
            I => \N__66221\
        );

    \I__15415\ : LocalMux
    port map (
            O => \N__66224\,
            I => \N__66217\
        );

    \I__15414\ : LocalMux
    port map (
            O => \N__66221\,
            I => \N__66214\
        );

    \I__15413\ : CascadeMux
    port map (
            O => \N__66220\,
            I => \N__66211\
        );

    \I__15412\ : Span4Mux_v
    port map (
            O => \N__66217\,
            I => \N__66208\
        );

    \I__15411\ : Span4Mux_v
    port map (
            O => \N__66214\,
            I => \N__66205\
        );

    \I__15410\ : InMux
    port map (
            O => \N__66211\,
            I => \N__66202\
        );

    \I__15409\ : Span4Mux_h
    port map (
            O => \N__66208\,
            I => \N__66199\
        );

    \I__15408\ : Span4Mux_v
    port map (
            O => \N__66205\,
            I => \N__66196\
        );

    \I__15407\ : LocalMux
    port map (
            O => \N__66202\,
            I => \c0.data_in_frame_18_4\
        );

    \I__15406\ : Odrv4
    port map (
            O => \N__66199\,
            I => \c0.data_in_frame_18_4\
        );

    \I__15405\ : Odrv4
    port map (
            O => \N__66196\,
            I => \c0.data_in_frame_18_4\
        );

    \I__15404\ : InMux
    port map (
            O => \N__66189\,
            I => \N__66186\
        );

    \I__15403\ : LocalMux
    port map (
            O => \N__66186\,
            I => \c0.n12_adj_4455\
        );

    \I__15402\ : CascadeMux
    port map (
            O => \N__66183\,
            I => \N__66180\
        );

    \I__15401\ : InMux
    port map (
            O => \N__66180\,
            I => \N__66177\
        );

    \I__15400\ : LocalMux
    port map (
            O => \N__66177\,
            I => \N__66174\
        );

    \I__15399\ : Span12Mux_h
    port map (
            O => \N__66174\,
            I => \N__66170\
        );

    \I__15398\ : InMux
    port map (
            O => \N__66173\,
            I => \N__66167\
        );

    \I__15397\ : Odrv12
    port map (
            O => \N__66170\,
            I => \c0.n22463\
        );

    \I__15396\ : LocalMux
    port map (
            O => \N__66167\,
            I => \c0.n22463\
        );

    \I__15395\ : InMux
    port map (
            O => \N__66162\,
            I => \N__66157\
        );

    \I__15394\ : InMux
    port map (
            O => \N__66161\,
            I => \N__66154\
        );

    \I__15393\ : InMux
    port map (
            O => \N__66160\,
            I => \N__66151\
        );

    \I__15392\ : LocalMux
    port map (
            O => \N__66157\,
            I => \N__66146\
        );

    \I__15391\ : LocalMux
    port map (
            O => \N__66154\,
            I => \N__66146\
        );

    \I__15390\ : LocalMux
    port map (
            O => \N__66151\,
            I => \N__66143\
        );

    \I__15389\ : Span4Mux_v
    port map (
            O => \N__66146\,
            I => \N__66138\
        );

    \I__15388\ : Span4Mux_v
    port map (
            O => \N__66143\,
            I => \N__66138\
        );

    \I__15387\ : Odrv4
    port map (
            O => \N__66138\,
            I => \c0.n24540\
        );

    \I__15386\ : InMux
    port map (
            O => \N__66135\,
            I => \N__66130\
        );

    \I__15385\ : InMux
    port map (
            O => \N__66134\,
            I => \N__66125\
        );

    \I__15384\ : InMux
    port map (
            O => \N__66133\,
            I => \N__66125\
        );

    \I__15383\ : LocalMux
    port map (
            O => \N__66130\,
            I => \N__66122\
        );

    \I__15382\ : LocalMux
    port map (
            O => \N__66125\,
            I => \c0.n23507\
        );

    \I__15381\ : Odrv4
    port map (
            O => \N__66122\,
            I => \c0.n23507\
        );

    \I__15380\ : CascadeMux
    port map (
            O => \N__66117\,
            I => \N__66113\
        );

    \I__15379\ : InMux
    port map (
            O => \N__66116\,
            I => \N__66110\
        );

    \I__15378\ : InMux
    port map (
            O => \N__66113\,
            I => \N__66107\
        );

    \I__15377\ : LocalMux
    port map (
            O => \N__66110\,
            I => \N__66102\
        );

    \I__15376\ : LocalMux
    port map (
            O => \N__66107\,
            I => \N__66102\
        );

    \I__15375\ : Odrv4
    port map (
            O => \N__66102\,
            I => data_in_frame_21_0
        );

    \I__15374\ : InMux
    port map (
            O => \N__66099\,
            I => \N__66093\
        );

    \I__15373\ : CascadeMux
    port map (
            O => \N__66098\,
            I => \N__66090\
        );

    \I__15372\ : InMux
    port map (
            O => \N__66097\,
            I => \N__66087\
        );

    \I__15371\ : InMux
    port map (
            O => \N__66096\,
            I => \N__66084\
        );

    \I__15370\ : LocalMux
    port map (
            O => \N__66093\,
            I => \N__66081\
        );

    \I__15369\ : InMux
    port map (
            O => \N__66090\,
            I => \N__66078\
        );

    \I__15368\ : LocalMux
    port map (
            O => \N__66087\,
            I => \N__66073\
        );

    \I__15367\ : LocalMux
    port map (
            O => \N__66084\,
            I => \N__66073\
        );

    \I__15366\ : Span4Mux_h
    port map (
            O => \N__66081\,
            I => \N__66070\
        );

    \I__15365\ : LocalMux
    port map (
            O => \N__66078\,
            I => \N__66063\
        );

    \I__15364\ : Span4Mux_v
    port map (
            O => \N__66073\,
            I => \N__66063\
        );

    \I__15363\ : Span4Mux_h
    port map (
            O => \N__66070\,
            I => \N__66063\
        );

    \I__15362\ : Odrv4
    port map (
            O => \N__66063\,
            I => \c0.data_in_frame_17_0\
        );

    \I__15361\ : InMux
    port map (
            O => \N__66060\,
            I => \N__66057\
        );

    \I__15360\ : LocalMux
    port map (
            O => \N__66057\,
            I => \N__66054\
        );

    \I__15359\ : Span4Mux_h
    port map (
            O => \N__66054\,
            I => \N__66049\
        );

    \I__15358\ : InMux
    port map (
            O => \N__66053\,
            I => \N__66044\
        );

    \I__15357\ : InMux
    port map (
            O => \N__66052\,
            I => \N__66044\
        );

    \I__15356\ : Span4Mux_h
    port map (
            O => \N__66049\,
            I => \N__66041\
        );

    \I__15355\ : LocalMux
    port map (
            O => \N__66044\,
            I => \N__66038\
        );

    \I__15354\ : Odrv4
    port map (
            O => \N__66041\,
            I => \c0.n23313\
        );

    \I__15353\ : Odrv4
    port map (
            O => \N__66038\,
            I => \c0.n23313\
        );

    \I__15352\ : InMux
    port map (
            O => \N__66033\,
            I => \N__66027\
        );

    \I__15351\ : InMux
    port map (
            O => \N__66032\,
            I => \N__66027\
        );

    \I__15350\ : LocalMux
    port map (
            O => \N__66027\,
            I => \N__66024\
        );

    \I__15349\ : Span4Mux_v
    port map (
            O => \N__66024\,
            I => \N__66021\
        );

    \I__15348\ : Odrv4
    port map (
            O => \N__66021\,
            I => \c0.n26_adj_4578\
        );

    \I__15347\ : InMux
    port map (
            O => \N__66018\,
            I => \N__66011\
        );

    \I__15346\ : InMux
    port map (
            O => \N__66017\,
            I => \N__66011\
        );

    \I__15345\ : CascadeMux
    port map (
            O => \N__66016\,
            I => \N__66007\
        );

    \I__15344\ : LocalMux
    port map (
            O => \N__66011\,
            I => \N__66003\
        );

    \I__15343\ : InMux
    port map (
            O => \N__66010\,
            I => \N__66000\
        );

    \I__15342\ : InMux
    port map (
            O => \N__66007\,
            I => \N__65995\
        );

    \I__15341\ : InMux
    port map (
            O => \N__66006\,
            I => \N__65995\
        );

    \I__15340\ : Odrv4
    port map (
            O => \N__66003\,
            I => \c0.data_in_frame_13_5\
        );

    \I__15339\ : LocalMux
    port map (
            O => \N__66000\,
            I => \c0.data_in_frame_13_5\
        );

    \I__15338\ : LocalMux
    port map (
            O => \N__65995\,
            I => \c0.data_in_frame_13_5\
        );

    \I__15337\ : InMux
    port map (
            O => \N__65988\,
            I => \N__65984\
        );

    \I__15336\ : CascadeMux
    port map (
            O => \N__65987\,
            I => \N__65981\
        );

    \I__15335\ : LocalMux
    port map (
            O => \N__65984\,
            I => \N__65977\
        );

    \I__15334\ : InMux
    port map (
            O => \N__65981\,
            I => \N__65972\
        );

    \I__15333\ : InMux
    port map (
            O => \N__65980\,
            I => \N__65972\
        );

    \I__15332\ : Span4Mux_v
    port map (
            O => \N__65977\,
            I => \N__65969\
        );

    \I__15331\ : LocalMux
    port map (
            O => \N__65972\,
            I => \c0.data_in_frame_17_7\
        );

    \I__15330\ : Odrv4
    port map (
            O => \N__65969\,
            I => \c0.data_in_frame_17_7\
        );

    \I__15329\ : InMux
    port map (
            O => \N__65964\,
            I => \N__65961\
        );

    \I__15328\ : LocalMux
    port map (
            O => \N__65961\,
            I => \N__65956\
        );

    \I__15327\ : CascadeMux
    port map (
            O => \N__65960\,
            I => \N__65953\
        );

    \I__15326\ : InMux
    port map (
            O => \N__65959\,
            I => \N__65950\
        );

    \I__15325\ : Span4Mux_h
    port map (
            O => \N__65956\,
            I => \N__65947\
        );

    \I__15324\ : InMux
    port map (
            O => \N__65953\,
            I => \N__65944\
        );

    \I__15323\ : LocalMux
    port map (
            O => \N__65950\,
            I => \N__65941\
        );

    \I__15322\ : Span4Mux_h
    port map (
            O => \N__65947\,
            I => \N__65938\
        );

    \I__15321\ : LocalMux
    port map (
            O => \N__65944\,
            I => \c0.data_in_frame_16_2\
        );

    \I__15320\ : Odrv12
    port map (
            O => \N__65941\,
            I => \c0.data_in_frame_16_2\
        );

    \I__15319\ : Odrv4
    port map (
            O => \N__65938\,
            I => \c0.data_in_frame_16_2\
        );

    \I__15318\ : InMux
    port map (
            O => \N__65931\,
            I => \N__65928\
        );

    \I__15317\ : LocalMux
    port map (
            O => \N__65928\,
            I => \N__65924\
        );

    \I__15316\ : InMux
    port map (
            O => \N__65927\,
            I => \N__65921\
        );

    \I__15315\ : Span4Mux_v
    port map (
            O => \N__65924\,
            I => \N__65918\
        );

    \I__15314\ : LocalMux
    port map (
            O => \N__65921\,
            I => \N__65915\
        );

    \I__15313\ : Span4Mux_h
    port map (
            O => \N__65918\,
            I => \N__65910\
        );

    \I__15312\ : Span4Mux_v
    port map (
            O => \N__65915\,
            I => \N__65910\
        );

    \I__15311\ : Span4Mux_v
    port map (
            O => \N__65910\,
            I => \N__65907\
        );

    \I__15310\ : Odrv4
    port map (
            O => \N__65907\,
            I => \c0.n24527\
        );

    \I__15309\ : InMux
    port map (
            O => \N__65904\,
            I => \N__65899\
        );

    \I__15308\ : InMux
    port map (
            O => \N__65903\,
            I => \N__65896\
        );

    \I__15307\ : CascadeMux
    port map (
            O => \N__65902\,
            I => \N__65893\
        );

    \I__15306\ : LocalMux
    port map (
            O => \N__65899\,
            I => \N__65888\
        );

    \I__15305\ : LocalMux
    port map (
            O => \N__65896\,
            I => \N__65888\
        );

    \I__15304\ : InMux
    port map (
            O => \N__65893\,
            I => \N__65885\
        );

    \I__15303\ : Span4Mux_h
    port map (
            O => \N__65888\,
            I => \N__65881\
        );

    \I__15302\ : LocalMux
    port map (
            O => \N__65885\,
            I => \N__65878\
        );

    \I__15301\ : InMux
    port map (
            O => \N__65884\,
            I => \N__65875\
        );

    \I__15300\ : Span4Mux_h
    port map (
            O => \N__65881\,
            I => \N__65872\
        );

    \I__15299\ : Span4Mux_h
    port map (
            O => \N__65878\,
            I => \N__65869\
        );

    \I__15298\ : LocalMux
    port map (
            O => \N__65875\,
            I => data_in_frame_21_3
        );

    \I__15297\ : Odrv4
    port map (
            O => \N__65872\,
            I => data_in_frame_21_3
        );

    \I__15296\ : Odrv4
    port map (
            O => \N__65869\,
            I => data_in_frame_21_3
        );

    \I__15295\ : InMux
    port map (
            O => \N__65862\,
            I => \N__65858\
        );

    \I__15294\ : InMux
    port map (
            O => \N__65861\,
            I => \N__65855\
        );

    \I__15293\ : LocalMux
    port map (
            O => \N__65858\,
            I => \N__65850\
        );

    \I__15292\ : LocalMux
    port map (
            O => \N__65855\,
            I => \N__65847\
        );

    \I__15291\ : InMux
    port map (
            O => \N__65854\,
            I => \N__65841\
        );

    \I__15290\ : InMux
    port map (
            O => \N__65853\,
            I => \N__65841\
        );

    \I__15289\ : Span4Mux_v
    port map (
            O => \N__65850\,
            I => \N__65836\
        );

    \I__15288\ : Span4Mux_h
    port map (
            O => \N__65847\,
            I => \N__65836\
        );

    \I__15287\ : InMux
    port map (
            O => \N__65846\,
            I => \N__65832\
        );

    \I__15286\ : LocalMux
    port map (
            O => \N__65841\,
            I => \N__65829\
        );

    \I__15285\ : Span4Mux_h
    port map (
            O => \N__65836\,
            I => \N__65826\
        );

    \I__15284\ : InMux
    port map (
            O => \N__65835\,
            I => \N__65823\
        );

    \I__15283\ : LocalMux
    port map (
            O => \N__65832\,
            I => \c0.n21344\
        );

    \I__15282\ : Odrv4
    port map (
            O => \N__65829\,
            I => \c0.n21344\
        );

    \I__15281\ : Odrv4
    port map (
            O => \N__65826\,
            I => \c0.n21344\
        );

    \I__15280\ : LocalMux
    port map (
            O => \N__65823\,
            I => \c0.n21344\
        );

    \I__15279\ : InMux
    port map (
            O => \N__65814\,
            I => \N__65811\
        );

    \I__15278\ : LocalMux
    port map (
            O => \N__65811\,
            I => \N__65808\
        );

    \I__15277\ : Odrv4
    port map (
            O => \N__65808\,
            I => \c0.n42_adj_4589\
        );

    \I__15276\ : InMux
    port map (
            O => \N__65805\,
            I => \N__65802\
        );

    \I__15275\ : LocalMux
    port map (
            O => \N__65802\,
            I => \N__65799\
        );

    \I__15274\ : Span4Mux_v
    port map (
            O => \N__65799\,
            I => \N__65795\
        );

    \I__15273\ : InMux
    port map (
            O => \N__65798\,
            I => \N__65792\
        );

    \I__15272\ : Odrv4
    port map (
            O => \N__65795\,
            I => \c0.n22_adj_4243\
        );

    \I__15271\ : LocalMux
    port map (
            O => \N__65792\,
            I => \c0.n22_adj_4243\
        );

    \I__15270\ : InMux
    port map (
            O => \N__65787\,
            I => \N__65783\
        );

    \I__15269\ : InMux
    port map (
            O => \N__65786\,
            I => \N__65780\
        );

    \I__15268\ : LocalMux
    port map (
            O => \N__65783\,
            I => \N__65776\
        );

    \I__15267\ : LocalMux
    port map (
            O => \N__65780\,
            I => \N__65773\
        );

    \I__15266\ : CascadeMux
    port map (
            O => \N__65779\,
            I => \N__65769\
        );

    \I__15265\ : Span4Mux_v
    port map (
            O => \N__65776\,
            I => \N__65766\
        );

    \I__15264\ : Span4Mux_h
    port map (
            O => \N__65773\,
            I => \N__65763\
        );

    \I__15263\ : InMux
    port map (
            O => \N__65772\,
            I => \N__65760\
        );

    \I__15262\ : InMux
    port map (
            O => \N__65769\,
            I => \N__65757\
        );

    \I__15261\ : Odrv4
    port map (
            O => \N__65766\,
            I => \c0.n13738\
        );

    \I__15260\ : Odrv4
    port map (
            O => \N__65763\,
            I => \c0.n13738\
        );

    \I__15259\ : LocalMux
    port map (
            O => \N__65760\,
            I => \c0.n13738\
        );

    \I__15258\ : LocalMux
    port map (
            O => \N__65757\,
            I => \c0.n13738\
        );

    \I__15257\ : CascadeMux
    port map (
            O => \N__65748\,
            I => \N__65744\
        );

    \I__15256\ : CascadeMux
    port map (
            O => \N__65747\,
            I => \N__65741\
        );

    \I__15255\ : InMux
    port map (
            O => \N__65744\,
            I => \N__65738\
        );

    \I__15254\ : InMux
    port map (
            O => \N__65741\,
            I => \N__65735\
        );

    \I__15253\ : LocalMux
    port map (
            O => \N__65738\,
            I => \N__65732\
        );

    \I__15252\ : LocalMux
    port map (
            O => \N__65735\,
            I => \N__65729\
        );

    \I__15251\ : Span4Mux_h
    port map (
            O => \N__65732\,
            I => \N__65726\
        );

    \I__15250\ : Odrv12
    port map (
            O => \N__65729\,
            I => \c0.n10_adj_4230\
        );

    \I__15249\ : Odrv4
    port map (
            O => \N__65726\,
            I => \c0.n10_adj_4230\
        );

    \I__15248\ : InMux
    port map (
            O => \N__65721\,
            I => \N__65718\
        );

    \I__15247\ : LocalMux
    port map (
            O => \N__65718\,
            I => \N__65714\
        );

    \I__15246\ : InMux
    port map (
            O => \N__65717\,
            I => \N__65711\
        );

    \I__15245\ : Odrv4
    port map (
            O => \N__65714\,
            I => \c0.n5_adj_4310\
        );

    \I__15244\ : LocalMux
    port map (
            O => \N__65711\,
            I => \c0.n5_adj_4310\
        );

    \I__15243\ : InMux
    port map (
            O => \N__65706\,
            I => \N__65698\
        );

    \I__15242\ : InMux
    port map (
            O => \N__65705\,
            I => \N__65698\
        );

    \I__15241\ : InMux
    port map (
            O => \N__65704\,
            I => \N__65691\
        );

    \I__15240\ : InMux
    port map (
            O => \N__65703\,
            I => \N__65691\
        );

    \I__15239\ : LocalMux
    port map (
            O => \N__65698\,
            I => \N__65688\
        );

    \I__15238\ : CascadeMux
    port map (
            O => \N__65697\,
            I => \N__65685\
        );

    \I__15237\ : CascadeMux
    port map (
            O => \N__65696\,
            I => \N__65682\
        );

    \I__15236\ : LocalMux
    port map (
            O => \N__65691\,
            I => \N__65679\
        );

    \I__15235\ : Span4Mux_v
    port map (
            O => \N__65688\,
            I => \N__65675\
        );

    \I__15234\ : InMux
    port map (
            O => \N__65685\,
            I => \N__65670\
        );

    \I__15233\ : InMux
    port map (
            O => \N__65682\,
            I => \N__65670\
        );

    \I__15232\ : Span4Mux_v
    port map (
            O => \N__65679\,
            I => \N__65667\
        );

    \I__15231\ : InMux
    port map (
            O => \N__65678\,
            I => \N__65664\
        );

    \I__15230\ : Odrv4
    port map (
            O => \N__65675\,
            I => \c0.data_in_frame_4_5\
        );

    \I__15229\ : LocalMux
    port map (
            O => \N__65670\,
            I => \c0.data_in_frame_4_5\
        );

    \I__15228\ : Odrv4
    port map (
            O => \N__65667\,
            I => \c0.data_in_frame_4_5\
        );

    \I__15227\ : LocalMux
    port map (
            O => \N__65664\,
            I => \c0.data_in_frame_4_5\
        );

    \I__15226\ : CascadeMux
    port map (
            O => \N__65655\,
            I => \N__65651\
        );

    \I__15225\ : InMux
    port map (
            O => \N__65654\,
            I => \N__65646\
        );

    \I__15224\ : InMux
    port map (
            O => \N__65651\,
            I => \N__65646\
        );

    \I__15223\ : LocalMux
    port map (
            O => \N__65646\,
            I => \N__65643\
        );

    \I__15222\ : Odrv12
    port map (
            O => \N__65643\,
            I => \c0.n23283\
        );

    \I__15221\ : InMux
    port map (
            O => \N__65640\,
            I => \N__65634\
        );

    \I__15220\ : InMux
    port map (
            O => \N__65639\,
            I => \N__65627\
        );

    \I__15219\ : InMux
    port map (
            O => \N__65638\,
            I => \N__65624\
        );

    \I__15218\ : InMux
    port map (
            O => \N__65637\,
            I => \N__65621\
        );

    \I__15217\ : LocalMux
    port map (
            O => \N__65634\,
            I => \N__65618\
        );

    \I__15216\ : InMux
    port map (
            O => \N__65633\,
            I => \N__65613\
        );

    \I__15215\ : InMux
    port map (
            O => \N__65632\,
            I => \N__65613\
        );

    \I__15214\ : InMux
    port map (
            O => \N__65631\,
            I => \N__65608\
        );

    \I__15213\ : InMux
    port map (
            O => \N__65630\,
            I => \N__65608\
        );

    \I__15212\ : LocalMux
    port map (
            O => \N__65627\,
            I => \c0.data_in_frame_8_7\
        );

    \I__15211\ : LocalMux
    port map (
            O => \N__65624\,
            I => \c0.data_in_frame_8_7\
        );

    \I__15210\ : LocalMux
    port map (
            O => \N__65621\,
            I => \c0.data_in_frame_8_7\
        );

    \I__15209\ : Odrv4
    port map (
            O => \N__65618\,
            I => \c0.data_in_frame_8_7\
        );

    \I__15208\ : LocalMux
    port map (
            O => \N__65613\,
            I => \c0.data_in_frame_8_7\
        );

    \I__15207\ : LocalMux
    port map (
            O => \N__65608\,
            I => \c0.data_in_frame_8_7\
        );

    \I__15206\ : InMux
    port map (
            O => \N__65595\,
            I => \N__65592\
        );

    \I__15205\ : LocalMux
    port map (
            O => \N__65592\,
            I => \N__65588\
        );

    \I__15204\ : InMux
    port map (
            O => \N__65591\,
            I => \N__65585\
        );

    \I__15203\ : Odrv12
    port map (
            O => \N__65588\,
            I => \c0.n20_adj_4260\
        );

    \I__15202\ : LocalMux
    port map (
            O => \N__65585\,
            I => \c0.n20_adj_4260\
        );

    \I__15201\ : CascadeMux
    port map (
            O => \N__65580\,
            I => \N__65577\
        );

    \I__15200\ : InMux
    port map (
            O => \N__65577\,
            I => \N__65573\
        );

    \I__15199\ : InMux
    port map (
            O => \N__65576\,
            I => \N__65570\
        );

    \I__15198\ : LocalMux
    port map (
            O => \N__65573\,
            I => \N__65567\
        );

    \I__15197\ : LocalMux
    port map (
            O => \N__65570\,
            I => \N__65564\
        );

    \I__15196\ : Span4Mux_h
    port map (
            O => \N__65567\,
            I => \N__65561\
        );

    \I__15195\ : Span4Mux_v
    port map (
            O => \N__65564\,
            I => \N__65558\
        );

    \I__15194\ : Odrv4
    port map (
            O => \N__65561\,
            I => \c0.n22803\
        );

    \I__15193\ : Odrv4
    port map (
            O => \N__65558\,
            I => \c0.n22803\
        );

    \I__15192\ : InMux
    port map (
            O => \N__65553\,
            I => \N__65550\
        );

    \I__15191\ : LocalMux
    port map (
            O => \N__65550\,
            I => \N__65546\
        );

    \I__15190\ : InMux
    port map (
            O => \N__65549\,
            I => \N__65543\
        );

    \I__15189\ : Odrv4
    port map (
            O => \N__65546\,
            I => \c0.n4_adj_4261\
        );

    \I__15188\ : LocalMux
    port map (
            O => \N__65543\,
            I => \c0.n4_adj_4261\
        );

    \I__15187\ : InMux
    port map (
            O => \N__65538\,
            I => \N__65535\
        );

    \I__15186\ : LocalMux
    port map (
            O => \N__65535\,
            I => \N__65532\
        );

    \I__15185\ : Span12Mux_h
    port map (
            O => \N__65532\,
            I => \N__65529\
        );

    \I__15184\ : Odrv12
    port map (
            O => \N__65529\,
            I => \c0.n31_adj_4743\
        );

    \I__15183\ : InMux
    port map (
            O => \N__65526\,
            I => \N__65522\
        );

    \I__15182\ : InMux
    port map (
            O => \N__65525\,
            I => \N__65519\
        );

    \I__15181\ : LocalMux
    port map (
            O => \N__65522\,
            I => \N__65516\
        );

    \I__15180\ : LocalMux
    port map (
            O => \N__65519\,
            I => \c0.n5813\
        );

    \I__15179\ : Odrv4
    port map (
            O => \N__65516\,
            I => \c0.n5813\
        );

    \I__15178\ : CascadeMux
    port map (
            O => \N__65511\,
            I => \N__65507\
        );

    \I__15177\ : CascadeMux
    port map (
            O => \N__65510\,
            I => \N__65504\
        );

    \I__15176\ : InMux
    port map (
            O => \N__65507\,
            I => \N__65501\
        );

    \I__15175\ : InMux
    port map (
            O => \N__65504\,
            I => \N__65498\
        );

    \I__15174\ : LocalMux
    port map (
            O => \N__65501\,
            I => \c0.n22602\
        );

    \I__15173\ : LocalMux
    port map (
            O => \N__65498\,
            I => \c0.n22602\
        );

    \I__15172\ : InMux
    port map (
            O => \N__65493\,
            I => \N__65489\
        );

    \I__15171\ : InMux
    port map (
            O => \N__65492\,
            I => \N__65486\
        );

    \I__15170\ : LocalMux
    port map (
            O => \N__65489\,
            I => \N__65481\
        );

    \I__15169\ : LocalMux
    port map (
            O => \N__65486\,
            I => \N__65481\
        );

    \I__15168\ : Span4Mux_v
    port map (
            O => \N__65481\,
            I => \N__65478\
        );

    \I__15167\ : Odrv4
    port map (
            O => \N__65478\,
            I => \c0.n11\
        );

    \I__15166\ : InMux
    port map (
            O => \N__65475\,
            I => \N__65472\
        );

    \I__15165\ : LocalMux
    port map (
            O => \N__65472\,
            I => \N__65469\
        );

    \I__15164\ : Odrv12
    port map (
            O => \N__65469\,
            I => \c0.n17_adj_4219\
        );

    \I__15163\ : CascadeMux
    port map (
            O => \N__65466\,
            I => \c0.n16_adj_4218_cascade_\
        );

    \I__15162\ : CascadeMux
    port map (
            O => \N__65463\,
            I => \c0.n13767_cascade_\
        );

    \I__15161\ : InMux
    port map (
            O => \N__65460\,
            I => \N__65457\
        );

    \I__15160\ : LocalMux
    port map (
            O => \N__65457\,
            I => \N__65454\
        );

    \I__15159\ : Span4Mux_v
    port map (
            O => \N__65454\,
            I => \N__65450\
        );

    \I__15158\ : InMux
    port map (
            O => \N__65453\,
            I => \N__65447\
        );

    \I__15157\ : Span4Mux_h
    port map (
            O => \N__65450\,
            I => \N__65444\
        );

    \I__15156\ : LocalMux
    port map (
            O => \N__65447\,
            I => \N__65441\
        );

    \I__15155\ : Odrv4
    port map (
            O => \N__65444\,
            I => \c0.n5965\
        );

    \I__15154\ : Odrv4
    port map (
            O => \N__65441\,
            I => \c0.n5965\
        );

    \I__15153\ : InMux
    port map (
            O => \N__65436\,
            I => \N__65430\
        );

    \I__15152\ : InMux
    port map (
            O => \N__65435\,
            I => \N__65430\
        );

    \I__15151\ : LocalMux
    port map (
            O => \N__65430\,
            I => \c0.n6_adj_4454\
        );

    \I__15150\ : InMux
    port map (
            O => \N__65427\,
            I => \N__65423\
        );

    \I__15149\ : CascadeMux
    port map (
            O => \N__65426\,
            I => \N__65420\
        );

    \I__15148\ : LocalMux
    port map (
            O => \N__65423\,
            I => \N__65416\
        );

    \I__15147\ : InMux
    port map (
            O => \N__65420\,
            I => \N__65413\
        );

    \I__15146\ : InMux
    port map (
            O => \N__65419\,
            I => \N__65410\
        );

    \I__15145\ : Span4Mux_v
    port map (
            O => \N__65416\,
            I => \N__65407\
        );

    \I__15144\ : LocalMux
    port map (
            O => \N__65413\,
            I => \N__65398\
        );

    \I__15143\ : LocalMux
    port map (
            O => \N__65410\,
            I => \N__65398\
        );

    \I__15142\ : Sp12to4
    port map (
            O => \N__65407\,
            I => \N__65398\
        );

    \I__15141\ : InMux
    port map (
            O => \N__65406\,
            I => \N__65395\
        );

    \I__15140\ : InMux
    port map (
            O => \N__65405\,
            I => \N__65392\
        );

    \I__15139\ : Odrv12
    port map (
            O => \N__65398\,
            I => \c0.data_in_frame_15_3\
        );

    \I__15138\ : LocalMux
    port map (
            O => \N__65395\,
            I => \c0.data_in_frame_15_3\
        );

    \I__15137\ : LocalMux
    port map (
            O => \N__65392\,
            I => \c0.data_in_frame_15_3\
        );

    \I__15136\ : InMux
    port map (
            O => \N__65385\,
            I => \N__65382\
        );

    \I__15135\ : LocalMux
    port map (
            O => \N__65382\,
            I => \N__65379\
        );

    \I__15134\ : Span4Mux_v
    port map (
            O => \N__65379\,
            I => \N__65376\
        );

    \I__15133\ : Span4Mux_v
    port map (
            O => \N__65376\,
            I => \N__65373\
        );

    \I__15132\ : Odrv4
    port map (
            O => \N__65373\,
            I => \c0.n23_adj_4665\
        );

    \I__15131\ : InMux
    port map (
            O => \N__65370\,
            I => \N__65365\
        );

    \I__15130\ : CascadeMux
    port map (
            O => \N__65369\,
            I => \N__65362\
        );

    \I__15129\ : CascadeMux
    port map (
            O => \N__65368\,
            I => \N__65359\
        );

    \I__15128\ : LocalMux
    port map (
            O => \N__65365\,
            I => \N__65356\
        );

    \I__15127\ : InMux
    port map (
            O => \N__65362\,
            I => \N__65353\
        );

    \I__15126\ : InMux
    port map (
            O => \N__65359\,
            I => \N__65350\
        );

    \I__15125\ : Span4Mux_h
    port map (
            O => \N__65356\,
            I => \N__65347\
        );

    \I__15124\ : LocalMux
    port map (
            O => \N__65353\,
            I => \N__65344\
        );

    \I__15123\ : LocalMux
    port map (
            O => \N__65350\,
            I => \c0.data_in_frame_15_2\
        );

    \I__15122\ : Odrv4
    port map (
            O => \N__65347\,
            I => \c0.data_in_frame_15_2\
        );

    \I__15121\ : Odrv4
    port map (
            O => \N__65344\,
            I => \c0.data_in_frame_15_2\
        );

    \I__15120\ : CascadeMux
    port map (
            O => \N__65337\,
            I => \N__65332\
        );

    \I__15119\ : InMux
    port map (
            O => \N__65336\,
            I => \N__65328\
        );

    \I__15118\ : InMux
    port map (
            O => \N__65335\,
            I => \N__65324\
        );

    \I__15117\ : InMux
    port map (
            O => \N__65332\,
            I => \N__65319\
        );

    \I__15116\ : InMux
    port map (
            O => \N__65331\,
            I => \N__65319\
        );

    \I__15115\ : LocalMux
    port map (
            O => \N__65328\,
            I => \N__65316\
        );

    \I__15114\ : InMux
    port map (
            O => \N__65327\,
            I => \N__65313\
        );

    \I__15113\ : LocalMux
    port map (
            O => \N__65324\,
            I => \c0.data_in_frame_8_5\
        );

    \I__15112\ : LocalMux
    port map (
            O => \N__65319\,
            I => \c0.data_in_frame_8_5\
        );

    \I__15111\ : Odrv4
    port map (
            O => \N__65316\,
            I => \c0.data_in_frame_8_5\
        );

    \I__15110\ : LocalMux
    port map (
            O => \N__65313\,
            I => \c0.data_in_frame_8_5\
        );

    \I__15109\ : CascadeMux
    port map (
            O => \N__65304\,
            I => \N__65301\
        );

    \I__15108\ : InMux
    port map (
            O => \N__65301\,
            I => \N__65298\
        );

    \I__15107\ : LocalMux
    port map (
            O => \N__65298\,
            I => \N__65292\
        );

    \I__15106\ : InMux
    port map (
            O => \N__65297\,
            I => \N__65287\
        );

    \I__15105\ : InMux
    port map (
            O => \N__65296\,
            I => \N__65287\
        );

    \I__15104\ : CascadeMux
    port map (
            O => \N__65295\,
            I => \N__65283\
        );

    \I__15103\ : Span4Mux_v
    port map (
            O => \N__65292\,
            I => \N__65278\
        );

    \I__15102\ : LocalMux
    port map (
            O => \N__65287\,
            I => \N__65278\
        );

    \I__15101\ : CascadeMux
    port map (
            O => \N__65286\,
            I => \N__65275\
        );

    \I__15100\ : InMux
    port map (
            O => \N__65283\,
            I => \N__65272\
        );

    \I__15099\ : Span4Mux_h
    port map (
            O => \N__65278\,
            I => \N__65269\
        );

    \I__15098\ : InMux
    port map (
            O => \N__65275\,
            I => \N__65266\
        );

    \I__15097\ : LocalMux
    port map (
            O => \N__65272\,
            I => \N__65263\
        );

    \I__15096\ : Span4Mux_h
    port map (
            O => \N__65269\,
            I => \N__65260\
        );

    \I__15095\ : LocalMux
    port map (
            O => \N__65266\,
            I => \c0.data_in_frame_11_1\
        );

    \I__15094\ : Odrv12
    port map (
            O => \N__65263\,
            I => \c0.data_in_frame_11_1\
        );

    \I__15093\ : Odrv4
    port map (
            O => \N__65260\,
            I => \c0.data_in_frame_11_1\
        );

    \I__15092\ : InMux
    port map (
            O => \N__65253\,
            I => \N__65250\
        );

    \I__15091\ : LocalMux
    port map (
            O => \N__65250\,
            I => \c0.n22176\
        );

    \I__15090\ : CascadeMux
    port map (
            O => \N__65247\,
            I => \c0.n28_adj_4637_cascade_\
        );

    \I__15089\ : InMux
    port map (
            O => \N__65244\,
            I => \N__65241\
        );

    \I__15088\ : LocalMux
    port map (
            O => \N__65241\,
            I => \c0.n24_adj_4636\
        );

    \I__15087\ : InMux
    port map (
            O => \N__65238\,
            I => \N__65235\
        );

    \I__15086\ : LocalMux
    port map (
            O => \N__65235\,
            I => \c0.n7_adj_4634\
        );

    \I__15085\ : InMux
    port map (
            O => \N__65232\,
            I => \N__65229\
        );

    \I__15084\ : LocalMux
    port map (
            O => \N__65229\,
            I => \c0.n16_adj_4635\
        );

    \I__15083\ : InMux
    port map (
            O => \N__65226\,
            I => \N__65223\
        );

    \I__15082\ : LocalMux
    port map (
            O => \N__65223\,
            I => \N__65217\
        );

    \I__15081\ : InMux
    port map (
            O => \N__65222\,
            I => \N__65214\
        );

    \I__15080\ : InMux
    port map (
            O => \N__65221\,
            I => \N__65209\
        );

    \I__15079\ : InMux
    port map (
            O => \N__65220\,
            I => \N__65209\
        );

    \I__15078\ : Odrv4
    port map (
            O => \N__65217\,
            I => \c0.n23406\
        );

    \I__15077\ : LocalMux
    port map (
            O => \N__65214\,
            I => \c0.n23406\
        );

    \I__15076\ : LocalMux
    port map (
            O => \N__65209\,
            I => \c0.n23406\
        );

    \I__15075\ : InMux
    port map (
            O => \N__65202\,
            I => \N__65197\
        );

    \I__15074\ : InMux
    port map (
            O => \N__65201\,
            I => \N__65194\
        );

    \I__15073\ : InMux
    port map (
            O => \N__65200\,
            I => \N__65190\
        );

    \I__15072\ : LocalMux
    port map (
            O => \N__65197\,
            I => \N__65185\
        );

    \I__15071\ : LocalMux
    port map (
            O => \N__65194\,
            I => \N__65185\
        );

    \I__15070\ : InMux
    port map (
            O => \N__65193\,
            I => \N__65181\
        );

    \I__15069\ : LocalMux
    port map (
            O => \N__65190\,
            I => \N__65178\
        );

    \I__15068\ : Span4Mux_h
    port map (
            O => \N__65185\,
            I => \N__65175\
        );

    \I__15067\ : InMux
    port map (
            O => \N__65184\,
            I => \N__65172\
        );

    \I__15066\ : LocalMux
    port map (
            O => \N__65181\,
            I => data_in_frame_6_4
        );

    \I__15065\ : Odrv12
    port map (
            O => \N__65178\,
            I => data_in_frame_6_4
        );

    \I__15064\ : Odrv4
    port map (
            O => \N__65175\,
            I => data_in_frame_6_4
        );

    \I__15063\ : LocalMux
    port map (
            O => \N__65172\,
            I => data_in_frame_6_4
        );

    \I__15062\ : CascadeMux
    port map (
            O => \N__65163\,
            I => \c0.n14_adj_4609_cascade_\
        );

    \I__15061\ : InMux
    port map (
            O => \N__65160\,
            I => \N__65157\
        );

    \I__15060\ : LocalMux
    port map (
            O => \N__65157\,
            I => \c0.n10_adj_4617\
        );

    \I__15059\ : InMux
    port map (
            O => \N__65154\,
            I => \N__65151\
        );

    \I__15058\ : LocalMux
    port map (
            O => \N__65151\,
            I => \N__65147\
        );

    \I__15057\ : InMux
    port map (
            O => \N__65150\,
            I => \N__65144\
        );

    \I__15056\ : Span4Mux_v
    port map (
            O => \N__65147\,
            I => \N__65140\
        );

    \I__15055\ : LocalMux
    port map (
            O => \N__65144\,
            I => \N__65137\
        );

    \I__15054\ : InMux
    port map (
            O => \N__65143\,
            I => \N__65134\
        );

    \I__15053\ : Odrv4
    port map (
            O => \N__65140\,
            I => \c0.n17\
        );

    \I__15052\ : Odrv12
    port map (
            O => \N__65137\,
            I => \c0.n17\
        );

    \I__15051\ : LocalMux
    port map (
            O => \N__65134\,
            I => \c0.n17\
        );

    \I__15050\ : InMux
    port map (
            O => \N__65127\,
            I => \N__65121\
        );

    \I__15049\ : InMux
    port map (
            O => \N__65126\,
            I => \N__65121\
        );

    \I__15048\ : LocalMux
    port map (
            O => \N__65121\,
            I => \N__65118\
        );

    \I__15047\ : Odrv12
    port map (
            O => \N__65118\,
            I => \c0.n8_adj_4216\
        );

    \I__15046\ : CascadeMux
    port map (
            O => \N__65115\,
            I => \c0.n12_cascade_\
        );

    \I__15045\ : InMux
    port map (
            O => \N__65112\,
            I => \N__65105\
        );

    \I__15044\ : InMux
    port map (
            O => \N__65111\,
            I => \N__65102\
        );

    \I__15043\ : InMux
    port map (
            O => \N__65110\,
            I => \N__65097\
        );

    \I__15042\ : InMux
    port map (
            O => \N__65109\,
            I => \N__65097\
        );

    \I__15041\ : InMux
    port map (
            O => \N__65108\,
            I => \N__65093\
        );

    \I__15040\ : LocalMux
    port map (
            O => \N__65105\,
            I => \N__65088\
        );

    \I__15039\ : LocalMux
    port map (
            O => \N__65102\,
            I => \N__65088\
        );

    \I__15038\ : LocalMux
    port map (
            O => \N__65097\,
            I => \N__65085\
        );

    \I__15037\ : InMux
    port map (
            O => \N__65096\,
            I => \N__65082\
        );

    \I__15036\ : LocalMux
    port map (
            O => \N__65093\,
            I => \N__65079\
        );

    \I__15035\ : Span4Mux_v
    port map (
            O => \N__65088\,
            I => \N__65074\
        );

    \I__15034\ : Span4Mux_h
    port map (
            O => \N__65085\,
            I => \N__65074\
        );

    \I__15033\ : LocalMux
    port map (
            O => \N__65082\,
            I => \N__65070\
        );

    \I__15032\ : Span12Mux_h
    port map (
            O => \N__65079\,
            I => \N__65065\
        );

    \I__15031\ : Span4Mux_h
    port map (
            O => \N__65074\,
            I => \N__65062\
        );

    \I__15030\ : InMux
    port map (
            O => \N__65073\,
            I => \N__65059\
        );

    \I__15029\ : Span4Mux_v
    port map (
            O => \N__65070\,
            I => \N__65056\
        );

    \I__15028\ : InMux
    port map (
            O => \N__65069\,
            I => \N__65051\
        );

    \I__15027\ : InMux
    port map (
            O => \N__65068\,
            I => \N__65051\
        );

    \I__15026\ : Odrv12
    port map (
            O => \N__65065\,
            I => \c0.data_in_frame_4_2\
        );

    \I__15025\ : Odrv4
    port map (
            O => \N__65062\,
            I => \c0.data_in_frame_4_2\
        );

    \I__15024\ : LocalMux
    port map (
            O => \N__65059\,
            I => \c0.data_in_frame_4_2\
        );

    \I__15023\ : Odrv4
    port map (
            O => \N__65056\,
            I => \c0.data_in_frame_4_2\
        );

    \I__15022\ : LocalMux
    port map (
            O => \N__65051\,
            I => \c0.data_in_frame_4_2\
        );

    \I__15021\ : CascadeMux
    port map (
            O => \N__65040\,
            I => \N__65036\
        );

    \I__15020\ : CascadeMux
    port map (
            O => \N__65039\,
            I => \N__65032\
        );

    \I__15019\ : InMux
    port map (
            O => \N__65036\,
            I => \N__65029\
        );

    \I__15018\ : CascadeMux
    port map (
            O => \N__65035\,
            I => \N__65026\
        );

    \I__15017\ : InMux
    port map (
            O => \N__65032\,
            I => \N__65023\
        );

    \I__15016\ : LocalMux
    port map (
            O => \N__65029\,
            I => \N__65020\
        );

    \I__15015\ : InMux
    port map (
            O => \N__65026\,
            I => \N__65017\
        );

    \I__15014\ : LocalMux
    port map (
            O => \N__65023\,
            I => \c0.data_in_frame_12_2\
        );

    \I__15013\ : Odrv4
    port map (
            O => \N__65020\,
            I => \c0.data_in_frame_12_2\
        );

    \I__15012\ : LocalMux
    port map (
            O => \N__65017\,
            I => \c0.data_in_frame_12_2\
        );

    \I__15011\ : InMux
    port map (
            O => \N__65010\,
            I => \N__65006\
        );

    \I__15010\ : InMux
    port map (
            O => \N__65009\,
            I => \N__65003\
        );

    \I__15009\ : LocalMux
    port map (
            O => \N__65006\,
            I => \N__65000\
        );

    \I__15008\ : LocalMux
    port map (
            O => \N__65003\,
            I => \N__64997\
        );

    \I__15007\ : Span4Mux_h
    port map (
            O => \N__65000\,
            I => \N__64994\
        );

    \I__15006\ : Odrv4
    port map (
            O => \N__64997\,
            I => \c0.n13809\
        );

    \I__15005\ : Odrv4
    port map (
            O => \N__64994\,
            I => \c0.n13809\
        );

    \I__15004\ : CascadeMux
    port map (
            O => \N__64989\,
            I => \N__64983\
        );

    \I__15003\ : InMux
    port map (
            O => \N__64988\,
            I => \N__64980\
        );

    \I__15002\ : CascadeMux
    port map (
            O => \N__64987\,
            I => \N__64977\
        );

    \I__15001\ : InMux
    port map (
            O => \N__64986\,
            I => \N__64974\
        );

    \I__15000\ : InMux
    port map (
            O => \N__64983\,
            I => \N__64971\
        );

    \I__14999\ : LocalMux
    port map (
            O => \N__64980\,
            I => \N__64968\
        );

    \I__14998\ : InMux
    port map (
            O => \N__64977\,
            I => \N__64962\
        );

    \I__14997\ : LocalMux
    port map (
            O => \N__64974\,
            I => \N__64959\
        );

    \I__14996\ : LocalMux
    port map (
            O => \N__64971\,
            I => \N__64956\
        );

    \I__14995\ : Span4Mux_v
    port map (
            O => \N__64968\,
            I => \N__64953\
        );

    \I__14994\ : InMux
    port map (
            O => \N__64967\,
            I => \N__64950\
        );

    \I__14993\ : CascadeMux
    port map (
            O => \N__64966\,
            I => \N__64947\
        );

    \I__14992\ : InMux
    port map (
            O => \N__64965\,
            I => \N__64944\
        );

    \I__14991\ : LocalMux
    port map (
            O => \N__64962\,
            I => \N__64939\
        );

    \I__14990\ : Span4Mux_v
    port map (
            O => \N__64959\,
            I => \N__64939\
        );

    \I__14989\ : Span4Mux_v
    port map (
            O => \N__64956\,
            I => \N__64936\
        );

    \I__14988\ : Span4Mux_h
    port map (
            O => \N__64953\,
            I => \N__64931\
        );

    \I__14987\ : LocalMux
    port map (
            O => \N__64950\,
            I => \N__64931\
        );

    \I__14986\ : InMux
    port map (
            O => \N__64947\,
            I => \N__64928\
        );

    \I__14985\ : LocalMux
    port map (
            O => \N__64944\,
            I => \N__64923\
        );

    \I__14984\ : Span4Mux_h
    port map (
            O => \N__64939\,
            I => \N__64923\
        );

    \I__14983\ : Odrv4
    port map (
            O => \N__64936\,
            I => \c0.data_in_frame_11_5\
        );

    \I__14982\ : Odrv4
    port map (
            O => \N__64931\,
            I => \c0.data_in_frame_11_5\
        );

    \I__14981\ : LocalMux
    port map (
            O => \N__64928\,
            I => \c0.data_in_frame_11_5\
        );

    \I__14980\ : Odrv4
    port map (
            O => \N__64923\,
            I => \c0.data_in_frame_11_5\
        );

    \I__14979\ : InMux
    port map (
            O => \N__64914\,
            I => \N__64911\
        );

    \I__14978\ : LocalMux
    port map (
            O => \N__64911\,
            I => \N__64908\
        );

    \I__14977\ : Span4Mux_v
    port map (
            O => \N__64908\,
            I => \N__64905\
        );

    \I__14976\ : Odrv4
    port map (
            O => \N__64905\,
            I => \c0.n22751\
        );

    \I__14975\ : CascadeMux
    port map (
            O => \N__64902\,
            I => \N__64898\
        );

    \I__14974\ : CascadeMux
    port map (
            O => \N__64901\,
            I => \N__64894\
        );

    \I__14973\ : InMux
    port map (
            O => \N__64898\,
            I => \N__64891\
        );

    \I__14972\ : InMux
    port map (
            O => \N__64897\,
            I => \N__64888\
        );

    \I__14971\ : InMux
    port map (
            O => \N__64894\,
            I => \N__64885\
        );

    \I__14970\ : LocalMux
    port map (
            O => \N__64891\,
            I => \N__64880\
        );

    \I__14969\ : LocalMux
    port map (
            O => \N__64888\,
            I => \N__64877\
        );

    \I__14968\ : LocalMux
    port map (
            O => \N__64885\,
            I => \N__64874\
        );

    \I__14967\ : InMux
    port map (
            O => \N__64884\,
            I => \N__64868\
        );

    \I__14966\ : InMux
    port map (
            O => \N__64883\,
            I => \N__64868\
        );

    \I__14965\ : Span4Mux_v
    port map (
            O => \N__64880\,
            I => \N__64863\
        );

    \I__14964\ : Span4Mux_h
    port map (
            O => \N__64877\,
            I => \N__64863\
        );

    \I__14963\ : Span4Mux_h
    port map (
            O => \N__64874\,
            I => \N__64860\
        );

    \I__14962\ : InMux
    port map (
            O => \N__64873\,
            I => \N__64857\
        );

    \I__14961\ : LocalMux
    port map (
            O => \N__64868\,
            I => \N__64854\
        );

    \I__14960\ : Span4Mux_h
    port map (
            O => \N__64863\,
            I => \N__64851\
        );

    \I__14959\ : Span4Mux_h
    port map (
            O => \N__64860\,
            I => \N__64848\
        );

    \I__14958\ : LocalMux
    port map (
            O => \N__64857\,
            I => data_in_frame_6_7
        );

    \I__14957\ : Odrv12
    port map (
            O => \N__64854\,
            I => data_in_frame_6_7
        );

    \I__14956\ : Odrv4
    port map (
            O => \N__64851\,
            I => data_in_frame_6_7
        );

    \I__14955\ : Odrv4
    port map (
            O => \N__64848\,
            I => data_in_frame_6_7
        );

    \I__14954\ : InMux
    port map (
            O => \N__64839\,
            I => \N__64835\
        );

    \I__14953\ : CascadeMux
    port map (
            O => \N__64838\,
            I => \N__64831\
        );

    \I__14952\ : LocalMux
    port map (
            O => \N__64835\,
            I => \N__64828\
        );

    \I__14951\ : InMux
    port map (
            O => \N__64834\,
            I => \N__64824\
        );

    \I__14950\ : InMux
    port map (
            O => \N__64831\,
            I => \N__64821\
        );

    \I__14949\ : Span4Mux_h
    port map (
            O => \N__64828\,
            I => \N__64814\
        );

    \I__14948\ : InMux
    port map (
            O => \N__64827\,
            I => \N__64811\
        );

    \I__14947\ : LocalMux
    port map (
            O => \N__64824\,
            I => \N__64808\
        );

    \I__14946\ : LocalMux
    port map (
            O => \N__64821\,
            I => \N__64805\
        );

    \I__14945\ : InMux
    port map (
            O => \N__64820\,
            I => \N__64796\
        );

    \I__14944\ : InMux
    port map (
            O => \N__64819\,
            I => \N__64796\
        );

    \I__14943\ : InMux
    port map (
            O => \N__64818\,
            I => \N__64796\
        );

    \I__14942\ : InMux
    port map (
            O => \N__64817\,
            I => \N__64796\
        );

    \I__14941\ : Span4Mux_h
    port map (
            O => \N__64814\,
            I => \N__64793\
        );

    \I__14940\ : LocalMux
    port map (
            O => \N__64811\,
            I => \N__64788\
        );

    \I__14939\ : Span12Mux_v
    port map (
            O => \N__64808\,
            I => \N__64788\
        );

    \I__14938\ : Odrv12
    port map (
            O => \N__64805\,
            I => \c0.data_in_frame_4_7\
        );

    \I__14937\ : LocalMux
    port map (
            O => \N__64796\,
            I => \c0.data_in_frame_4_7\
        );

    \I__14936\ : Odrv4
    port map (
            O => \N__64793\,
            I => \c0.data_in_frame_4_7\
        );

    \I__14935\ : Odrv12
    port map (
            O => \N__64788\,
            I => \c0.data_in_frame_4_7\
        );

    \I__14934\ : InMux
    port map (
            O => \N__64779\,
            I => \N__64774\
        );

    \I__14933\ : InMux
    port map (
            O => \N__64778\,
            I => \N__64769\
        );

    \I__14932\ : InMux
    port map (
            O => \N__64777\,
            I => \N__64765\
        );

    \I__14931\ : LocalMux
    port map (
            O => \N__64774\,
            I => \N__64761\
        );

    \I__14930\ : InMux
    port map (
            O => \N__64773\,
            I => \N__64756\
        );

    \I__14929\ : InMux
    port map (
            O => \N__64772\,
            I => \N__64756\
        );

    \I__14928\ : LocalMux
    port map (
            O => \N__64769\,
            I => \N__64752\
        );

    \I__14927\ : InMux
    port map (
            O => \N__64768\,
            I => \N__64749\
        );

    \I__14926\ : LocalMux
    port map (
            O => \N__64765\,
            I => \N__64746\
        );

    \I__14925\ : InMux
    port map (
            O => \N__64764\,
            I => \N__64743\
        );

    \I__14924\ : Span4Mux_v
    port map (
            O => \N__64761\,
            I => \N__64738\
        );

    \I__14923\ : LocalMux
    port map (
            O => \N__64756\,
            I => \N__64738\
        );

    \I__14922\ : CascadeMux
    port map (
            O => \N__64755\,
            I => \N__64734\
        );

    \I__14921\ : Span4Mux_h
    port map (
            O => \N__64752\,
            I => \N__64728\
        );

    \I__14920\ : LocalMux
    port map (
            O => \N__64749\,
            I => \N__64728\
        );

    \I__14919\ : Span4Mux_h
    port map (
            O => \N__64746\,
            I => \N__64725\
        );

    \I__14918\ : LocalMux
    port map (
            O => \N__64743\,
            I => \N__64719\
        );

    \I__14917\ : Span4Mux_h
    port map (
            O => \N__64738\,
            I => \N__64719\
        );

    \I__14916\ : InMux
    port map (
            O => \N__64737\,
            I => \N__64716\
        );

    \I__14915\ : InMux
    port map (
            O => \N__64734\,
            I => \N__64713\
        );

    \I__14914\ : InMux
    port map (
            O => \N__64733\,
            I => \N__64710\
        );

    \I__14913\ : Span4Mux_h
    port map (
            O => \N__64728\,
            I => \N__64705\
        );

    \I__14912\ : Span4Mux_h
    port map (
            O => \N__64725\,
            I => \N__64705\
        );

    \I__14911\ : InMux
    port map (
            O => \N__64724\,
            I => \N__64702\
        );

    \I__14910\ : Sp12to4
    port map (
            O => \N__64719\,
            I => \N__64697\
        );

    \I__14909\ : LocalMux
    port map (
            O => \N__64716\,
            I => \N__64697\
        );

    \I__14908\ : LocalMux
    port map (
            O => \N__64713\,
            I => \c0.data_in_frame_2_7\
        );

    \I__14907\ : LocalMux
    port map (
            O => \N__64710\,
            I => \c0.data_in_frame_2_7\
        );

    \I__14906\ : Odrv4
    port map (
            O => \N__64705\,
            I => \c0.data_in_frame_2_7\
        );

    \I__14905\ : LocalMux
    port map (
            O => \N__64702\,
            I => \c0.data_in_frame_2_7\
        );

    \I__14904\ : Odrv12
    port map (
            O => \N__64697\,
            I => \c0.data_in_frame_2_7\
        );

    \I__14903\ : CascadeMux
    port map (
            O => \N__64686\,
            I => \N__64683\
        );

    \I__14902\ : InMux
    port map (
            O => \N__64683\,
            I => \N__64680\
        );

    \I__14901\ : LocalMux
    port map (
            O => \N__64680\,
            I => \c0.n49\
        );

    \I__14900\ : InMux
    port map (
            O => \N__64677\,
            I => \N__64674\
        );

    \I__14899\ : LocalMux
    port map (
            O => \N__64674\,
            I => \N__64670\
        );

    \I__14898\ : InMux
    port map (
            O => \N__64673\,
            I => \N__64667\
        );

    \I__14897\ : Odrv12
    port map (
            O => \N__64670\,
            I => \c0.n23528\
        );

    \I__14896\ : LocalMux
    port map (
            O => \N__64667\,
            I => \c0.n23528\
        );

    \I__14895\ : InMux
    port map (
            O => \N__64662\,
            I => \N__64659\
        );

    \I__14894\ : LocalMux
    port map (
            O => \N__64659\,
            I => \N__64656\
        );

    \I__14893\ : Span4Mux_v
    port map (
            O => \N__64656\,
            I => \N__64652\
        );

    \I__14892\ : InMux
    port map (
            O => \N__64655\,
            I => \N__64649\
        );

    \I__14891\ : Span4Mux_h
    port map (
            O => \N__64652\,
            I => \N__64644\
        );

    \I__14890\ : LocalMux
    port map (
            O => \N__64649\,
            I => \N__64644\
        );

    \I__14889\ : Span4Mux_v
    port map (
            O => \N__64644\,
            I => \N__64641\
        );

    \I__14888\ : Odrv4
    port map (
            O => \N__64641\,
            I => \c0.n7_adj_4229\
        );

    \I__14887\ : InMux
    port map (
            O => \N__64638\,
            I => \N__64635\
        );

    \I__14886\ : LocalMux
    port map (
            O => \N__64635\,
            I => \N__64630\
        );

    \I__14885\ : InMux
    port map (
            O => \N__64634\,
            I => \N__64625\
        );

    \I__14884\ : InMux
    port map (
            O => \N__64633\,
            I => \N__64625\
        );

    \I__14883\ : Span12Mux_v
    port map (
            O => \N__64630\,
            I => \N__64622\
        );

    \I__14882\ : LocalMux
    port map (
            O => \N__64625\,
            I => \N__64619\
        );

    \I__14881\ : Odrv12
    port map (
            O => \N__64622\,
            I => \c0.data_out_frame_0__7__N_2743\
        );

    \I__14880\ : Odrv4
    port map (
            O => \N__64619\,
            I => \c0.data_out_frame_0__7__N_2743\
        );

    \I__14879\ : InMux
    port map (
            O => \N__64614\,
            I => \N__64610\
        );

    \I__14878\ : InMux
    port map (
            O => \N__64613\,
            I => \N__64607\
        );

    \I__14877\ : LocalMux
    port map (
            O => \N__64610\,
            I => \N__64602\
        );

    \I__14876\ : LocalMux
    port map (
            O => \N__64607\,
            I => \N__64599\
        );

    \I__14875\ : InMux
    port map (
            O => \N__64606\,
            I => \N__64596\
        );

    \I__14874\ : InMux
    port map (
            O => \N__64605\,
            I => \N__64593\
        );

    \I__14873\ : Span4Mux_v
    port map (
            O => \N__64602\,
            I => \N__64590\
        );

    \I__14872\ : Span4Mux_v
    port map (
            O => \N__64599\,
            I => \N__64585\
        );

    \I__14871\ : LocalMux
    port map (
            O => \N__64596\,
            I => \N__64585\
        );

    \I__14870\ : LocalMux
    port map (
            O => \N__64593\,
            I => \N__64582\
        );

    \I__14869\ : Span4Mux_h
    port map (
            O => \N__64590\,
            I => \N__64578\
        );

    \I__14868\ : Span4Mux_v
    port map (
            O => \N__64585\,
            I => \N__64573\
        );

    \I__14867\ : Span4Mux_v
    port map (
            O => \N__64582\,
            I => \N__64573\
        );

    \I__14866\ : InMux
    port map (
            O => \N__64581\,
            I => \N__64570\
        );

    \I__14865\ : Odrv4
    port map (
            O => \N__64578\,
            I => \c0.n13523\
        );

    \I__14864\ : Odrv4
    port map (
            O => \N__64573\,
            I => \c0.n13523\
        );

    \I__14863\ : LocalMux
    port map (
            O => \N__64570\,
            I => \c0.n13523\
        );

    \I__14862\ : InMux
    port map (
            O => \N__64563\,
            I => \N__64557\
        );

    \I__14861\ : InMux
    port map (
            O => \N__64562\,
            I => \N__64557\
        );

    \I__14860\ : LocalMux
    port map (
            O => \N__64557\,
            I => \c0.n47\
        );

    \I__14859\ : CascadeMux
    port map (
            O => \N__64554\,
            I => \N__64551\
        );

    \I__14858\ : InMux
    port map (
            O => \N__64551\,
            I => \N__64548\
        );

    \I__14857\ : LocalMux
    port map (
            O => \N__64548\,
            I => \c0.n10_adj_4664\
        );

    \I__14856\ : InMux
    port map (
            O => \N__64545\,
            I => \N__64541\
        );

    \I__14855\ : CascadeMux
    port map (
            O => \N__64544\,
            I => \N__64538\
        );

    \I__14854\ : LocalMux
    port map (
            O => \N__64541\,
            I => \N__64535\
        );

    \I__14853\ : InMux
    port map (
            O => \N__64538\,
            I => \N__64532\
        );

    \I__14852\ : Span4Mux_v
    port map (
            O => \N__64535\,
            I => \N__64524\
        );

    \I__14851\ : LocalMux
    port map (
            O => \N__64532\,
            I => \N__64524\
        );

    \I__14850\ : InMux
    port map (
            O => \N__64531\,
            I => \N__64521\
        );

    \I__14849\ : InMux
    port map (
            O => \N__64530\,
            I => \N__64516\
        );

    \I__14848\ : InMux
    port map (
            O => \N__64529\,
            I => \N__64516\
        );

    \I__14847\ : Span4Mux_v
    port map (
            O => \N__64524\,
            I => \N__64513\
        );

    \I__14846\ : LocalMux
    port map (
            O => \N__64521\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14845\ : LocalMux
    port map (
            O => \N__64516\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14844\ : Odrv4
    port map (
            O => \N__64513\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14843\ : InMux
    port map (
            O => \N__64506\,
            I => \N__64503\
        );

    \I__14842\ : LocalMux
    port map (
            O => \N__64503\,
            I => \N__64498\
        );

    \I__14841\ : CascadeMux
    port map (
            O => \N__64502\,
            I => \N__64495\
        );

    \I__14840\ : InMux
    port map (
            O => \N__64501\,
            I => \N__64492\
        );

    \I__14839\ : Span4Mux_v
    port map (
            O => \N__64498\,
            I => \N__64487\
        );

    \I__14838\ : InMux
    port map (
            O => \N__64495\,
            I => \N__64484\
        );

    \I__14837\ : LocalMux
    port map (
            O => \N__64492\,
            I => \N__64481\
        );

    \I__14836\ : InMux
    port map (
            O => \N__64491\,
            I => \N__64478\
        );

    \I__14835\ : InMux
    port map (
            O => \N__64490\,
            I => \N__64475\
        );

    \I__14834\ : Span4Mux_h
    port map (
            O => \N__64487\,
            I => \N__64472\
        );

    \I__14833\ : LocalMux
    port map (
            O => \N__64484\,
            I => \N__64465\
        );

    \I__14832\ : Span4Mux_v
    port map (
            O => \N__64481\,
            I => \N__64465\
        );

    \I__14831\ : LocalMux
    port map (
            O => \N__64478\,
            I => \N__64465\
        );

    \I__14830\ : LocalMux
    port map (
            O => \N__64475\,
            I => \c0.data_in_frame_7_0\
        );

    \I__14829\ : Odrv4
    port map (
            O => \N__64472\,
            I => \c0.data_in_frame_7_0\
        );

    \I__14828\ : Odrv4
    port map (
            O => \N__64465\,
            I => \c0.data_in_frame_7_0\
        );

    \I__14827\ : CascadeMux
    port map (
            O => \N__64458\,
            I => \N__64454\
        );

    \I__14826\ : InMux
    port map (
            O => \N__64457\,
            I => \N__64451\
        );

    \I__14825\ : InMux
    port map (
            O => \N__64454\,
            I => \N__64447\
        );

    \I__14824\ : LocalMux
    port map (
            O => \N__64451\,
            I => \N__64444\
        );

    \I__14823\ : CascadeMux
    port map (
            O => \N__64450\,
            I => \N__64441\
        );

    \I__14822\ : LocalMux
    port map (
            O => \N__64447\,
            I => \N__64437\
        );

    \I__14821\ : Span4Mux_h
    port map (
            O => \N__64444\,
            I => \N__64434\
        );

    \I__14820\ : InMux
    port map (
            O => \N__64441\,
            I => \N__64431\
        );

    \I__14819\ : InMux
    port map (
            O => \N__64440\,
            I => \N__64428\
        );

    \I__14818\ : Span4Mux_v
    port map (
            O => \N__64437\,
            I => \N__64423\
        );

    \I__14817\ : Span4Mux_h
    port map (
            O => \N__64434\,
            I => \N__64423\
        );

    \I__14816\ : LocalMux
    port map (
            O => \N__64431\,
            I => \c0.data_in_frame_7_5\
        );

    \I__14815\ : LocalMux
    port map (
            O => \N__64428\,
            I => \c0.data_in_frame_7_5\
        );

    \I__14814\ : Odrv4
    port map (
            O => \N__64423\,
            I => \c0.data_in_frame_7_5\
        );

    \I__14813\ : CascadeMux
    port map (
            O => \N__64416\,
            I => \c0.n22417_cascade_\
        );

    \I__14812\ : InMux
    port map (
            O => \N__64413\,
            I => \N__64410\
        );

    \I__14811\ : LocalMux
    port map (
            O => \N__64410\,
            I => \N__64406\
        );

    \I__14810\ : InMux
    port map (
            O => \N__64409\,
            I => \N__64403\
        );

    \I__14809\ : Span4Mux_h
    port map (
            O => \N__64406\,
            I => \N__64400\
        );

    \I__14808\ : LocalMux
    port map (
            O => \N__64403\,
            I => \N__64397\
        );

    \I__14807\ : Span4Mux_h
    port map (
            O => \N__64400\,
            I => \N__64394\
        );

    \I__14806\ : Odrv4
    port map (
            O => \N__64397\,
            I => \c0.n4_adj_4333\
        );

    \I__14805\ : Odrv4
    port map (
            O => \N__64394\,
            I => \c0.n4_adj_4333\
        );

    \I__14804\ : InMux
    port map (
            O => \N__64389\,
            I => \N__64386\
        );

    \I__14803\ : LocalMux
    port map (
            O => \N__64386\,
            I => \N__64383\
        );

    \I__14802\ : Span4Mux_h
    port map (
            O => \N__64383\,
            I => \N__64380\
        );

    \I__14801\ : Odrv4
    port map (
            O => \N__64380\,
            I => \c0.n86\
        );

    \I__14800\ : InMux
    port map (
            O => \N__64377\,
            I => \N__64374\
        );

    \I__14799\ : LocalMux
    port map (
            O => \N__64374\,
            I => \N__64370\
        );

    \I__14798\ : InMux
    port map (
            O => \N__64373\,
            I => \N__64367\
        );

    \I__14797\ : Span4Mux_h
    port map (
            O => \N__64370\,
            I => \N__64364\
        );

    \I__14796\ : LocalMux
    port map (
            O => \N__64367\,
            I => \N__64361\
        );

    \I__14795\ : Span4Mux_h
    port map (
            O => \N__64364\,
            I => \N__64355\
        );

    \I__14794\ : Span4Mux_v
    port map (
            O => \N__64361\,
            I => \N__64355\
        );

    \I__14793\ : InMux
    port map (
            O => \N__64360\,
            I => \N__64352\
        );

    \I__14792\ : Odrv4
    port map (
            O => \N__64355\,
            I => \c0.n13085\
        );

    \I__14791\ : LocalMux
    port map (
            O => \N__64352\,
            I => \c0.n13085\
        );

    \I__14790\ : InMux
    port map (
            O => \N__64347\,
            I => \N__64342\
        );

    \I__14789\ : InMux
    port map (
            O => \N__64346\,
            I => \N__64337\
        );

    \I__14788\ : InMux
    port map (
            O => \N__64345\,
            I => \N__64334\
        );

    \I__14787\ : LocalMux
    port map (
            O => \N__64342\,
            I => \N__64331\
        );

    \I__14786\ : InMux
    port map (
            O => \N__64341\,
            I => \N__64328\
        );

    \I__14785\ : InMux
    port map (
            O => \N__64340\,
            I => \N__64325\
        );

    \I__14784\ : LocalMux
    port map (
            O => \N__64337\,
            I => \N__64322\
        );

    \I__14783\ : LocalMux
    port map (
            O => \N__64334\,
            I => \N__64317\
        );

    \I__14782\ : Span4Mux_h
    port map (
            O => \N__64331\,
            I => \N__64317\
        );

    \I__14781\ : LocalMux
    port map (
            O => \N__64328\,
            I => \N__64314\
        );

    \I__14780\ : LocalMux
    port map (
            O => \N__64325\,
            I => \N__64311\
        );

    \I__14779\ : Span4Mux_v
    port map (
            O => \N__64322\,
            I => \N__64306\
        );

    \I__14778\ : Span4Mux_v
    port map (
            O => \N__64317\,
            I => \N__64306\
        );

    \I__14777\ : Span4Mux_h
    port map (
            O => \N__64314\,
            I => \N__64303\
        );

    \I__14776\ : Span4Mux_v
    port map (
            O => \N__64311\,
            I => \N__64300\
        );

    \I__14775\ : Odrv4
    port map (
            O => \N__64306\,
            I => \c0.n7_adj_4282\
        );

    \I__14774\ : Odrv4
    port map (
            O => \N__64303\,
            I => \c0.n7_adj_4282\
        );

    \I__14773\ : Odrv4
    port map (
            O => \N__64300\,
            I => \c0.n7_adj_4282\
        );

    \I__14772\ : InMux
    port map (
            O => \N__64293\,
            I => \N__64290\
        );

    \I__14771\ : LocalMux
    port map (
            O => \N__64290\,
            I => \c0.n50\
        );

    \I__14770\ : CascadeMux
    port map (
            O => \N__64287\,
            I => \n22121_cascade_\
        );

    \I__14769\ : CascadeMux
    port map (
            O => \N__64284\,
            I => \N__64280\
        );

    \I__14768\ : InMux
    port map (
            O => \N__64283\,
            I => \N__64275\
        );

    \I__14767\ : InMux
    port map (
            O => \N__64280\,
            I => \N__64275\
        );

    \I__14766\ : LocalMux
    port map (
            O => \N__64275\,
            I => data_in_frame_6_6
        );

    \I__14765\ : InMux
    port map (
            O => \N__64272\,
            I => \N__64269\
        );

    \I__14764\ : LocalMux
    port map (
            O => \N__64269\,
            I => \N__64266\
        );

    \I__14763\ : Span4Mux_h
    port map (
            O => \N__64266\,
            I => \N__64263\
        );

    \I__14762\ : Span4Mux_v
    port map (
            O => \N__64263\,
            I => \N__64256\
        );

    \I__14761\ : InMux
    port map (
            O => \N__64262\,
            I => \N__64251\
        );

    \I__14760\ : InMux
    port map (
            O => \N__64261\,
            I => \N__64251\
        );

    \I__14759\ : InMux
    port map (
            O => \N__64260\,
            I => \N__64246\
        );

    \I__14758\ : InMux
    port map (
            O => \N__64259\,
            I => \N__64246\
        );

    \I__14757\ : Odrv4
    port map (
            O => \N__64256\,
            I => \c0.data_in_frame_2_2\
        );

    \I__14756\ : LocalMux
    port map (
            O => \N__64251\,
            I => \c0.data_in_frame_2_2\
        );

    \I__14755\ : LocalMux
    port map (
            O => \N__64246\,
            I => \c0.data_in_frame_2_2\
        );

    \I__14754\ : CascadeMux
    port map (
            O => \N__64239\,
            I => \N__64236\
        );

    \I__14753\ : InMux
    port map (
            O => \N__64236\,
            I => \N__64233\
        );

    \I__14752\ : LocalMux
    port map (
            O => \N__64233\,
            I => \N__64230\
        );

    \I__14751\ : Span4Mux_v
    port map (
            O => \N__64230\,
            I => \N__64226\
        );

    \I__14750\ : CascadeMux
    port map (
            O => \N__64229\,
            I => \N__64223\
        );

    \I__14749\ : Span4Mux_h
    port map (
            O => \N__64226\,
            I => \N__64220\
        );

    \I__14748\ : InMux
    port map (
            O => \N__64223\,
            I => \N__64217\
        );

    \I__14747\ : Odrv4
    port map (
            O => \N__64220\,
            I => \c0.n4_adj_4211\
        );

    \I__14746\ : LocalMux
    port map (
            O => \N__64217\,
            I => \c0.n4_adj_4211\
        );

    \I__14745\ : InMux
    port map (
            O => \N__64212\,
            I => \N__64206\
        );

    \I__14744\ : InMux
    port map (
            O => \N__64211\,
            I => \N__64206\
        );

    \I__14743\ : LocalMux
    port map (
            O => \N__64206\,
            I => \c0.n22647\
        );

    \I__14742\ : CascadeMux
    port map (
            O => \N__64203\,
            I => \c0.n13904_cascade_\
        );

    \I__14741\ : InMux
    port map (
            O => \N__64200\,
            I => \N__64197\
        );

    \I__14740\ : LocalMux
    port map (
            O => \N__64197\,
            I => \c0.n21_adj_4327\
        );

    \I__14739\ : CascadeMux
    port map (
            O => \N__64194\,
            I => \c0.n19_adj_4324_cascade_\
        );

    \I__14738\ : InMux
    port map (
            O => \N__64191\,
            I => \N__64188\
        );

    \I__14737\ : LocalMux
    port map (
            O => \N__64188\,
            I => \N__64185\
        );

    \I__14736\ : Span4Mux_h
    port map (
            O => \N__64185\,
            I => \N__64182\
        );

    \I__14735\ : Odrv4
    port map (
            O => \N__64182\,
            I => \c0.n22417\
        );

    \I__14734\ : CascadeMux
    port map (
            O => \N__64179\,
            I => \N__64174\
        );

    \I__14733\ : InMux
    port map (
            O => \N__64178\,
            I => \N__64169\
        );

    \I__14732\ : InMux
    port map (
            O => \N__64177\,
            I => \N__64169\
        );

    \I__14731\ : InMux
    port map (
            O => \N__64174\,
            I => \N__64165\
        );

    \I__14730\ : LocalMux
    port map (
            O => \N__64169\,
            I => \N__64162\
        );

    \I__14729\ : CascadeMux
    port map (
            O => \N__64168\,
            I => \N__64159\
        );

    \I__14728\ : LocalMux
    port map (
            O => \N__64165\,
            I => \N__64153\
        );

    \I__14727\ : Span4Mux_v
    port map (
            O => \N__64162\,
            I => \N__64153\
        );

    \I__14726\ : InMux
    port map (
            O => \N__64159\,
            I => \N__64148\
        );

    \I__14725\ : InMux
    port map (
            O => \N__64158\,
            I => \N__64148\
        );

    \I__14724\ : Odrv4
    port map (
            O => \N__64153\,
            I => \c0.data_in_frame_24_1\
        );

    \I__14723\ : LocalMux
    port map (
            O => \N__64148\,
            I => \c0.data_in_frame_24_1\
        );

    \I__14722\ : InMux
    port map (
            O => \N__64143\,
            I => \N__64140\
        );

    \I__14721\ : LocalMux
    port map (
            O => \N__64140\,
            I => \N__64135\
        );

    \I__14720\ : CascadeMux
    port map (
            O => \N__64139\,
            I => \N__64130\
        );

    \I__14719\ : InMux
    port map (
            O => \N__64138\,
            I => \N__64127\
        );

    \I__14718\ : Span4Mux_v
    port map (
            O => \N__64135\,
            I => \N__64124\
        );

    \I__14717\ : InMux
    port map (
            O => \N__64134\,
            I => \N__64121\
        );

    \I__14716\ : InMux
    port map (
            O => \N__64133\,
            I => \N__64118\
        );

    \I__14715\ : InMux
    port map (
            O => \N__64130\,
            I => \N__64115\
        );

    \I__14714\ : LocalMux
    port map (
            O => \N__64127\,
            I => \N__64112\
        );

    \I__14713\ : Sp12to4
    port map (
            O => \N__64124\,
            I => \N__64107\
        );

    \I__14712\ : LocalMux
    port map (
            O => \N__64121\,
            I => \N__64107\
        );

    \I__14711\ : LocalMux
    port map (
            O => \N__64118\,
            I => \N__64104\
        );

    \I__14710\ : LocalMux
    port map (
            O => \N__64115\,
            I => \N__64099\
        );

    \I__14709\ : Span4Mux_h
    port map (
            O => \N__64112\,
            I => \N__64099\
        );

    \I__14708\ : Span12Mux_h
    port map (
            O => \N__64107\,
            I => \N__64096\
        );

    \I__14707\ : Odrv12
    port map (
            O => \N__64104\,
            I => \c0.data_in_frame_27_1\
        );

    \I__14706\ : Odrv4
    port map (
            O => \N__64099\,
            I => \c0.data_in_frame_27_1\
        );

    \I__14705\ : Odrv12
    port map (
            O => \N__64096\,
            I => \c0.data_in_frame_27_1\
        );

    \I__14704\ : InMux
    port map (
            O => \N__64089\,
            I => \N__64086\
        );

    \I__14703\ : LocalMux
    port map (
            O => \N__64086\,
            I => \N__64082\
        );

    \I__14702\ : InMux
    port map (
            O => \N__64085\,
            I => \N__64079\
        );

    \I__14701\ : Span4Mux_h
    port map (
            O => \N__64082\,
            I => \N__64076\
        );

    \I__14700\ : LocalMux
    port map (
            O => \N__64079\,
            I => \N__64073\
        );

    \I__14699\ : Odrv4
    port map (
            O => \N__64076\,
            I => \c0.n39_adj_4515\
        );

    \I__14698\ : Odrv4
    port map (
            O => \N__64073\,
            I => \c0.n39_adj_4515\
        );

    \I__14697\ : InMux
    port map (
            O => \N__64068\,
            I => \N__64065\
        );

    \I__14696\ : LocalMux
    port map (
            O => \N__64065\,
            I => \N__64062\
        );

    \I__14695\ : Odrv4
    port map (
            O => \N__64062\,
            I => \c0.n10_adj_4675\
        );

    \I__14694\ : CascadeMux
    port map (
            O => \N__64059\,
            I => \N__64056\
        );

    \I__14693\ : InMux
    port map (
            O => \N__64056\,
            I => \N__64053\
        );

    \I__14692\ : LocalMux
    port map (
            O => \N__64053\,
            I => \N__64050\
        );

    \I__14691\ : Span4Mux_v
    port map (
            O => \N__64050\,
            I => \N__64045\
        );

    \I__14690\ : InMux
    port map (
            O => \N__64049\,
            I => \N__64042\
        );

    \I__14689\ : CascadeMux
    port map (
            O => \N__64048\,
            I => \N__64039\
        );

    \I__14688\ : Span4Mux_v
    port map (
            O => \N__64045\,
            I => \N__64034\
        );

    \I__14687\ : LocalMux
    port map (
            O => \N__64042\,
            I => \N__64034\
        );

    \I__14686\ : InMux
    port map (
            O => \N__64039\,
            I => \N__64030\
        );

    \I__14685\ : Span4Mux_h
    port map (
            O => \N__64034\,
            I => \N__64027\
        );

    \I__14684\ : InMux
    port map (
            O => \N__64033\,
            I => \N__64024\
        );

    \I__14683\ : LocalMux
    port map (
            O => \N__64030\,
            I => \c0.data_in_frame_11_0\
        );

    \I__14682\ : Odrv4
    port map (
            O => \N__64027\,
            I => \c0.data_in_frame_11_0\
        );

    \I__14681\ : LocalMux
    port map (
            O => \N__64024\,
            I => \c0.data_in_frame_11_0\
        );

    \I__14680\ : InMux
    port map (
            O => \N__64017\,
            I => \N__64014\
        );

    \I__14679\ : LocalMux
    port map (
            O => \N__64014\,
            I => \N__64009\
        );

    \I__14678\ : CascadeMux
    port map (
            O => \N__64013\,
            I => \N__64003\
        );

    \I__14677\ : InMux
    port map (
            O => \N__64012\,
            I => \N__64000\
        );

    \I__14676\ : Span4Mux_h
    port map (
            O => \N__64009\,
            I => \N__63997\
        );

    \I__14675\ : InMux
    port map (
            O => \N__64008\,
            I => \N__63994\
        );

    \I__14674\ : InMux
    port map (
            O => \N__64007\,
            I => \N__63989\
        );

    \I__14673\ : InMux
    port map (
            O => \N__64006\,
            I => \N__63989\
        );

    \I__14672\ : InMux
    port map (
            O => \N__64003\,
            I => \N__63986\
        );

    \I__14671\ : LocalMux
    port map (
            O => \N__64000\,
            I => \N__63983\
        );

    \I__14670\ : Odrv4
    port map (
            O => \N__63997\,
            I => \c0.data_in_frame_4_6\
        );

    \I__14669\ : LocalMux
    port map (
            O => \N__63994\,
            I => \c0.data_in_frame_4_6\
        );

    \I__14668\ : LocalMux
    port map (
            O => \N__63989\,
            I => \c0.data_in_frame_4_6\
        );

    \I__14667\ : LocalMux
    port map (
            O => \N__63986\,
            I => \c0.data_in_frame_4_6\
        );

    \I__14666\ : Odrv4
    port map (
            O => \N__63983\,
            I => \c0.data_in_frame_4_6\
        );

    \I__14665\ : InMux
    port map (
            O => \N__63972\,
            I => \N__63969\
        );

    \I__14664\ : LocalMux
    port map (
            O => \N__63969\,
            I => \N__63966\
        );

    \I__14663\ : Span4Mux_h
    port map (
            O => \N__63966\,
            I => \N__63962\
        );

    \I__14662\ : InMux
    port map (
            O => \N__63965\,
            I => \N__63958\
        );

    \I__14661\ : Span4Mux_h
    port map (
            O => \N__63962\,
            I => \N__63955\
        );

    \I__14660\ : InMux
    port map (
            O => \N__63961\,
            I => \N__63952\
        );

    \I__14659\ : LocalMux
    port map (
            O => \N__63958\,
            I => \c0.data_in_frame_23_7\
        );

    \I__14658\ : Odrv4
    port map (
            O => \N__63955\,
            I => \c0.data_in_frame_23_7\
        );

    \I__14657\ : LocalMux
    port map (
            O => \N__63952\,
            I => \c0.data_in_frame_23_7\
        );

    \I__14656\ : CascadeMux
    port map (
            O => \N__63945\,
            I => \c0.n7_adj_4364_cascade_\
        );

    \I__14655\ : InMux
    port map (
            O => \N__63942\,
            I => \N__63939\
        );

    \I__14654\ : LocalMux
    port map (
            O => \N__63939\,
            I => \N__63936\
        );

    \I__14653\ : Span4Mux_h
    port map (
            O => \N__63936\,
            I => \N__63933\
        );

    \I__14652\ : Span4Mux_h
    port map (
            O => \N__63933\,
            I => \N__63929\
        );

    \I__14651\ : InMux
    port map (
            O => \N__63932\,
            I => \N__63926\
        );

    \I__14650\ : Odrv4
    port map (
            O => \N__63929\,
            I => \c0.n21426\
        );

    \I__14649\ : LocalMux
    port map (
            O => \N__63926\,
            I => \c0.n21426\
        );

    \I__14648\ : CascadeMux
    port map (
            O => \N__63921\,
            I => \c0.n23031_cascade_\
        );

    \I__14647\ : InMux
    port map (
            O => \N__63918\,
            I => \N__63914\
        );

    \I__14646\ : CascadeMux
    port map (
            O => \N__63917\,
            I => \N__63911\
        );

    \I__14645\ : LocalMux
    port map (
            O => \N__63914\,
            I => \N__63908\
        );

    \I__14644\ : InMux
    port map (
            O => \N__63911\,
            I => \N__63903\
        );

    \I__14643\ : Span4Mux_v
    port map (
            O => \N__63908\,
            I => \N__63900\
        );

    \I__14642\ : InMux
    port map (
            O => \N__63907\,
            I => \N__63895\
        );

    \I__14641\ : InMux
    port map (
            O => \N__63906\,
            I => \N__63895\
        );

    \I__14640\ : LocalMux
    port map (
            O => \N__63903\,
            I => \c0.data_in_frame_25_7\
        );

    \I__14639\ : Odrv4
    port map (
            O => \N__63900\,
            I => \c0.data_in_frame_25_7\
        );

    \I__14638\ : LocalMux
    port map (
            O => \N__63895\,
            I => \c0.data_in_frame_25_7\
        );

    \I__14637\ : CascadeMux
    port map (
            O => \N__63888\,
            I => \N__63885\
        );

    \I__14636\ : InMux
    port map (
            O => \N__63885\,
            I => \N__63882\
        );

    \I__14635\ : LocalMux
    port map (
            O => \N__63882\,
            I => \N__63879\
        );

    \I__14634\ : Span4Mux_h
    port map (
            O => \N__63879\,
            I => \N__63874\
        );

    \I__14633\ : CascadeMux
    port map (
            O => \N__63878\,
            I => \N__63871\
        );

    \I__14632\ : CascadeMux
    port map (
            O => \N__63877\,
            I => \N__63868\
        );

    \I__14631\ : Span4Mux_h
    port map (
            O => \N__63874\,
            I => \N__63865\
        );

    \I__14630\ : InMux
    port map (
            O => \N__63871\,
            I => \N__63860\
        );

    \I__14629\ : InMux
    port map (
            O => \N__63868\,
            I => \N__63860\
        );

    \I__14628\ : Odrv4
    port map (
            O => \N__63865\,
            I => \c0.data_in_frame_26_5\
        );

    \I__14627\ : LocalMux
    port map (
            O => \N__63860\,
            I => \c0.data_in_frame_26_5\
        );

    \I__14626\ : InMux
    port map (
            O => \N__63855\,
            I => \N__63852\
        );

    \I__14625\ : LocalMux
    port map (
            O => \N__63852\,
            I => \c0.n24482\
        );

    \I__14624\ : InMux
    port map (
            O => \N__63849\,
            I => \N__63843\
        );

    \I__14623\ : InMux
    port map (
            O => \N__63848\,
            I => \N__63838\
        );

    \I__14622\ : InMux
    port map (
            O => \N__63847\,
            I => \N__63838\
        );

    \I__14621\ : InMux
    port map (
            O => \N__63846\,
            I => \N__63835\
        );

    \I__14620\ : LocalMux
    port map (
            O => \N__63843\,
            I => \c0.n23031\
        );

    \I__14619\ : LocalMux
    port map (
            O => \N__63838\,
            I => \c0.n23031\
        );

    \I__14618\ : LocalMux
    port map (
            O => \N__63835\,
            I => \c0.n23031\
        );

    \I__14617\ : CascadeMux
    port map (
            O => \N__63828\,
            I => \N__63825\
        );

    \I__14616\ : InMux
    port map (
            O => \N__63825\,
            I => \N__63821\
        );

    \I__14615\ : InMux
    port map (
            O => \N__63824\,
            I => \N__63818\
        );

    \I__14614\ : LocalMux
    port map (
            O => \N__63821\,
            I => \c0.data_in_frame_28_2\
        );

    \I__14613\ : LocalMux
    port map (
            O => \N__63818\,
            I => \c0.data_in_frame_28_2\
        );

    \I__14612\ : CascadeMux
    port map (
            O => \N__63813\,
            I => \c0.n36_adj_4460_cascade_\
        );

    \I__14611\ : InMux
    port map (
            O => \N__63810\,
            I => \N__63807\
        );

    \I__14610\ : LocalMux
    port map (
            O => \N__63807\,
            I => \c0.n41_adj_4511\
        );

    \I__14609\ : InMux
    port map (
            O => \N__63804\,
            I => \N__63798\
        );

    \I__14608\ : InMux
    port map (
            O => \N__63803\,
            I => \N__63798\
        );

    \I__14607\ : LocalMux
    port map (
            O => \N__63798\,
            I => \N__63795\
        );

    \I__14606\ : Odrv4
    port map (
            O => \N__63795\,
            I => \c0.n6_adj_4459\
        );

    \I__14605\ : InMux
    port map (
            O => \N__63792\,
            I => \N__63783\
        );

    \I__14604\ : InMux
    port map (
            O => \N__63791\,
            I => \N__63779\
        );

    \I__14603\ : InMux
    port map (
            O => \N__63790\,
            I => \N__63776\
        );

    \I__14602\ : InMux
    port map (
            O => \N__63789\,
            I => \N__63771\
        );

    \I__14601\ : InMux
    port map (
            O => \N__63788\,
            I => \N__63771\
        );

    \I__14600\ : InMux
    port map (
            O => \N__63787\,
            I => \N__63768\
        );

    \I__14599\ : InMux
    port map (
            O => \N__63786\,
            I => \N__63765\
        );

    \I__14598\ : LocalMux
    port map (
            O => \N__63783\,
            I => \N__63762\
        );

    \I__14597\ : InMux
    port map (
            O => \N__63782\,
            I => \N__63759\
        );

    \I__14596\ : LocalMux
    port map (
            O => \N__63779\,
            I => \N__63750\
        );

    \I__14595\ : LocalMux
    port map (
            O => \N__63776\,
            I => \N__63750\
        );

    \I__14594\ : LocalMux
    port map (
            O => \N__63771\,
            I => \N__63750\
        );

    \I__14593\ : LocalMux
    port map (
            O => \N__63768\,
            I => \N__63750\
        );

    \I__14592\ : LocalMux
    port map (
            O => \N__63765\,
            I => \c0.n22426\
        );

    \I__14591\ : Odrv4
    port map (
            O => \N__63762\,
            I => \c0.n22426\
        );

    \I__14590\ : LocalMux
    port map (
            O => \N__63759\,
            I => \c0.n22426\
        );

    \I__14589\ : Odrv4
    port map (
            O => \N__63750\,
            I => \c0.n22426\
        );

    \I__14588\ : CascadeMux
    port map (
            O => \N__63741\,
            I => \N__63736\
        );

    \I__14587\ : CascadeMux
    port map (
            O => \N__63740\,
            I => \N__63732\
        );

    \I__14586\ : CascadeMux
    port map (
            O => \N__63739\,
            I => \N__63728\
        );

    \I__14585\ : InMux
    port map (
            O => \N__63736\,
            I => \N__63724\
        );

    \I__14584\ : InMux
    port map (
            O => \N__63735\,
            I => \N__63719\
        );

    \I__14583\ : InMux
    port map (
            O => \N__63732\,
            I => \N__63719\
        );

    \I__14582\ : CascadeMux
    port map (
            O => \N__63731\,
            I => \N__63716\
        );

    \I__14581\ : InMux
    port map (
            O => \N__63728\,
            I => \N__63713\
        );

    \I__14580\ : InMux
    port map (
            O => \N__63727\,
            I => \N__63710\
        );

    \I__14579\ : LocalMux
    port map (
            O => \N__63724\,
            I => \N__63705\
        );

    \I__14578\ : LocalMux
    port map (
            O => \N__63719\,
            I => \N__63705\
        );

    \I__14577\ : InMux
    port map (
            O => \N__63716\,
            I => \N__63702\
        );

    \I__14576\ : LocalMux
    port map (
            O => \N__63713\,
            I => \N__63697\
        );

    \I__14575\ : LocalMux
    port map (
            O => \N__63710\,
            I => \N__63697\
        );

    \I__14574\ : Span4Mux_h
    port map (
            O => \N__63705\,
            I => \N__63694\
        );

    \I__14573\ : LocalMux
    port map (
            O => \N__63702\,
            I => \c0.data_in_frame_26_1\
        );

    \I__14572\ : Odrv4
    port map (
            O => \N__63697\,
            I => \c0.data_in_frame_26_1\
        );

    \I__14571\ : Odrv4
    port map (
            O => \N__63694\,
            I => \c0.data_in_frame_26_1\
        );

    \I__14570\ : CascadeMux
    port map (
            O => \N__63687\,
            I => \N__63681\
        );

    \I__14569\ : InMux
    port map (
            O => \N__63686\,
            I => \N__63677\
        );

    \I__14568\ : InMux
    port map (
            O => \N__63685\,
            I => \N__63672\
        );

    \I__14567\ : InMux
    port map (
            O => \N__63684\,
            I => \N__63672\
        );

    \I__14566\ : InMux
    port map (
            O => \N__63681\,
            I => \N__63669\
        );

    \I__14565\ : InMux
    port map (
            O => \N__63680\,
            I => \N__63666\
        );

    \I__14564\ : LocalMux
    port map (
            O => \N__63677\,
            I => \c0.n22340\
        );

    \I__14563\ : LocalMux
    port map (
            O => \N__63672\,
            I => \c0.n22340\
        );

    \I__14562\ : LocalMux
    port map (
            O => \N__63669\,
            I => \c0.n22340\
        );

    \I__14561\ : LocalMux
    port map (
            O => \N__63666\,
            I => \c0.n22340\
        );

    \I__14560\ : CascadeMux
    port map (
            O => \N__63657\,
            I => \c0.n5_adj_4472_cascade_\
        );

    \I__14559\ : InMux
    port map (
            O => \N__63654\,
            I => \N__63650\
        );

    \I__14558\ : InMux
    port map (
            O => \N__63653\,
            I => \N__63647\
        );

    \I__14557\ : LocalMux
    port map (
            O => \N__63650\,
            I => \c0.n21010\
        );

    \I__14556\ : LocalMux
    port map (
            O => \N__63647\,
            I => \c0.n21010\
        );

    \I__14555\ : InMux
    port map (
            O => \N__63642\,
            I => \N__63639\
        );

    \I__14554\ : LocalMux
    port map (
            O => \N__63639\,
            I => \c0.n24_adj_4496\
        );

    \I__14553\ : InMux
    port map (
            O => \N__63636\,
            I => \N__63631\
        );

    \I__14552\ : InMux
    port map (
            O => \N__63635\,
            I => \N__63626\
        );

    \I__14551\ : InMux
    port map (
            O => \N__63634\,
            I => \N__63626\
        );

    \I__14550\ : LocalMux
    port map (
            O => \N__63631\,
            I => \c0.n34_adj_4361\
        );

    \I__14549\ : LocalMux
    port map (
            O => \N__63626\,
            I => \c0.n34_adj_4361\
        );

    \I__14548\ : CascadeMux
    port map (
            O => \N__63621\,
            I => \c0.n57_cascade_\
        );

    \I__14547\ : InMux
    port map (
            O => \N__63618\,
            I => \N__63615\
        );

    \I__14546\ : LocalMux
    port map (
            O => \N__63615\,
            I => \c0.n48_adj_4365\
        );

    \I__14545\ : CascadeMux
    port map (
            O => \N__63612\,
            I => \c0.n21426_cascade_\
        );

    \I__14544\ : InMux
    port map (
            O => \N__63609\,
            I => \N__63606\
        );

    \I__14543\ : LocalMux
    port map (
            O => \N__63606\,
            I => \N__63603\
        );

    \I__14542\ : Span4Mux_h
    port map (
            O => \N__63603\,
            I => \N__63600\
        );

    \I__14541\ : Span4Mux_h
    port map (
            O => \N__63600\,
            I => \N__63595\
        );

    \I__14540\ : InMux
    port map (
            O => \N__63599\,
            I => \N__63592\
        );

    \I__14539\ : InMux
    port map (
            O => \N__63598\,
            I => \N__63589\
        );

    \I__14538\ : Odrv4
    port map (
            O => \N__63595\,
            I => \c0.n23032\
        );

    \I__14537\ : LocalMux
    port map (
            O => \N__63592\,
            I => \c0.n23032\
        );

    \I__14536\ : LocalMux
    port map (
            O => \N__63589\,
            I => \c0.n23032\
        );

    \I__14535\ : CascadeMux
    port map (
            O => \N__63582\,
            I => \c0.n23032_cascade_\
        );

    \I__14534\ : InMux
    port map (
            O => \N__63579\,
            I => \N__63576\
        );

    \I__14533\ : LocalMux
    port map (
            O => \N__63576\,
            I => \N__63573\
        );

    \I__14532\ : Odrv4
    port map (
            O => \N__63573\,
            I => \c0.n25456\
        );

    \I__14531\ : CascadeMux
    port map (
            O => \N__63570\,
            I => \c0.n23209_cascade_\
        );

    \I__14530\ : InMux
    port map (
            O => \N__63567\,
            I => \N__63564\
        );

    \I__14529\ : LocalMux
    port map (
            O => \N__63564\,
            I => \c0.n56_adj_4479\
        );

    \I__14528\ : InMux
    port map (
            O => \N__63561\,
            I => \N__63557\
        );

    \I__14527\ : InMux
    port map (
            O => \N__63560\,
            I => \N__63554\
        );

    \I__14526\ : LocalMux
    port map (
            O => \N__63557\,
            I => \N__63551\
        );

    \I__14525\ : LocalMux
    port map (
            O => \N__63554\,
            I => \N__63548\
        );

    \I__14524\ : Odrv12
    port map (
            O => \N__63551\,
            I => \c0.n21299\
        );

    \I__14523\ : Odrv12
    port map (
            O => \N__63548\,
            I => \c0.n21299\
        );

    \I__14522\ : InMux
    port map (
            O => \N__63543\,
            I => \N__63539\
        );

    \I__14521\ : InMux
    port map (
            O => \N__63542\,
            I => \N__63536\
        );

    \I__14520\ : LocalMux
    port map (
            O => \N__63539\,
            I => \N__63533\
        );

    \I__14519\ : LocalMux
    port map (
            O => \N__63536\,
            I => \N__63530\
        );

    \I__14518\ : Span4Mux_h
    port map (
            O => \N__63533\,
            I => \N__63527\
        );

    \I__14517\ : Span4Mux_v
    port map (
            O => \N__63530\,
            I => \N__63524\
        );

    \I__14516\ : Span4Mux_v
    port map (
            O => \N__63527\,
            I => \N__63517\
        );

    \I__14515\ : Span4Mux_h
    port map (
            O => \N__63524\,
            I => \N__63517\
        );

    \I__14514\ : InMux
    port map (
            O => \N__63523\,
            I => \N__63512\
        );

    \I__14513\ : InMux
    port map (
            O => \N__63522\,
            I => \N__63512\
        );

    \I__14512\ : Odrv4
    port map (
            O => \N__63517\,
            I => data_in_frame_22_6
        );

    \I__14511\ : LocalMux
    port map (
            O => \N__63512\,
            I => data_in_frame_22_6
        );

    \I__14510\ : InMux
    port map (
            O => \N__63507\,
            I => \N__63503\
        );

    \I__14509\ : InMux
    port map (
            O => \N__63506\,
            I => \N__63500\
        );

    \I__14508\ : LocalMux
    port map (
            O => \N__63503\,
            I => \N__63496\
        );

    \I__14507\ : LocalMux
    port map (
            O => \N__63500\,
            I => \N__63493\
        );

    \I__14506\ : InMux
    port map (
            O => \N__63499\,
            I => \N__63490\
        );

    \I__14505\ : Span4Mux_h
    port map (
            O => \N__63496\,
            I => \N__63487\
        );

    \I__14504\ : Span4Mux_h
    port map (
            O => \N__63493\,
            I => \N__63484\
        );

    \I__14503\ : LocalMux
    port map (
            O => \N__63490\,
            I => \N__63479\
        );

    \I__14502\ : Span4Mux_h
    port map (
            O => \N__63487\,
            I => \N__63479\
        );

    \I__14501\ : Odrv4
    port map (
            O => \N__63484\,
            I => data_in_frame_22_0
        );

    \I__14500\ : Odrv4
    port map (
            O => \N__63479\,
            I => data_in_frame_22_0
        );

    \I__14499\ : CascadeMux
    port map (
            O => \N__63474\,
            I => \c0.n12559_cascade_\
        );

    \I__14498\ : InMux
    port map (
            O => \N__63471\,
            I => \N__63468\
        );

    \I__14497\ : LocalMux
    port map (
            O => \N__63468\,
            I => \N__63465\
        );

    \I__14496\ : Span12Mux_v
    port map (
            O => \N__63465\,
            I => \N__63461\
        );

    \I__14495\ : InMux
    port map (
            O => \N__63464\,
            I => \N__63458\
        );

    \I__14494\ : Odrv12
    port map (
            O => \N__63461\,
            I => \c0.n22375\
        );

    \I__14493\ : LocalMux
    port map (
            O => \N__63458\,
            I => \c0.n22375\
        );

    \I__14492\ : InMux
    port map (
            O => \N__63453\,
            I => \N__63450\
        );

    \I__14491\ : LocalMux
    port map (
            O => \N__63450\,
            I => \N__63447\
        );

    \I__14490\ : Span4Mux_h
    port map (
            O => \N__63447\,
            I => \N__63444\
        );

    \I__14489\ : Odrv4
    port map (
            O => \N__63444\,
            I => \c0.n24451\
        );

    \I__14488\ : CascadeMux
    port map (
            O => \N__63441\,
            I => \N__63437\
        );

    \I__14487\ : InMux
    port map (
            O => \N__63440\,
            I => \N__63434\
        );

    \I__14486\ : InMux
    port map (
            O => \N__63437\,
            I => \N__63431\
        );

    \I__14485\ : LocalMux
    port map (
            O => \N__63434\,
            I => \N__63427\
        );

    \I__14484\ : LocalMux
    port map (
            O => \N__63431\,
            I => \N__63424\
        );

    \I__14483\ : InMux
    port map (
            O => \N__63430\,
            I => \N__63421\
        );

    \I__14482\ : Span4Mux_h
    port map (
            O => \N__63427\,
            I => \N__63418\
        );

    \I__14481\ : Span4Mux_h
    port map (
            O => \N__63424\,
            I => \N__63413\
        );

    \I__14480\ : LocalMux
    port map (
            O => \N__63421\,
            I => \N__63413\
        );

    \I__14479\ : Span4Mux_h
    port map (
            O => \N__63418\,
            I => \N__63409\
        );

    \I__14478\ : Span4Mux_v
    port map (
            O => \N__63413\,
            I => \N__63406\
        );

    \I__14477\ : CascadeMux
    port map (
            O => \N__63412\,
            I => \N__63403\
        );

    \I__14476\ : Sp12to4
    port map (
            O => \N__63409\,
            I => \N__63400\
        );

    \I__14475\ : Span4Mux_h
    port map (
            O => \N__63406\,
            I => \N__63397\
        );

    \I__14474\ : InMux
    port map (
            O => \N__63403\,
            I => \N__63394\
        );

    \I__14473\ : Span12Mux_v
    port map (
            O => \N__63400\,
            I => \N__63391\
        );

    \I__14472\ : Span4Mux_v
    port map (
            O => \N__63397\,
            I => \N__63388\
        );

    \I__14471\ : LocalMux
    port map (
            O => \N__63394\,
            I => \c0.data_in_frame_19_1\
        );

    \I__14470\ : Odrv12
    port map (
            O => \N__63391\,
            I => \c0.data_in_frame_19_1\
        );

    \I__14469\ : Odrv4
    port map (
            O => \N__63388\,
            I => \c0.data_in_frame_19_1\
        );

    \I__14468\ : InMux
    port map (
            O => \N__63381\,
            I => \N__63375\
        );

    \I__14467\ : InMux
    port map (
            O => \N__63380\,
            I => \N__63372\
        );

    \I__14466\ : InMux
    port map (
            O => \N__63379\,
            I => \N__63367\
        );

    \I__14465\ : InMux
    port map (
            O => \N__63378\,
            I => \N__63367\
        );

    \I__14464\ : LocalMux
    port map (
            O => \N__63375\,
            I => \N__63364\
        );

    \I__14463\ : LocalMux
    port map (
            O => \N__63372\,
            I => \N__63359\
        );

    \I__14462\ : LocalMux
    port map (
            O => \N__63367\,
            I => \N__63359\
        );

    \I__14461\ : Span4Mux_v
    port map (
            O => \N__63364\,
            I => \N__63356\
        );

    \I__14460\ : Span4Mux_v
    port map (
            O => \N__63359\,
            I => \N__63353\
        );

    \I__14459\ : Odrv4
    port map (
            O => \N__63356\,
            I => \c0.n6215\
        );

    \I__14458\ : Odrv4
    port map (
            O => \N__63353\,
            I => \c0.n6215\
        );

    \I__14457\ : CascadeMux
    port map (
            O => \N__63348\,
            I => \N__63342\
        );

    \I__14456\ : InMux
    port map (
            O => \N__63347\,
            I => \N__63339\
        );

    \I__14455\ : InMux
    port map (
            O => \N__63346\,
            I => \N__63332\
        );

    \I__14454\ : InMux
    port map (
            O => \N__63345\,
            I => \N__63332\
        );

    \I__14453\ : InMux
    port map (
            O => \N__63342\,
            I => \N__63332\
        );

    \I__14452\ : LocalMux
    port map (
            O => \N__63339\,
            I => \N__63329\
        );

    \I__14451\ : LocalMux
    port map (
            O => \N__63332\,
            I => \N__63325\
        );

    \I__14450\ : Span4Mux_h
    port map (
            O => \N__63329\,
            I => \N__63322\
        );

    \I__14449\ : InMux
    port map (
            O => \N__63328\,
            I => \N__63319\
        );

    \I__14448\ : Sp12to4
    port map (
            O => \N__63325\,
            I => \N__63316\
        );

    \I__14447\ : Span4Mux_h
    port map (
            O => \N__63322\,
            I => \N__63313\
        );

    \I__14446\ : LocalMux
    port map (
            O => \N__63319\,
            I => \c0.data_in_frame_19_2\
        );

    \I__14445\ : Odrv12
    port map (
            O => \N__63316\,
            I => \c0.data_in_frame_19_2\
        );

    \I__14444\ : Odrv4
    port map (
            O => \N__63313\,
            I => \c0.data_in_frame_19_2\
        );

    \I__14443\ : InMux
    port map (
            O => \N__63306\,
            I => \N__63303\
        );

    \I__14442\ : LocalMux
    port map (
            O => \N__63303\,
            I => \N__63300\
        );

    \I__14441\ : Span4Mux_h
    port map (
            O => \N__63300\,
            I => \N__63296\
        );

    \I__14440\ : InMux
    port map (
            O => \N__63299\,
            I => \N__63292\
        );

    \I__14439\ : Span4Mux_h
    port map (
            O => \N__63296\,
            I => \N__63289\
        );

    \I__14438\ : InMux
    port map (
            O => \N__63295\,
            I => \N__63286\
        );

    \I__14437\ : LocalMux
    port map (
            O => \N__63292\,
            I => \c0.n21275\
        );

    \I__14436\ : Odrv4
    port map (
            O => \N__63289\,
            I => \c0.n21275\
        );

    \I__14435\ : LocalMux
    port map (
            O => \N__63286\,
            I => \c0.n21275\
        );

    \I__14434\ : CascadeMux
    port map (
            O => \N__63279\,
            I => \c0.n21275_cascade_\
        );

    \I__14433\ : InMux
    port map (
            O => \N__63276\,
            I => \N__63273\
        );

    \I__14432\ : LocalMux
    port map (
            O => \N__63273\,
            I => \N__63270\
        );

    \I__14431\ : Span4Mux_v
    port map (
            O => \N__63270\,
            I => \N__63267\
        );

    \I__14430\ : Odrv4
    port map (
            O => \N__63267\,
            I => \c0.n14_adj_4440\
        );

    \I__14429\ : InMux
    port map (
            O => \N__63264\,
            I => \N__63260\
        );

    \I__14428\ : InMux
    port map (
            O => \N__63263\,
            I => \N__63257\
        );

    \I__14427\ : LocalMux
    port map (
            O => \N__63260\,
            I => \N__63254\
        );

    \I__14426\ : LocalMux
    port map (
            O => \N__63257\,
            I => \N__63251\
        );

    \I__14425\ : Span4Mux_h
    port map (
            O => \N__63254\,
            I => \N__63246\
        );

    \I__14424\ : Span4Mux_v
    port map (
            O => \N__63251\,
            I => \N__63246\
        );

    \I__14423\ : Odrv4
    port map (
            O => \N__63246\,
            I => \c0.n63_adj_4516\
        );

    \I__14422\ : InMux
    port map (
            O => \N__63243\,
            I => \N__63237\
        );

    \I__14421\ : InMux
    port map (
            O => \N__63242\,
            I => \N__63234\
        );

    \I__14420\ : InMux
    port map (
            O => \N__63241\,
            I => \N__63231\
        );

    \I__14419\ : InMux
    port map (
            O => \N__63240\,
            I => \N__63227\
        );

    \I__14418\ : LocalMux
    port map (
            O => \N__63237\,
            I => \N__63223\
        );

    \I__14417\ : LocalMux
    port map (
            O => \N__63234\,
            I => \N__63218\
        );

    \I__14416\ : LocalMux
    port map (
            O => \N__63231\,
            I => \N__63218\
        );

    \I__14415\ : InMux
    port map (
            O => \N__63230\,
            I => \N__63215\
        );

    \I__14414\ : LocalMux
    port map (
            O => \N__63227\,
            I => \N__63212\
        );

    \I__14413\ : InMux
    port map (
            O => \N__63226\,
            I => \N__63208\
        );

    \I__14412\ : Span4Mux_v
    port map (
            O => \N__63223\,
            I => \N__63203\
        );

    \I__14411\ : Span4Mux_v
    port map (
            O => \N__63218\,
            I => \N__63203\
        );

    \I__14410\ : LocalMux
    port map (
            O => \N__63215\,
            I => \N__63198\
        );

    \I__14409\ : Span4Mux_v
    port map (
            O => \N__63212\,
            I => \N__63198\
        );

    \I__14408\ : InMux
    port map (
            O => \N__63211\,
            I => \N__63195\
        );

    \I__14407\ : LocalMux
    port map (
            O => \N__63208\,
            I => \N__63192\
        );

    \I__14406\ : Span4Mux_h
    port map (
            O => \N__63203\,
            I => \N__63185\
        );

    \I__14405\ : Span4Mux_h
    port map (
            O => \N__63198\,
            I => \N__63185\
        );

    \I__14404\ : LocalMux
    port map (
            O => \N__63195\,
            I => \N__63185\
        );

    \I__14403\ : Span4Mux_h
    port map (
            O => \N__63192\,
            I => \N__63182\
        );

    \I__14402\ : Span4Mux_v
    port map (
            O => \N__63185\,
            I => \N__63179\
        );

    \I__14401\ : Odrv4
    port map (
            O => \N__63182\,
            I => \c0.n14189\
        );

    \I__14400\ : Odrv4
    port map (
            O => \N__63179\,
            I => \c0.n14189\
        );

    \I__14399\ : CascadeMux
    port map (
            O => \N__63174\,
            I => \N__63171\
        );

    \I__14398\ : InMux
    port map (
            O => \N__63171\,
            I => \N__63167\
        );

    \I__14397\ : InMux
    port map (
            O => \N__63170\,
            I => \N__63164\
        );

    \I__14396\ : LocalMux
    port map (
            O => \N__63167\,
            I => \c0.n46\
        );

    \I__14395\ : LocalMux
    port map (
            O => \N__63164\,
            I => \c0.n46\
        );

    \I__14394\ : CascadeMux
    port map (
            O => \N__63159\,
            I => \c0.n46_cascade_\
        );

    \I__14393\ : CascadeMux
    port map (
            O => \N__63156\,
            I => \N__63153\
        );

    \I__14392\ : InMux
    port map (
            O => \N__63153\,
            I => \N__63149\
        );

    \I__14391\ : InMux
    port map (
            O => \N__63152\,
            I => \N__63145\
        );

    \I__14390\ : LocalMux
    port map (
            O => \N__63149\,
            I => \N__63142\
        );

    \I__14389\ : InMux
    port map (
            O => \N__63148\,
            I => \N__63138\
        );

    \I__14388\ : LocalMux
    port map (
            O => \N__63145\,
            I => \N__63135\
        );

    \I__14387\ : Span4Mux_h
    port map (
            O => \N__63142\,
            I => \N__63132\
        );

    \I__14386\ : InMux
    port map (
            O => \N__63141\,
            I => \N__63129\
        );

    \I__14385\ : LocalMux
    port map (
            O => \N__63138\,
            I => \c0.data_in_frame_12_7\
        );

    \I__14384\ : Odrv4
    port map (
            O => \N__63135\,
            I => \c0.data_in_frame_12_7\
        );

    \I__14383\ : Odrv4
    port map (
            O => \N__63132\,
            I => \c0.data_in_frame_12_7\
        );

    \I__14382\ : LocalMux
    port map (
            O => \N__63129\,
            I => \c0.data_in_frame_12_7\
        );

    \I__14381\ : InMux
    port map (
            O => \N__63120\,
            I => \N__63117\
        );

    \I__14380\ : LocalMux
    port map (
            O => \N__63117\,
            I => \c0.n25_adj_4579\
        );

    \I__14379\ : CascadeMux
    port map (
            O => \N__63114\,
            I => \c0.n25_adj_4579_cascade_\
        );

    \I__14378\ : CascadeMux
    port map (
            O => \N__63111\,
            I => \c0.n23433_cascade_\
        );

    \I__14377\ : InMux
    port map (
            O => \N__63108\,
            I => \N__63102\
        );

    \I__14376\ : InMux
    port map (
            O => \N__63107\,
            I => \N__63102\
        );

    \I__14375\ : LocalMux
    port map (
            O => \N__63102\,
            I => \N__63099\
        );

    \I__14374\ : Odrv12
    port map (
            O => \N__63099\,
            I => \c0.n18_adj_4580\
        );

    \I__14373\ : InMux
    port map (
            O => \N__63096\,
            I => \N__63093\
        );

    \I__14372\ : LocalMux
    port map (
            O => \N__63093\,
            I => \c0.n24_adj_4655\
        );

    \I__14371\ : InMux
    port map (
            O => \N__63090\,
            I => \N__63086\
        );

    \I__14370\ : CascadeMux
    port map (
            O => \N__63089\,
            I => \N__63083\
        );

    \I__14369\ : LocalMux
    port map (
            O => \N__63086\,
            I => \N__63080\
        );

    \I__14368\ : InMux
    port map (
            O => \N__63083\,
            I => \N__63077\
        );

    \I__14367\ : Span4Mux_h
    port map (
            O => \N__63080\,
            I => \N__63074\
        );

    \I__14366\ : LocalMux
    port map (
            O => \N__63077\,
            I => \c0.n41_adj_4592\
        );

    \I__14365\ : Odrv4
    port map (
            O => \N__63074\,
            I => \c0.n41_adj_4592\
        );

    \I__14364\ : InMux
    port map (
            O => \N__63069\,
            I => \N__63066\
        );

    \I__14363\ : LocalMux
    port map (
            O => \N__63066\,
            I => \c0.n43_adj_4661\
        );

    \I__14362\ : CascadeMux
    port map (
            O => \N__63063\,
            I => \N__63060\
        );

    \I__14361\ : InMux
    port map (
            O => \N__63060\,
            I => \N__63057\
        );

    \I__14360\ : LocalMux
    port map (
            O => \N__63057\,
            I => \N__63054\
        );

    \I__14359\ : Odrv4
    port map (
            O => \N__63054\,
            I => \c0.n44_adj_4588\
        );

    \I__14358\ : InMux
    port map (
            O => \N__63051\,
            I => \N__63048\
        );

    \I__14357\ : LocalMux
    port map (
            O => \N__63048\,
            I => \N__63045\
        );

    \I__14356\ : Span4Mux_h
    port map (
            O => \N__63045\,
            I => \N__63042\
        );

    \I__14355\ : Odrv4
    port map (
            O => \N__63042\,
            I => \c0.n39_adj_4341\
        );

    \I__14354\ : InMux
    port map (
            O => \N__63039\,
            I => \N__63036\
        );

    \I__14353\ : LocalMux
    port map (
            O => \N__63036\,
            I => \N__63033\
        );

    \I__14352\ : Span4Mux_v
    port map (
            O => \N__63033\,
            I => \N__63029\
        );

    \I__14351\ : InMux
    port map (
            O => \N__63032\,
            I => \N__63026\
        );

    \I__14350\ : Odrv4
    port map (
            O => \N__63029\,
            I => \c0.n22205\
        );

    \I__14349\ : LocalMux
    port map (
            O => \N__63026\,
            I => \c0.n22205\
        );

    \I__14348\ : CascadeMux
    port map (
            O => \N__63021\,
            I => \c0.n50_adj_4340_cascade_\
        );

    \I__14347\ : InMux
    port map (
            O => \N__63018\,
            I => \N__63015\
        );

    \I__14346\ : LocalMux
    port map (
            O => \N__63015\,
            I => \N__63012\
        );

    \I__14345\ : Span4Mux_v
    port map (
            O => \N__63012\,
            I => \N__63008\
        );

    \I__14344\ : InMux
    port map (
            O => \N__63011\,
            I => \N__63005\
        );

    \I__14343\ : Span4Mux_h
    port map (
            O => \N__63008\,
            I => \N__63002\
        );

    \I__14342\ : LocalMux
    port map (
            O => \N__63005\,
            I => \N__62999\
        );

    \I__14341\ : Odrv4
    port map (
            O => \N__63002\,
            I => \c0.n5_adj_4486\
        );

    \I__14340\ : Odrv4
    port map (
            O => \N__62999\,
            I => \c0.n5_adj_4486\
        );

    \I__14339\ : InMux
    port map (
            O => \N__62994\,
            I => \N__62991\
        );

    \I__14338\ : LocalMux
    port map (
            O => \N__62991\,
            I => \N__62988\
        );

    \I__14337\ : Odrv4
    port map (
            O => \N__62988\,
            I => \c0.n20467\
        );

    \I__14336\ : CascadeMux
    port map (
            O => \N__62985\,
            I => \c0.n20467_cascade_\
        );

    \I__14335\ : CascadeMux
    port map (
            O => \N__62982\,
            I => \N__62977\
        );

    \I__14334\ : InMux
    port map (
            O => \N__62981\,
            I => \N__62974\
        );

    \I__14333\ : CascadeMux
    port map (
            O => \N__62980\,
            I => \N__62971\
        );

    \I__14332\ : InMux
    port map (
            O => \N__62977\,
            I => \N__62968\
        );

    \I__14331\ : LocalMux
    port map (
            O => \N__62974\,
            I => \N__62965\
        );

    \I__14330\ : InMux
    port map (
            O => \N__62971\,
            I => \N__62962\
        );

    \I__14329\ : LocalMux
    port map (
            O => \N__62968\,
            I => \N__62959\
        );

    \I__14328\ : Span4Mux_h
    port map (
            O => \N__62965\,
            I => \N__62956\
        );

    \I__14327\ : LocalMux
    port map (
            O => \N__62962\,
            I => \N__62953\
        );

    \I__14326\ : Span4Mux_v
    port map (
            O => \N__62959\,
            I => \N__62948\
        );

    \I__14325\ : Span4Mux_v
    port map (
            O => \N__62956\,
            I => \N__62948\
        );

    \I__14324\ : Odrv4
    port map (
            O => \N__62953\,
            I => \c0.n6404\
        );

    \I__14323\ : Odrv4
    port map (
            O => \N__62948\,
            I => \c0.n6404\
        );

    \I__14322\ : CascadeMux
    port map (
            O => \N__62943\,
            I => \c0.n17_adj_4354_cascade_\
        );

    \I__14321\ : InMux
    port map (
            O => \N__62940\,
            I => \N__62934\
        );

    \I__14320\ : InMux
    port map (
            O => \N__62939\,
            I => \N__62934\
        );

    \I__14319\ : LocalMux
    port map (
            O => \N__62934\,
            I => \c0.n10_adj_4630\
        );

    \I__14318\ : InMux
    port map (
            O => \N__62931\,
            I => \N__62928\
        );

    \I__14317\ : LocalMux
    port map (
            O => \N__62928\,
            I => \N__62924\
        );

    \I__14316\ : CascadeMux
    port map (
            O => \N__62927\,
            I => \N__62921\
        );

    \I__14315\ : Span4Mux_h
    port map (
            O => \N__62924\,
            I => \N__62916\
        );

    \I__14314\ : InMux
    port map (
            O => \N__62921\,
            I => \N__62911\
        );

    \I__14313\ : InMux
    port map (
            O => \N__62920\,
            I => \N__62911\
        );

    \I__14312\ : InMux
    port map (
            O => \N__62919\,
            I => \N__62908\
        );

    \I__14311\ : Span4Mux_v
    port map (
            O => \N__62916\,
            I => \N__62905\
        );

    \I__14310\ : LocalMux
    port map (
            O => \N__62911\,
            I => \N__62900\
        );

    \I__14309\ : LocalMux
    port map (
            O => \N__62908\,
            I => \N__62900\
        );

    \I__14308\ : Odrv4
    port map (
            O => \N__62905\,
            I => \c0.n23523\
        );

    \I__14307\ : Odrv12
    port map (
            O => \N__62900\,
            I => \c0.n23523\
        );

    \I__14306\ : InMux
    port map (
            O => \N__62895\,
            I => \N__62891\
        );

    \I__14305\ : InMux
    port map (
            O => \N__62894\,
            I => \N__62888\
        );

    \I__14304\ : LocalMux
    port map (
            O => \N__62891\,
            I => \N__62881\
        );

    \I__14303\ : LocalMux
    port map (
            O => \N__62888\,
            I => \N__62881\
        );

    \I__14302\ : InMux
    port map (
            O => \N__62887\,
            I => \N__62876\
        );

    \I__14301\ : InMux
    port map (
            O => \N__62886\,
            I => \N__62876\
        );

    \I__14300\ : Span4Mux_v
    port map (
            O => \N__62881\,
            I => \N__62872\
        );

    \I__14299\ : LocalMux
    port map (
            O => \N__62876\,
            I => \N__62869\
        );

    \I__14298\ : InMux
    port map (
            O => \N__62875\,
            I => \N__62866\
        );

    \I__14297\ : Odrv4
    port map (
            O => \N__62872\,
            I => \c0.n6_adj_4209\
        );

    \I__14296\ : Odrv12
    port map (
            O => \N__62869\,
            I => \c0.n6_adj_4209\
        );

    \I__14295\ : LocalMux
    port map (
            O => \N__62866\,
            I => \c0.n6_adj_4209\
        );

    \I__14294\ : CascadeMux
    port map (
            O => \N__62859\,
            I => \N__62855\
        );

    \I__14293\ : InMux
    port map (
            O => \N__62858\,
            I => \N__62849\
        );

    \I__14292\ : InMux
    port map (
            O => \N__62855\,
            I => \N__62849\
        );

    \I__14291\ : InMux
    port map (
            O => \N__62854\,
            I => \N__62844\
        );

    \I__14290\ : LocalMux
    port map (
            O => \N__62849\,
            I => \N__62841\
        );

    \I__14289\ : InMux
    port map (
            O => \N__62848\,
            I => \N__62838\
        );

    \I__14288\ : CascadeMux
    port map (
            O => \N__62847\,
            I => \N__62835\
        );

    \I__14287\ : LocalMux
    port map (
            O => \N__62844\,
            I => \N__62832\
        );

    \I__14286\ : Span4Mux_v
    port map (
            O => \N__62841\,
            I => \N__62829\
        );

    \I__14285\ : LocalMux
    port map (
            O => \N__62838\,
            I => \N__62826\
        );

    \I__14284\ : InMux
    port map (
            O => \N__62835\,
            I => \N__62823\
        );

    \I__14283\ : Span12Mux_v
    port map (
            O => \N__62832\,
            I => \N__62820\
        );

    \I__14282\ : Span4Mux_v
    port map (
            O => \N__62829\,
            I => \N__62815\
        );

    \I__14281\ : Span4Mux_h
    port map (
            O => \N__62826\,
            I => \N__62815\
        );

    \I__14280\ : LocalMux
    port map (
            O => \N__62823\,
            I => \c0.data_in_frame_13_7\
        );

    \I__14279\ : Odrv12
    port map (
            O => \N__62820\,
            I => \c0.data_in_frame_13_7\
        );

    \I__14278\ : Odrv4
    port map (
            O => \N__62815\,
            I => \c0.data_in_frame_13_7\
        );

    \I__14277\ : InMux
    port map (
            O => \N__62808\,
            I => \N__62803\
        );

    \I__14276\ : CascadeMux
    port map (
            O => \N__62807\,
            I => \N__62800\
        );

    \I__14275\ : CascadeMux
    port map (
            O => \N__62806\,
            I => \N__62796\
        );

    \I__14274\ : LocalMux
    port map (
            O => \N__62803\,
            I => \N__62792\
        );

    \I__14273\ : InMux
    port map (
            O => \N__62800\,
            I => \N__62787\
        );

    \I__14272\ : InMux
    port map (
            O => \N__62799\,
            I => \N__62787\
        );

    \I__14271\ : InMux
    port map (
            O => \N__62796\,
            I => \N__62784\
        );

    \I__14270\ : InMux
    port map (
            O => \N__62795\,
            I => \N__62781\
        );

    \I__14269\ : Span4Mux_h
    port map (
            O => \N__62792\,
            I => \N__62774\
        );

    \I__14268\ : LocalMux
    port map (
            O => \N__62787\,
            I => \N__62774\
        );

    \I__14267\ : LocalMux
    port map (
            O => \N__62784\,
            I => \N__62774\
        );

    \I__14266\ : LocalMux
    port map (
            O => \N__62781\,
            I => \c0.data_in_frame_12_6\
        );

    \I__14265\ : Odrv4
    port map (
            O => \N__62774\,
            I => \c0.data_in_frame_12_6\
        );

    \I__14264\ : InMux
    port map (
            O => \N__62769\,
            I => \N__62759\
        );

    \I__14263\ : InMux
    port map (
            O => \N__62768\,
            I => \N__62759\
        );

    \I__14262\ : InMux
    port map (
            O => \N__62767\,
            I => \N__62759\
        );

    \I__14261\ : InMux
    port map (
            O => \N__62766\,
            I => \N__62753\
        );

    \I__14260\ : LocalMux
    port map (
            O => \N__62759\,
            I => \N__62750\
        );

    \I__14259\ : InMux
    port map (
            O => \N__62758\,
            I => \N__62743\
        );

    \I__14258\ : InMux
    port map (
            O => \N__62757\,
            I => \N__62743\
        );

    \I__14257\ : InMux
    port map (
            O => \N__62756\,
            I => \N__62743\
        );

    \I__14256\ : LocalMux
    port map (
            O => \N__62753\,
            I => \N__62735\
        );

    \I__14255\ : Span4Mux_v
    port map (
            O => \N__62750\,
            I => \N__62735\
        );

    \I__14254\ : LocalMux
    port map (
            O => \N__62743\,
            I => \N__62735\
        );

    \I__14253\ : InMux
    port map (
            O => \N__62742\,
            I => \N__62732\
        );

    \I__14252\ : Odrv4
    port map (
            O => \N__62735\,
            I => \c0.n22782\
        );

    \I__14251\ : LocalMux
    port map (
            O => \N__62732\,
            I => \c0.n22782\
        );

    \I__14250\ : InMux
    port map (
            O => \N__62727\,
            I => \N__62724\
        );

    \I__14249\ : LocalMux
    port map (
            O => \N__62724\,
            I => \c0.n12_adj_4246\
        );

    \I__14248\ : InMux
    port map (
            O => \N__62721\,
            I => \N__62715\
        );

    \I__14247\ : InMux
    port map (
            O => \N__62720\,
            I => \N__62715\
        );

    \I__14246\ : LocalMux
    port map (
            O => \N__62715\,
            I => \c0.n23453\
        );

    \I__14245\ : InMux
    port map (
            O => \N__62712\,
            I => \N__62705\
        );

    \I__14244\ : InMux
    port map (
            O => \N__62711\,
            I => \N__62705\
        );

    \I__14243\ : InMux
    port map (
            O => \N__62710\,
            I => \N__62702\
        );

    \I__14242\ : LocalMux
    port map (
            O => \N__62705\,
            I => \N__62699\
        );

    \I__14241\ : LocalMux
    port map (
            O => \N__62702\,
            I => \N__62696\
        );

    \I__14240\ : Span4Mux_h
    port map (
            O => \N__62699\,
            I => \N__62693\
        );

    \I__14239\ : Odrv4
    port map (
            O => \N__62696\,
            I => \c0.n22540\
        );

    \I__14238\ : Odrv4
    port map (
            O => \N__62693\,
            I => \c0.n22540\
        );

    \I__14237\ : InMux
    port map (
            O => \N__62688\,
            I => \N__62683\
        );

    \I__14236\ : InMux
    port map (
            O => \N__62687\,
            I => \N__62677\
        );

    \I__14235\ : InMux
    port map (
            O => \N__62686\,
            I => \N__62677\
        );

    \I__14234\ : LocalMux
    port map (
            O => \N__62683\,
            I => \N__62674\
        );

    \I__14233\ : InMux
    port map (
            O => \N__62682\,
            I => \N__62671\
        );

    \I__14232\ : LocalMux
    port map (
            O => \N__62677\,
            I => \N__62668\
        );

    \I__14231\ : Span4Mux_v
    port map (
            O => \N__62674\,
            I => \N__62663\
        );

    \I__14230\ : LocalMux
    port map (
            O => \N__62671\,
            I => \N__62658\
        );

    \I__14229\ : Span4Mux_h
    port map (
            O => \N__62668\,
            I => \N__62658\
        );

    \I__14228\ : InMux
    port map (
            O => \N__62667\,
            I => \N__62655\
        );

    \I__14227\ : InMux
    port map (
            O => \N__62666\,
            I => \N__62652\
        );

    \I__14226\ : Odrv4
    port map (
            O => \N__62663\,
            I => \c0.n24333\
        );

    \I__14225\ : Odrv4
    port map (
            O => \N__62658\,
            I => \c0.n24333\
        );

    \I__14224\ : LocalMux
    port map (
            O => \N__62655\,
            I => \c0.n24333\
        );

    \I__14223\ : LocalMux
    port map (
            O => \N__62652\,
            I => \c0.n24333\
        );

    \I__14222\ : CascadeMux
    port map (
            O => \N__62643\,
            I => \N__62640\
        );

    \I__14221\ : InMux
    port map (
            O => \N__62640\,
            I => \N__62635\
        );

    \I__14220\ : InMux
    port map (
            O => \N__62639\,
            I => \N__62632\
        );

    \I__14219\ : InMux
    port map (
            O => \N__62638\,
            I => \N__62629\
        );

    \I__14218\ : LocalMux
    port map (
            O => \N__62635\,
            I => \N__62624\
        );

    \I__14217\ : LocalMux
    port map (
            O => \N__62632\,
            I => \N__62624\
        );

    \I__14216\ : LocalMux
    port map (
            O => \N__62629\,
            I => \N__62621\
        );

    \I__14215\ : Odrv4
    port map (
            O => \N__62624\,
            I => \c0.n22822\
        );

    \I__14214\ : Odrv4
    port map (
            O => \N__62621\,
            I => \c0.n22822\
        );

    \I__14213\ : CascadeMux
    port map (
            O => \N__62616\,
            I => \N__62610\
        );

    \I__14212\ : CascadeMux
    port map (
            O => \N__62615\,
            I => \N__62607\
        );

    \I__14211\ : InMux
    port map (
            O => \N__62614\,
            I => \N__62604\
        );

    \I__14210\ : InMux
    port map (
            O => \N__62613\,
            I => \N__62598\
        );

    \I__14209\ : InMux
    port map (
            O => \N__62610\,
            I => \N__62598\
        );

    \I__14208\ : InMux
    port map (
            O => \N__62607\,
            I => \N__62595\
        );

    \I__14207\ : LocalMux
    port map (
            O => \N__62604\,
            I => \N__62592\
        );

    \I__14206\ : CascadeMux
    port map (
            O => \N__62603\,
            I => \N__62588\
        );

    \I__14205\ : LocalMux
    port map (
            O => \N__62598\,
            I => \N__62585\
        );

    \I__14204\ : LocalMux
    port map (
            O => \N__62595\,
            I => \N__62582\
        );

    \I__14203\ : Span4Mux_v
    port map (
            O => \N__62592\,
            I => \N__62579\
        );

    \I__14202\ : InMux
    port map (
            O => \N__62591\,
            I => \N__62574\
        );

    \I__14201\ : InMux
    port map (
            O => \N__62588\,
            I => \N__62574\
        );

    \I__14200\ : Span4Mux_v
    port map (
            O => \N__62585\,
            I => \N__62571\
        );

    \I__14199\ : Span4Mux_v
    port map (
            O => \N__62582\,
            I => \N__62566\
        );

    \I__14198\ : Span4Mux_h
    port map (
            O => \N__62579\,
            I => \N__62566\
        );

    \I__14197\ : LocalMux
    port map (
            O => \N__62574\,
            I => data_in_frame_14_7
        );

    \I__14196\ : Odrv4
    port map (
            O => \N__62571\,
            I => data_in_frame_14_7
        );

    \I__14195\ : Odrv4
    port map (
            O => \N__62566\,
            I => data_in_frame_14_7
        );

    \I__14194\ : CascadeMux
    port map (
            O => \N__62559\,
            I => \c0.n12_adj_4246_cascade_\
        );

    \I__14193\ : CascadeMux
    port map (
            O => \N__62556\,
            I => \c0.n23691_cascade_\
        );

    \I__14192\ : InMux
    port map (
            O => \N__62553\,
            I => \N__62550\
        );

    \I__14191\ : LocalMux
    port map (
            O => \N__62550\,
            I => \N__62546\
        );

    \I__14190\ : InMux
    port map (
            O => \N__62549\,
            I => \N__62543\
        );

    \I__14189\ : Span4Mux_v
    port map (
            O => \N__62546\,
            I => \N__62538\
        );

    \I__14188\ : LocalMux
    port map (
            O => \N__62543\,
            I => \N__62538\
        );

    \I__14187\ : Span4Mux_h
    port map (
            O => \N__62538\,
            I => \N__62535\
        );

    \I__14186\ : Odrv4
    port map (
            O => \N__62535\,
            I => \c0.n20543\
        );

    \I__14185\ : InMux
    port map (
            O => \N__62532\,
            I => \N__62529\
        );

    \I__14184\ : LocalMux
    port map (
            O => \N__62529\,
            I => \N__62523\
        );

    \I__14183\ : InMux
    port map (
            O => \N__62528\,
            I => \N__62518\
        );

    \I__14182\ : InMux
    port map (
            O => \N__62527\,
            I => \N__62518\
        );

    \I__14181\ : CascadeMux
    port map (
            O => \N__62526\,
            I => \N__62515\
        );

    \I__14180\ : Span4Mux_h
    port map (
            O => \N__62523\,
            I => \N__62512\
        );

    \I__14179\ : LocalMux
    port map (
            O => \N__62518\,
            I => \N__62509\
        );

    \I__14178\ : InMux
    port map (
            O => \N__62515\,
            I => \N__62506\
        );

    \I__14177\ : Span4Mux_h
    port map (
            O => \N__62512\,
            I => \N__62503\
        );

    \I__14176\ : Span4Mux_v
    port map (
            O => \N__62509\,
            I => \N__62500\
        );

    \I__14175\ : LocalMux
    port map (
            O => \N__62506\,
            I => \c0.data_in_frame_16_5\
        );

    \I__14174\ : Odrv4
    port map (
            O => \N__62503\,
            I => \c0.data_in_frame_16_5\
        );

    \I__14173\ : Odrv4
    port map (
            O => \N__62500\,
            I => \c0.data_in_frame_16_5\
        );

    \I__14172\ : InMux
    port map (
            O => \N__62493\,
            I => \N__62490\
        );

    \I__14171\ : LocalMux
    port map (
            O => \N__62490\,
            I => \c0.n10_adj_4602\
        );

    \I__14170\ : InMux
    port map (
            O => \N__62487\,
            I => \N__62484\
        );

    \I__14169\ : LocalMux
    port map (
            O => \N__62484\,
            I => \N__62480\
        );

    \I__14168\ : InMux
    port map (
            O => \N__62483\,
            I => \N__62477\
        );

    \I__14167\ : Span4Mux_h
    port map (
            O => \N__62480\,
            I => \N__62471\
        );

    \I__14166\ : LocalMux
    port map (
            O => \N__62477\,
            I => \N__62471\
        );

    \I__14165\ : InMux
    port map (
            O => \N__62476\,
            I => \N__62468\
        );

    \I__14164\ : Odrv4
    port map (
            O => \N__62471\,
            I => \c0.n22644\
        );

    \I__14163\ : LocalMux
    port map (
            O => \N__62468\,
            I => \c0.n22644\
        );

    \I__14162\ : InMux
    port map (
            O => \N__62463\,
            I => \N__62460\
        );

    \I__14161\ : LocalMux
    port map (
            O => \N__62460\,
            I => \N__62455\
        );

    \I__14160\ : CascadeMux
    port map (
            O => \N__62459\,
            I => \N__62452\
        );

    \I__14159\ : InMux
    port map (
            O => \N__62458\,
            I => \N__62449\
        );

    \I__14158\ : Span4Mux_h
    port map (
            O => \N__62455\,
            I => \N__62446\
        );

    \I__14157\ : InMux
    port map (
            O => \N__62452\,
            I => \N__62442\
        );

    \I__14156\ : LocalMux
    port map (
            O => \N__62449\,
            I => \N__62439\
        );

    \I__14155\ : Span4Mux_h
    port map (
            O => \N__62446\,
            I => \N__62436\
        );

    \I__14154\ : InMux
    port map (
            O => \N__62445\,
            I => \N__62433\
        );

    \I__14153\ : LocalMux
    port map (
            O => \N__62442\,
            I => \c0.data_in_frame_15_1\
        );

    \I__14152\ : Odrv4
    port map (
            O => \N__62439\,
            I => \c0.data_in_frame_15_1\
        );

    \I__14151\ : Odrv4
    port map (
            O => \N__62436\,
            I => \c0.data_in_frame_15_1\
        );

    \I__14150\ : LocalMux
    port map (
            O => \N__62433\,
            I => \c0.data_in_frame_15_1\
        );

    \I__14149\ : InMux
    port map (
            O => \N__62424\,
            I => \N__62420\
        );

    \I__14148\ : InMux
    port map (
            O => \N__62423\,
            I => \N__62417\
        );

    \I__14147\ : LocalMux
    port map (
            O => \N__62420\,
            I => \c0.n14165\
        );

    \I__14146\ : LocalMux
    port map (
            O => \N__62417\,
            I => \c0.n14165\
        );

    \I__14145\ : CascadeMux
    port map (
            O => \N__62412\,
            I => \N__62408\
        );

    \I__14144\ : InMux
    port map (
            O => \N__62411\,
            I => \N__62404\
        );

    \I__14143\ : InMux
    port map (
            O => \N__62408\,
            I => \N__62401\
        );

    \I__14142\ : InMux
    port map (
            O => \N__62407\,
            I => \N__62398\
        );

    \I__14141\ : LocalMux
    port map (
            O => \N__62404\,
            I => \N__62389\
        );

    \I__14140\ : LocalMux
    port map (
            O => \N__62401\,
            I => \N__62389\
        );

    \I__14139\ : LocalMux
    port map (
            O => \N__62398\,
            I => \N__62389\
        );

    \I__14138\ : InMux
    port map (
            O => \N__62397\,
            I => \N__62386\
        );

    \I__14137\ : InMux
    port map (
            O => \N__62396\,
            I => \N__62383\
        );

    \I__14136\ : Span4Mux_v
    port map (
            O => \N__62389\,
            I => \N__62380\
        );

    \I__14135\ : LocalMux
    port map (
            O => \N__62386\,
            I => \N__62376\
        );

    \I__14134\ : LocalMux
    port map (
            O => \N__62383\,
            I => \N__62371\
        );

    \I__14133\ : Span4Mux_h
    port map (
            O => \N__62380\,
            I => \N__62371\
        );

    \I__14132\ : InMux
    port map (
            O => \N__62379\,
            I => \N__62368\
        );

    \I__14131\ : Odrv4
    port map (
            O => \N__62376\,
            I => data_in_frame_14_5
        );

    \I__14130\ : Odrv4
    port map (
            O => \N__62371\,
            I => data_in_frame_14_5
        );

    \I__14129\ : LocalMux
    port map (
            O => \N__62368\,
            I => data_in_frame_14_5
        );

    \I__14128\ : CascadeMux
    port map (
            O => \N__62361\,
            I => \N__62357\
        );

    \I__14127\ : InMux
    port map (
            O => \N__62360\,
            I => \N__62350\
        );

    \I__14126\ : InMux
    port map (
            O => \N__62357\,
            I => \N__62345\
        );

    \I__14125\ : InMux
    port map (
            O => \N__62356\,
            I => \N__62345\
        );

    \I__14124\ : InMux
    port map (
            O => \N__62355\,
            I => \N__62338\
        );

    \I__14123\ : InMux
    port map (
            O => \N__62354\,
            I => \N__62338\
        );

    \I__14122\ : InMux
    port map (
            O => \N__62353\,
            I => \N__62338\
        );

    \I__14121\ : LocalMux
    port map (
            O => \N__62350\,
            I => \c0.n24444\
        );

    \I__14120\ : LocalMux
    port map (
            O => \N__62345\,
            I => \c0.n24444\
        );

    \I__14119\ : LocalMux
    port map (
            O => \N__62338\,
            I => \c0.n24444\
        );

    \I__14118\ : CascadeMux
    port map (
            O => \N__62331\,
            I => \N__62328\
        );

    \I__14117\ : InMux
    port map (
            O => \N__62328\,
            I => \N__62325\
        );

    \I__14116\ : LocalMux
    port map (
            O => \N__62325\,
            I => \N__62322\
        );

    \I__14115\ : Odrv4
    port map (
            O => \N__62322\,
            I => \c0.n7_adj_4581\
        );

    \I__14114\ : InMux
    port map (
            O => \N__62319\,
            I => \N__62313\
        );

    \I__14113\ : InMux
    port map (
            O => \N__62318\,
            I => \N__62310\
        );

    \I__14112\ : InMux
    port map (
            O => \N__62317\,
            I => \N__62306\
        );

    \I__14111\ : InMux
    port map (
            O => \N__62316\,
            I => \N__62303\
        );

    \I__14110\ : LocalMux
    port map (
            O => \N__62313\,
            I => \N__62300\
        );

    \I__14109\ : LocalMux
    port map (
            O => \N__62310\,
            I => \N__62297\
        );

    \I__14108\ : InMux
    port map (
            O => \N__62309\,
            I => \N__62291\
        );

    \I__14107\ : LocalMux
    port map (
            O => \N__62306\,
            I => \N__62286\
        );

    \I__14106\ : LocalMux
    port map (
            O => \N__62303\,
            I => \N__62286\
        );

    \I__14105\ : Span4Mux_h
    port map (
            O => \N__62300\,
            I => \N__62281\
        );

    \I__14104\ : Span4Mux_v
    port map (
            O => \N__62297\,
            I => \N__62281\
        );

    \I__14103\ : InMux
    port map (
            O => \N__62296\,
            I => \N__62278\
        );

    \I__14102\ : InMux
    port map (
            O => \N__62295\,
            I => \N__62275\
        );

    \I__14101\ : InMux
    port map (
            O => \N__62294\,
            I => \N__62272\
        );

    \I__14100\ : LocalMux
    port map (
            O => \N__62291\,
            I => \N__62268\
        );

    \I__14099\ : Span4Mux_v
    port map (
            O => \N__62286\,
            I => \N__62265\
        );

    \I__14098\ : Span4Mux_v
    port map (
            O => \N__62281\,
            I => \N__62262\
        );

    \I__14097\ : LocalMux
    port map (
            O => \N__62278\,
            I => \N__62259\
        );

    \I__14096\ : LocalMux
    port map (
            O => \N__62275\,
            I => \N__62254\
        );

    \I__14095\ : LocalMux
    port map (
            O => \N__62272\,
            I => \N__62254\
        );

    \I__14094\ : InMux
    port map (
            O => \N__62271\,
            I => \N__62250\
        );

    \I__14093\ : Span4Mux_h
    port map (
            O => \N__62268\,
            I => \N__62245\
        );

    \I__14092\ : Span4Mux_v
    port map (
            O => \N__62265\,
            I => \N__62245\
        );

    \I__14091\ : Span4Mux_v
    port map (
            O => \N__62262\,
            I => \N__62241\
        );

    \I__14090\ : Span4Mux_h
    port map (
            O => \N__62259\,
            I => \N__62236\
        );

    \I__14089\ : Span4Mux_h
    port map (
            O => \N__62254\,
            I => \N__62236\
        );

    \I__14088\ : InMux
    port map (
            O => \N__62253\,
            I => \N__62233\
        );

    \I__14087\ : LocalMux
    port map (
            O => \N__62250\,
            I => \N__62228\
        );

    \I__14086\ : Span4Mux_h
    port map (
            O => \N__62245\,
            I => \N__62228\
        );

    \I__14085\ : InMux
    port map (
            O => \N__62244\,
            I => \N__62225\
        );

    \I__14084\ : Span4Mux_v
    port map (
            O => \N__62241\,
            I => \N__62222\
        );

    \I__14083\ : Span4Mux_v
    port map (
            O => \N__62236\,
            I => \N__62219\
        );

    \I__14082\ : LocalMux
    port map (
            O => \N__62233\,
            I => \N__62216\
        );

    \I__14081\ : Span4Mux_v
    port map (
            O => \N__62228\,
            I => \N__62213\
        );

    \I__14080\ : LocalMux
    port map (
            O => \N__62225\,
            I => \N__62210\
        );

    \I__14079\ : Span4Mux_v
    port map (
            O => \N__62222\,
            I => \N__62207\
        );

    \I__14078\ : Span4Mux_v
    port map (
            O => \N__62219\,
            I => \N__62204\
        );

    \I__14077\ : Span12Mux_v
    port map (
            O => \N__62216\,
            I => \N__62201\
        );

    \I__14076\ : Span4Mux_v
    port map (
            O => \N__62213\,
            I => \N__62198\
        );

    \I__14075\ : Span12Mux_h
    port map (
            O => \N__62210\,
            I => \N__62194\
        );

    \I__14074\ : Span4Mux_h
    port map (
            O => \N__62207\,
            I => \N__62191\
        );

    \I__14073\ : Span4Mux_v
    port map (
            O => \N__62204\,
            I => \N__62188\
        );

    \I__14072\ : Span12Mux_v
    port map (
            O => \N__62201\,
            I => \N__62185\
        );

    \I__14071\ : Span4Mux_v
    port map (
            O => \N__62198\,
            I => \N__62182\
        );

    \I__14070\ : InMux
    port map (
            O => \N__62197\,
            I => \N__62179\
        );

    \I__14069\ : Odrv12
    port map (
            O => \N__62194\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__14068\ : Odrv4
    port map (
            O => \N__62191\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__14067\ : Odrv4
    port map (
            O => \N__62188\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__14066\ : Odrv12
    port map (
            O => \N__62185\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__14065\ : Odrv4
    port map (
            O => \N__62182\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__14064\ : LocalMux
    port map (
            O => \N__62179\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__14063\ : SRMux
    port map (
            O => \N__62166\,
            I => \N__62163\
        );

    \I__14062\ : LocalMux
    port map (
            O => \N__62163\,
            I => \N__62160\
        );

    \I__14061\ : Span12Mux_s5_v
    port map (
            O => \N__62160\,
            I => \N__62157\
        );

    \I__14060\ : Span12Mux_v
    port map (
            O => \N__62157\,
            I => \N__62154\
        );

    \I__14059\ : Odrv12
    port map (
            O => \N__62154\,
            I => \c0.n3_adj_4430\
        );

    \I__14058\ : InMux
    port map (
            O => \N__62151\,
            I => \N__62148\
        );

    \I__14057\ : LocalMux
    port map (
            O => \N__62148\,
            I => \N__62145\
        );

    \I__14056\ : Odrv12
    port map (
            O => \N__62145\,
            I => \c0.n124\
        );

    \I__14055\ : InMux
    port map (
            O => \N__62142\,
            I => \N__62136\
        );

    \I__14054\ : InMux
    port map (
            O => \N__62141\,
            I => \N__62136\
        );

    \I__14053\ : LocalMux
    port map (
            O => \N__62136\,
            I => \c0.n10_adj_4247\
        );

    \I__14052\ : InMux
    port map (
            O => \N__62133\,
            I => \N__62127\
        );

    \I__14051\ : InMux
    port map (
            O => \N__62132\,
            I => \N__62127\
        );

    \I__14050\ : LocalMux
    port map (
            O => \N__62127\,
            I => \c0.n22547\
        );

    \I__14049\ : InMux
    port map (
            O => \N__62124\,
            I => \N__62120\
        );

    \I__14048\ : InMux
    port map (
            O => \N__62123\,
            I => \N__62116\
        );

    \I__14047\ : LocalMux
    port map (
            O => \N__62120\,
            I => \N__62113\
        );

    \I__14046\ : InMux
    port map (
            O => \N__62119\,
            I => \N__62110\
        );

    \I__14045\ : LocalMux
    port map (
            O => \N__62116\,
            I => \N__62107\
        );

    \I__14044\ : Span4Mux_v
    port map (
            O => \N__62113\,
            I => \N__62102\
        );

    \I__14043\ : LocalMux
    port map (
            O => \N__62110\,
            I => \N__62102\
        );

    \I__14042\ : Span4Mux_v
    port map (
            O => \N__62107\,
            I => \N__62099\
        );

    \I__14041\ : Span4Mux_v
    port map (
            O => \N__62102\,
            I => \N__62096\
        );

    \I__14040\ : Odrv4
    port map (
            O => \N__62099\,
            I => \c0.n13998\
        );

    \I__14039\ : Odrv4
    port map (
            O => \N__62096\,
            I => \c0.n13998\
        );

    \I__14038\ : InMux
    port map (
            O => \N__62091\,
            I => \N__62088\
        );

    \I__14037\ : LocalMux
    port map (
            O => \N__62088\,
            I => \N__62085\
        );

    \I__14036\ : Span4Mux_v
    port map (
            O => \N__62085\,
            I => \N__62081\
        );

    \I__14035\ : InMux
    port map (
            O => \N__62084\,
            I => \N__62078\
        );

    \I__14034\ : Span4Mux_v
    port map (
            O => \N__62081\,
            I => \N__62075\
        );

    \I__14033\ : LocalMux
    port map (
            O => \N__62078\,
            I => \N__62072\
        );

    \I__14032\ : Span4Mux_h
    port map (
            O => \N__62075\,
            I => \N__62064\
        );

    \I__14031\ : Span4Mux_v
    port map (
            O => \N__62072\,
            I => \N__62064\
        );

    \I__14030\ : InMux
    port map (
            O => \N__62071\,
            I => \N__62057\
        );

    \I__14029\ : InMux
    port map (
            O => \N__62070\,
            I => \N__62057\
        );

    \I__14028\ : InMux
    port map (
            O => \N__62069\,
            I => \N__62057\
        );

    \I__14027\ : Odrv4
    port map (
            O => \N__62064\,
            I => \c0.n23156\
        );

    \I__14026\ : LocalMux
    port map (
            O => \N__62057\,
            I => \c0.n23156\
        );

    \I__14025\ : InMux
    port map (
            O => \N__62052\,
            I => \N__62049\
        );

    \I__14024\ : LocalMux
    port map (
            O => \N__62049\,
            I => \N__62046\
        );

    \I__14023\ : Span4Mux_v
    port map (
            O => \N__62046\,
            I => \N__62043\
        );

    \I__14022\ : Span4Mux_h
    port map (
            O => \N__62043\,
            I => \N__62040\
        );

    \I__14021\ : Odrv4
    port map (
            O => \N__62040\,
            I => \c0.n65\
        );

    \I__14020\ : InMux
    port map (
            O => \N__62037\,
            I => \N__62034\
        );

    \I__14019\ : LocalMux
    port map (
            O => \N__62034\,
            I => \N__62030\
        );

    \I__14018\ : InMux
    port map (
            O => \N__62033\,
            I => \N__62027\
        );

    \I__14017\ : Odrv12
    port map (
            O => \N__62030\,
            I => \c0.n60\
        );

    \I__14016\ : LocalMux
    port map (
            O => \N__62027\,
            I => \c0.n60\
        );

    \I__14015\ : CascadeMux
    port map (
            O => \N__62022\,
            I => \c0.n59_cascade_\
        );

    \I__14014\ : InMux
    port map (
            O => \N__62019\,
            I => \N__62016\
        );

    \I__14013\ : LocalMux
    port map (
            O => \N__62016\,
            I => \c0.n70\
        );

    \I__14012\ : CascadeMux
    port map (
            O => \N__62013\,
            I => \c0.n24444_cascade_\
        );

    \I__14011\ : InMux
    port map (
            O => \N__62010\,
            I => \N__62006\
        );

    \I__14010\ : InMux
    port map (
            O => \N__62009\,
            I => \N__62003\
        );

    \I__14009\ : LocalMux
    port map (
            O => \N__62006\,
            I => \N__62000\
        );

    \I__14008\ : LocalMux
    port map (
            O => \N__62003\,
            I => \c0.n21282\
        );

    \I__14007\ : Odrv4
    port map (
            O => \N__62000\,
            I => \c0.n21282\
        );

    \I__14006\ : InMux
    port map (
            O => \N__61995\,
            I => \N__61992\
        );

    \I__14005\ : LocalMux
    port map (
            O => \N__61992\,
            I => \N__61988\
        );

    \I__14004\ : CascadeMux
    port map (
            O => \N__61991\,
            I => \N__61984\
        );

    \I__14003\ : Span4Mux_h
    port map (
            O => \N__61988\,
            I => \N__61981\
        );

    \I__14002\ : CascadeMux
    port map (
            O => \N__61987\,
            I => \N__61978\
        );

    \I__14001\ : InMux
    port map (
            O => \N__61984\,
            I => \N__61975\
        );

    \I__14000\ : Span4Mux_v
    port map (
            O => \N__61981\,
            I => \N__61972\
        );

    \I__13999\ : InMux
    port map (
            O => \N__61978\,
            I => \N__61969\
        );

    \I__13998\ : LocalMux
    port map (
            O => \N__61975\,
            I => \c0.data_in_frame_15_7\
        );

    \I__13997\ : Odrv4
    port map (
            O => \N__61972\,
            I => \c0.data_in_frame_15_7\
        );

    \I__13996\ : LocalMux
    port map (
            O => \N__61969\,
            I => \c0.data_in_frame_15_7\
        );

    \I__13995\ : CascadeMux
    port map (
            O => \N__61962\,
            I => \N__61959\
        );

    \I__13994\ : InMux
    port map (
            O => \N__61959\,
            I => \N__61956\
        );

    \I__13993\ : LocalMux
    port map (
            O => \N__61956\,
            I => \N__61953\
        );

    \I__13992\ : Span4Mux_h
    port map (
            O => \N__61953\,
            I => \N__61950\
        );

    \I__13991\ : Span4Mux_h
    port map (
            O => \N__61950\,
            I => \N__61946\
        );

    \I__13990\ : InMux
    port map (
            O => \N__61949\,
            I => \N__61943\
        );

    \I__13989\ : Odrv4
    port map (
            O => \N__61946\,
            I => \c0.n22514\
        );

    \I__13988\ : LocalMux
    port map (
            O => \N__61943\,
            I => \c0.n22514\
        );

    \I__13987\ : CascadeMux
    port map (
            O => \N__61938\,
            I => \c0.n23224_cascade_\
        );

    \I__13986\ : InMux
    port map (
            O => \N__61935\,
            I => \N__61931\
        );

    \I__13985\ : InMux
    port map (
            O => \N__61934\,
            I => \N__61928\
        );

    \I__13984\ : LocalMux
    port map (
            O => \N__61931\,
            I => \N__61921\
        );

    \I__13983\ : LocalMux
    port map (
            O => \N__61928\,
            I => \N__61921\
        );

    \I__13982\ : InMux
    port map (
            O => \N__61927\,
            I => \N__61916\
        );

    \I__13981\ : InMux
    port map (
            O => \N__61926\,
            I => \N__61916\
        );

    \I__13980\ : Span4Mux_v
    port map (
            O => \N__61921\,
            I => \N__61913\
        );

    \I__13979\ : LocalMux
    port map (
            O => \N__61916\,
            I => \N__61910\
        );

    \I__13978\ : Span4Mux_h
    port map (
            O => \N__61913\,
            I => \N__61905\
        );

    \I__13977\ : Span4Mux_v
    port map (
            O => \N__61910\,
            I => \N__61905\
        );

    \I__13976\ : Odrv4
    port map (
            O => \N__61905\,
            I => \c0.n21409\
        );

    \I__13975\ : InMux
    port map (
            O => \N__61902\,
            I => \N__61898\
        );

    \I__13974\ : InMux
    port map (
            O => \N__61901\,
            I => \N__61894\
        );

    \I__13973\ : LocalMux
    port map (
            O => \N__61898\,
            I => \N__61891\
        );

    \I__13972\ : CascadeMux
    port map (
            O => \N__61897\,
            I => \N__61887\
        );

    \I__13971\ : LocalMux
    port map (
            O => \N__61894\,
            I => \N__61884\
        );

    \I__13970\ : Span4Mux_v
    port map (
            O => \N__61891\,
            I => \N__61881\
        );

    \I__13969\ : InMux
    port map (
            O => \N__61890\,
            I => \N__61878\
        );

    \I__13968\ : InMux
    port map (
            O => \N__61887\,
            I => \N__61875\
        );

    \I__13967\ : Span4Mux_h
    port map (
            O => \N__61884\,
            I => \N__61872\
        );

    \I__13966\ : Sp12to4
    port map (
            O => \N__61881\,
            I => \N__61867\
        );

    \I__13965\ : LocalMux
    port map (
            O => \N__61878\,
            I => \N__61867\
        );

    \I__13964\ : LocalMux
    port map (
            O => \N__61875\,
            I => \c0.data_in_frame_18_6\
        );

    \I__13963\ : Odrv4
    port map (
            O => \N__61872\,
            I => \c0.data_in_frame_18_6\
        );

    \I__13962\ : Odrv12
    port map (
            O => \N__61867\,
            I => \c0.data_in_frame_18_6\
        );

    \I__13961\ : InMux
    port map (
            O => \N__61860\,
            I => \N__61856\
        );

    \I__13960\ : InMux
    port map (
            O => \N__61859\,
            I => \N__61853\
        );

    \I__13959\ : LocalMux
    port map (
            O => \N__61856\,
            I => \N__61846\
        );

    \I__13958\ : LocalMux
    port map (
            O => \N__61853\,
            I => \N__61846\
        );

    \I__13957\ : InMux
    port map (
            O => \N__61852\,
            I => \N__61841\
        );

    \I__13956\ : InMux
    port map (
            O => \N__61851\,
            I => \N__61841\
        );

    \I__13955\ : Span4Mux_h
    port map (
            O => \N__61846\,
            I => \N__61838\
        );

    \I__13954\ : LocalMux
    port map (
            O => \N__61841\,
            I => \c0.n13128\
        );

    \I__13953\ : Odrv4
    port map (
            O => \N__61838\,
            I => \c0.n13128\
        );

    \I__13952\ : CascadeMux
    port map (
            O => \N__61833\,
            I => \N__61830\
        );

    \I__13951\ : InMux
    port map (
            O => \N__61830\,
            I => \N__61827\
        );

    \I__13950\ : LocalMux
    port map (
            O => \N__61827\,
            I => \N__61824\
        );

    \I__13949\ : Span4Mux_v
    port map (
            O => \N__61824\,
            I => \N__61821\
        );

    \I__13948\ : Span4Mux_v
    port map (
            O => \N__61821\,
            I => \N__61818\
        );

    \I__13947\ : Odrv4
    port map (
            O => \N__61818\,
            I => \c0.n7_adj_4603\
        );

    \I__13946\ : InMux
    port map (
            O => \N__61815\,
            I => \N__61812\
        );

    \I__13945\ : LocalMux
    port map (
            O => \N__61812\,
            I => \N__61808\
        );

    \I__13944\ : InMux
    port map (
            O => \N__61811\,
            I => \N__61805\
        );

    \I__13943\ : Odrv4
    port map (
            O => \N__61808\,
            I => \c0.n22589\
        );

    \I__13942\ : LocalMux
    port map (
            O => \N__61805\,
            I => \c0.n22589\
        );

    \I__13941\ : CascadeMux
    port map (
            O => \N__61800\,
            I => \c0.n13738_cascade_\
        );

    \I__13940\ : InMux
    port map (
            O => \N__61797\,
            I => \N__61793\
        );

    \I__13939\ : InMux
    port map (
            O => \N__61796\,
            I => \N__61789\
        );

    \I__13938\ : LocalMux
    port map (
            O => \N__61793\,
            I => \N__61786\
        );

    \I__13937\ : InMux
    port map (
            O => \N__61792\,
            I => \N__61783\
        );

    \I__13936\ : LocalMux
    port map (
            O => \N__61789\,
            I => \N__61774\
        );

    \I__13935\ : Span4Mux_v
    port map (
            O => \N__61786\,
            I => \N__61774\
        );

    \I__13934\ : LocalMux
    port map (
            O => \N__61783\,
            I => \N__61774\
        );

    \I__13933\ : InMux
    port map (
            O => \N__61782\,
            I => \N__61771\
        );

    \I__13932\ : CascadeMux
    port map (
            O => \N__61781\,
            I => \N__61768\
        );

    \I__13931\ : Span4Mux_v
    port map (
            O => \N__61774\,
            I => \N__61762\
        );

    \I__13930\ : LocalMux
    port map (
            O => \N__61771\,
            I => \N__61762\
        );

    \I__13929\ : InMux
    port map (
            O => \N__61768\,
            I => \N__61759\
        );

    \I__13928\ : InMux
    port map (
            O => \N__61767\,
            I => \N__61756\
        );

    \I__13927\ : Span4Mux_v
    port map (
            O => \N__61762\,
            I => \N__61753\
        );

    \I__13926\ : LocalMux
    port map (
            O => \N__61759\,
            I => \c0.data_in_frame_10_6\
        );

    \I__13925\ : LocalMux
    port map (
            O => \N__61756\,
            I => \c0.data_in_frame_10_6\
        );

    \I__13924\ : Odrv4
    port map (
            O => \N__61753\,
            I => \c0.data_in_frame_10_6\
        );

    \I__13923\ : InMux
    port map (
            O => \N__61746\,
            I => \N__61742\
        );

    \I__13922\ : CascadeMux
    port map (
            O => \N__61745\,
            I => \N__61735\
        );

    \I__13921\ : LocalMux
    port map (
            O => \N__61742\,
            I => \N__61732\
        );

    \I__13920\ : InMux
    port map (
            O => \N__61741\,
            I => \N__61725\
        );

    \I__13919\ : InMux
    port map (
            O => \N__61740\,
            I => \N__61725\
        );

    \I__13918\ : InMux
    port map (
            O => \N__61739\,
            I => \N__61725\
        );

    \I__13917\ : InMux
    port map (
            O => \N__61738\,
            I => \N__61720\
        );

    \I__13916\ : InMux
    port map (
            O => \N__61735\,
            I => \N__61720\
        );

    \I__13915\ : Span4Mux_v
    port map (
            O => \N__61732\,
            I => \N__61716\
        );

    \I__13914\ : LocalMux
    port map (
            O => \N__61725\,
            I => \N__61711\
        );

    \I__13913\ : LocalMux
    port map (
            O => \N__61720\,
            I => \N__61711\
        );

    \I__13912\ : InMux
    port map (
            O => \N__61719\,
            I => \N__61708\
        );

    \I__13911\ : Sp12to4
    port map (
            O => \N__61716\,
            I => \N__61703\
        );

    \I__13910\ : Span12Mux_v
    port map (
            O => \N__61711\,
            I => \N__61703\
        );

    \I__13909\ : LocalMux
    port map (
            O => \N__61708\,
            I => \c0.data_in_frame_10_7\
        );

    \I__13908\ : Odrv12
    port map (
            O => \N__61703\,
            I => \c0.data_in_frame_10_7\
        );

    \I__13907\ : InMux
    port map (
            O => \N__61698\,
            I => \N__61695\
        );

    \I__13906\ : LocalMux
    port map (
            O => \N__61695\,
            I => \N__61692\
        );

    \I__13905\ : Span4Mux_h
    port map (
            O => \N__61692\,
            I => \N__61688\
        );

    \I__13904\ : InMux
    port map (
            O => \N__61691\,
            I => \N__61685\
        );

    \I__13903\ : Odrv4
    port map (
            O => \N__61688\,
            I => \c0.n13734\
        );

    \I__13902\ : LocalMux
    port map (
            O => \N__61685\,
            I => \c0.n13734\
        );

    \I__13901\ : CascadeMux
    port map (
            O => \N__61680\,
            I => \c0.n39_adj_4708_cascade_\
        );

    \I__13900\ : InMux
    port map (
            O => \N__61677\,
            I => \N__61674\
        );

    \I__13899\ : LocalMux
    port map (
            O => \N__61674\,
            I => \N__61671\
        );

    \I__13898\ : Span4Mux_h
    port map (
            O => \N__61671\,
            I => \N__61668\
        );

    \I__13897\ : Span4Mux_v
    port map (
            O => \N__61668\,
            I => \N__61665\
        );

    \I__13896\ : Odrv4
    port map (
            O => \N__61665\,
            I => \c0.n63\
        );

    \I__13895\ : CascadeMux
    port map (
            O => \N__61662\,
            I => \c0.n64_cascade_\
        );

    \I__13894\ : CascadeMux
    port map (
            O => \N__61659\,
            I => \N__61655\
        );

    \I__13893\ : InMux
    port map (
            O => \N__61658\,
            I => \N__61652\
        );

    \I__13892\ : InMux
    port map (
            O => \N__61655\,
            I => \N__61649\
        );

    \I__13891\ : LocalMux
    port map (
            O => \N__61652\,
            I => \N__61645\
        );

    \I__13890\ : LocalMux
    port map (
            O => \N__61649\,
            I => \N__61642\
        );

    \I__13889\ : InMux
    port map (
            O => \N__61648\,
            I => \N__61639\
        );

    \I__13888\ : Span4Mux_h
    port map (
            O => \N__61645\,
            I => \N__61634\
        );

    \I__13887\ : Span4Mux_h
    port map (
            O => \N__61642\,
            I => \N__61634\
        );

    \I__13886\ : LocalMux
    port map (
            O => \N__61639\,
            I => \c0.n13721\
        );

    \I__13885\ : Odrv4
    port map (
            O => \N__61634\,
            I => \c0.n13721\
        );

    \I__13884\ : InMux
    port map (
            O => \N__61629\,
            I => \N__61626\
        );

    \I__13883\ : LocalMux
    port map (
            O => \N__61626\,
            I => \c0.n55_adj_4709\
        );

    \I__13882\ : CascadeMux
    port map (
            O => \N__61623\,
            I => \N__61620\
        );

    \I__13881\ : InMux
    port map (
            O => \N__61620\,
            I => \N__61617\
        );

    \I__13880\ : LocalMux
    port map (
            O => \N__61617\,
            I => \N__61613\
        );

    \I__13879\ : InMux
    port map (
            O => \N__61616\,
            I => \N__61610\
        );

    \I__13878\ : Span4Mux_v
    port map (
            O => \N__61613\,
            I => \N__61607\
        );

    \I__13877\ : LocalMux
    port map (
            O => \N__61610\,
            I => \N__61604\
        );

    \I__13876\ : Span4Mux_h
    port map (
            O => \N__61607\,
            I => \N__61601\
        );

    \I__13875\ : Odrv4
    port map (
            O => \N__61604\,
            I => \c0.n13186\
        );

    \I__13874\ : Odrv4
    port map (
            O => \N__61601\,
            I => \c0.n13186\
        );

    \I__13873\ : CascadeMux
    port map (
            O => \N__61596\,
            I => \N__61593\
        );

    \I__13872\ : InMux
    port map (
            O => \N__61593\,
            I => \N__61590\
        );

    \I__13871\ : LocalMux
    port map (
            O => \N__61590\,
            I => \N__61586\
        );

    \I__13870\ : InMux
    port map (
            O => \N__61589\,
            I => \N__61583\
        );

    \I__13869\ : Span4Mux_v
    port map (
            O => \N__61586\,
            I => \N__61579\
        );

    \I__13868\ : LocalMux
    port map (
            O => \N__61583\,
            I => \N__61576\
        );

    \I__13867\ : InMux
    port map (
            O => \N__61582\,
            I => \N__61573\
        );

    \I__13866\ : Span4Mux_h
    port map (
            O => \N__61579\,
            I => \N__61570\
        );

    \I__13865\ : Span12Mux_h
    port map (
            O => \N__61576\,
            I => \N__61567\
        );

    \I__13864\ : LocalMux
    port map (
            O => \N__61573\,
            I => \c0.data_in_frame_10_5\
        );

    \I__13863\ : Odrv4
    port map (
            O => \N__61570\,
            I => \c0.data_in_frame_10_5\
        );

    \I__13862\ : Odrv12
    port map (
            O => \N__61567\,
            I => \c0.data_in_frame_10_5\
        );

    \I__13861\ : CascadeMux
    port map (
            O => \N__61560\,
            I => \c0.n96_cascade_\
        );

    \I__13860\ : InMux
    port map (
            O => \N__61557\,
            I => \N__61554\
        );

    \I__13859\ : LocalMux
    port map (
            O => \N__61554\,
            I => \N__61549\
        );

    \I__13858\ : InMux
    port map (
            O => \N__61553\,
            I => \N__61545\
        );

    \I__13857\ : InMux
    port map (
            O => \N__61552\,
            I => \N__61542\
        );

    \I__13856\ : Span4Mux_h
    port map (
            O => \N__61549\,
            I => \N__61538\
        );

    \I__13855\ : CascadeMux
    port map (
            O => \N__61548\,
            I => \N__61535\
        );

    \I__13854\ : LocalMux
    port map (
            O => \N__61545\,
            I => \N__61530\
        );

    \I__13853\ : LocalMux
    port map (
            O => \N__61542\,
            I => \N__61530\
        );

    \I__13852\ : CascadeMux
    port map (
            O => \N__61541\,
            I => \N__61527\
        );

    \I__13851\ : Span4Mux_h
    port map (
            O => \N__61538\,
            I => \N__61524\
        );

    \I__13850\ : InMux
    port map (
            O => \N__61535\,
            I => \N__61521\
        );

    \I__13849\ : Span4Mux_v
    port map (
            O => \N__61530\,
            I => \N__61518\
        );

    \I__13848\ : InMux
    port map (
            O => \N__61527\,
            I => \N__61515\
        );

    \I__13847\ : Span4Mux_v
    port map (
            O => \N__61524\,
            I => \N__61512\
        );

    \I__13846\ : LocalMux
    port map (
            O => \N__61521\,
            I => \c0.data_in_frame_8_0\
        );

    \I__13845\ : Odrv4
    port map (
            O => \N__61518\,
            I => \c0.data_in_frame_8_0\
        );

    \I__13844\ : LocalMux
    port map (
            O => \N__61515\,
            I => \c0.data_in_frame_8_0\
        );

    \I__13843\ : Odrv4
    port map (
            O => \N__61512\,
            I => \c0.data_in_frame_8_0\
        );

    \I__13842\ : CascadeMux
    port map (
            O => \N__61503\,
            I => \N__61500\
        );

    \I__13841\ : InMux
    port map (
            O => \N__61500\,
            I => \N__61497\
        );

    \I__13840\ : LocalMux
    port map (
            O => \N__61497\,
            I => \N__61494\
        );

    \I__13839\ : Span4Mux_v
    port map (
            O => \N__61494\,
            I => \N__61491\
        );

    \I__13838\ : Odrv4
    port map (
            O => \N__61491\,
            I => \c0.n104\
        );

    \I__13837\ : InMux
    port map (
            O => \N__61488\,
            I => \N__61482\
        );

    \I__13836\ : InMux
    port map (
            O => \N__61487\,
            I => \N__61482\
        );

    \I__13835\ : LocalMux
    port map (
            O => \N__61482\,
            I => \c0.n7_adj_4253\
        );

    \I__13834\ : CascadeMux
    port map (
            O => \N__61479\,
            I => \N__61476\
        );

    \I__13833\ : InMux
    port map (
            O => \N__61476\,
            I => \N__61470\
        );

    \I__13832\ : InMux
    port map (
            O => \N__61475\,
            I => \N__61470\
        );

    \I__13831\ : LocalMux
    port map (
            O => \N__61470\,
            I => \c0.n5_adj_4252\
        );

    \I__13830\ : InMux
    port map (
            O => \N__61467\,
            I => \N__61463\
        );

    \I__13829\ : InMux
    port map (
            O => \N__61466\,
            I => \N__61460\
        );

    \I__13828\ : LocalMux
    port map (
            O => \N__61463\,
            I => \N__61457\
        );

    \I__13827\ : LocalMux
    port map (
            O => \N__61460\,
            I => \N__61454\
        );

    \I__13826\ : Span4Mux_h
    port map (
            O => \N__61457\,
            I => \N__61451\
        );

    \I__13825\ : Span4Mux_v
    port map (
            O => \N__61454\,
            I => \N__61448\
        );

    \I__13824\ : Span4Mux_h
    port map (
            O => \N__61451\,
            I => \N__61443\
        );

    \I__13823\ : Span4Mux_h
    port map (
            O => \N__61448\,
            I => \N__61443\
        );

    \I__13822\ : Odrv4
    port map (
            O => \N__61443\,
            I => \c0.n5_adj_4443\
        );

    \I__13821\ : CascadeMux
    port map (
            O => \N__61440\,
            I => \c0.n13734_cascade_\
        );

    \I__13820\ : InMux
    port map (
            O => \N__61437\,
            I => \N__61434\
        );

    \I__13819\ : LocalMux
    port map (
            O => \N__61434\,
            I => \N__61430\
        );

    \I__13818\ : InMux
    port map (
            O => \N__61433\,
            I => \N__61426\
        );

    \I__13817\ : Span4Mux_v
    port map (
            O => \N__61430\,
            I => \N__61421\
        );

    \I__13816\ : InMux
    port map (
            O => \N__61429\,
            I => \N__61418\
        );

    \I__13815\ : LocalMux
    port map (
            O => \N__61426\,
            I => \N__61415\
        );

    \I__13814\ : InMux
    port map (
            O => \N__61425\,
            I => \N__61412\
        );

    \I__13813\ : InMux
    port map (
            O => \N__61424\,
            I => \N__61409\
        );

    \I__13812\ : Sp12to4
    port map (
            O => \N__61421\,
            I => \N__61404\
        );

    \I__13811\ : LocalMux
    port map (
            O => \N__61418\,
            I => \N__61404\
        );

    \I__13810\ : Span4Mux_v
    port map (
            O => \N__61415\,
            I => \N__61399\
        );

    \I__13809\ : LocalMux
    port map (
            O => \N__61412\,
            I => \N__61399\
        );

    \I__13808\ : LocalMux
    port map (
            O => \N__61409\,
            I => \c0.n17734\
        );

    \I__13807\ : Odrv12
    port map (
            O => \N__61404\,
            I => \c0.n17734\
        );

    \I__13806\ : Odrv4
    port map (
            O => \N__61399\,
            I => \c0.n17734\
        );

    \I__13805\ : InMux
    port map (
            O => \N__61392\,
            I => \N__61388\
        );

    \I__13804\ : InMux
    port map (
            O => \N__61391\,
            I => \N__61385\
        );

    \I__13803\ : LocalMux
    port map (
            O => \N__61388\,
            I => \N__61381\
        );

    \I__13802\ : LocalMux
    port map (
            O => \N__61385\,
            I => \N__61377\
        );

    \I__13801\ : InMux
    port map (
            O => \N__61384\,
            I => \N__61374\
        );

    \I__13800\ : Span4Mux_v
    port map (
            O => \N__61381\,
            I => \N__61371\
        );

    \I__13799\ : InMux
    port map (
            O => \N__61380\,
            I => \N__61368\
        );

    \I__13798\ : Span4Mux_v
    port map (
            O => \N__61377\,
            I => \N__61363\
        );

    \I__13797\ : LocalMux
    port map (
            O => \N__61374\,
            I => \N__61363\
        );

    \I__13796\ : Sp12to4
    port map (
            O => \N__61371\,
            I => \N__61360\
        );

    \I__13795\ : LocalMux
    port map (
            O => \N__61368\,
            I => \N__61357\
        );

    \I__13794\ : Sp12to4
    port map (
            O => \N__61363\,
            I => \N__61352\
        );

    \I__13793\ : Span12Mux_h
    port map (
            O => \N__61360\,
            I => \N__61352\
        );

    \I__13792\ : Odrv4
    port map (
            O => \N__61357\,
            I => \c0.n12973\
        );

    \I__13791\ : Odrv12
    port map (
            O => \N__61352\,
            I => \c0.n12973\
        );

    \I__13790\ : CascadeMux
    port map (
            O => \N__61347\,
            I => \c0.n30_adj_4705_cascade_\
        );

    \I__13789\ : CascadeMux
    port map (
            O => \N__61344\,
            I => \c0.n23523_cascade_\
        );

    \I__13788\ : InMux
    port map (
            O => \N__61341\,
            I => \N__61338\
        );

    \I__13787\ : LocalMux
    port map (
            O => \N__61338\,
            I => \c0.n30\
        );

    \I__13786\ : InMux
    port map (
            O => \N__61335\,
            I => \N__61330\
        );

    \I__13785\ : InMux
    port map (
            O => \N__61334\,
            I => \N__61327\
        );

    \I__13784\ : InMux
    port map (
            O => \N__61333\,
            I => \N__61324\
        );

    \I__13783\ : LocalMux
    port map (
            O => \N__61330\,
            I => \N__61321\
        );

    \I__13782\ : LocalMux
    port map (
            O => \N__61327\,
            I => \N__61316\
        );

    \I__13781\ : LocalMux
    port map (
            O => \N__61324\,
            I => \N__61316\
        );

    \I__13780\ : Span12Mux_h
    port map (
            O => \N__61321\,
            I => \N__61313\
        );

    \I__13779\ : Span12Mux_h
    port map (
            O => \N__61316\,
            I => \N__61310\
        );

    \I__13778\ : Odrv12
    port map (
            O => \N__61313\,
            I => \c0.n13075\
        );

    \I__13777\ : Odrv12
    port map (
            O => \N__61310\,
            I => \c0.n13075\
        );

    \I__13776\ : CascadeMux
    port map (
            O => \N__61305\,
            I => \c0.n7_adj_4634_cascade_\
        );

    \I__13775\ : InMux
    port map (
            O => \N__61302\,
            I => \N__61299\
        );

    \I__13774\ : LocalMux
    port map (
            O => \N__61299\,
            I => \N__61295\
        );

    \I__13773\ : CascadeMux
    port map (
            O => \N__61298\,
            I => \N__61289\
        );

    \I__13772\ : Span4Mux_h
    port map (
            O => \N__61295\,
            I => \N__61285\
        );

    \I__13771\ : InMux
    port map (
            O => \N__61294\,
            I => \N__61282\
        );

    \I__13770\ : InMux
    port map (
            O => \N__61293\,
            I => \N__61277\
        );

    \I__13769\ : InMux
    port map (
            O => \N__61292\,
            I => \N__61277\
        );

    \I__13768\ : InMux
    port map (
            O => \N__61289\,
            I => \N__61272\
        );

    \I__13767\ : InMux
    port map (
            O => \N__61288\,
            I => \N__61272\
        );

    \I__13766\ : Odrv4
    port map (
            O => \N__61285\,
            I => \c0.n22230\
        );

    \I__13765\ : LocalMux
    port map (
            O => \N__61282\,
            I => \c0.n22230\
        );

    \I__13764\ : LocalMux
    port map (
            O => \N__61277\,
            I => \c0.n22230\
        );

    \I__13763\ : LocalMux
    port map (
            O => \N__61272\,
            I => \c0.n22230\
        );

    \I__13762\ : InMux
    port map (
            O => \N__61263\,
            I => \N__61259\
        );

    \I__13761\ : InMux
    port map (
            O => \N__61262\,
            I => \N__61256\
        );

    \I__13760\ : LocalMux
    port map (
            O => \N__61259\,
            I => \N__61252\
        );

    \I__13759\ : LocalMux
    port map (
            O => \N__61256\,
            I => \N__61249\
        );

    \I__13758\ : InMux
    port map (
            O => \N__61255\,
            I => \N__61246\
        );

    \I__13757\ : Span4Mux_v
    port map (
            O => \N__61252\,
            I => \N__61242\
        );

    \I__13756\ : Span4Mux_v
    port map (
            O => \N__61249\,
            I => \N__61239\
        );

    \I__13755\ : LocalMux
    port map (
            O => \N__61246\,
            I => \N__61236\
        );

    \I__13754\ : InMux
    port map (
            O => \N__61245\,
            I => \N__61232\
        );

    \I__13753\ : Span4Mux_v
    port map (
            O => \N__61242\,
            I => \N__61227\
        );

    \I__13752\ : Span4Mux_v
    port map (
            O => \N__61239\,
            I => \N__61227\
        );

    \I__13751\ : Span4Mux_h
    port map (
            O => \N__61236\,
            I => \N__61224\
        );

    \I__13750\ : InMux
    port map (
            O => \N__61235\,
            I => \N__61221\
        );

    \I__13749\ : LocalMux
    port map (
            O => \N__61232\,
            I => \c0.data_in_frame_9_4\
        );

    \I__13748\ : Odrv4
    port map (
            O => \N__61227\,
            I => \c0.data_in_frame_9_4\
        );

    \I__13747\ : Odrv4
    port map (
            O => \N__61224\,
            I => \c0.data_in_frame_9_4\
        );

    \I__13746\ : LocalMux
    port map (
            O => \N__61221\,
            I => \c0.data_in_frame_9_4\
        );

    \I__13745\ : CascadeMux
    port map (
            O => \N__61212\,
            I => \N__61209\
        );

    \I__13744\ : InMux
    port map (
            O => \N__61209\,
            I => \N__61206\
        );

    \I__13743\ : LocalMux
    port map (
            O => \N__61206\,
            I => \N__61203\
        );

    \I__13742\ : Span4Mux_h
    port map (
            O => \N__61203\,
            I => \N__61200\
        );

    \I__13741\ : Span4Mux_v
    port map (
            O => \N__61200\,
            I => \N__61197\
        );

    \I__13740\ : Odrv4
    port map (
            O => \N__61197\,
            I => \c0.n150\
        );

    \I__13739\ : InMux
    port map (
            O => \N__61194\,
            I => \N__61191\
        );

    \I__13738\ : LocalMux
    port map (
            O => \N__61191\,
            I => \N__61188\
        );

    \I__13737\ : Span4Mux_v
    port map (
            O => \N__61188\,
            I => \N__61185\
        );

    \I__13736\ : Span4Mux_h
    port map (
            O => \N__61185\,
            I => \N__61182\
        );

    \I__13735\ : Span4Mux_h
    port map (
            O => \N__61182\,
            I => \N__61179\
        );

    \I__13734\ : Odrv4
    port map (
            O => \N__61179\,
            I => \c0.n13651\
        );

    \I__13733\ : CascadeMux
    port map (
            O => \N__61176\,
            I => \N__61172\
        );

    \I__13732\ : InMux
    port map (
            O => \N__61175\,
            I => \N__61169\
        );

    \I__13731\ : InMux
    port map (
            O => \N__61172\,
            I => \N__61166\
        );

    \I__13730\ : LocalMux
    port map (
            O => \N__61169\,
            I => \N__61163\
        );

    \I__13729\ : LocalMux
    port map (
            O => \N__61166\,
            I => \N__61160\
        );

    \I__13728\ : Span4Mux_v
    port map (
            O => \N__61163\,
            I => \N__61157\
        );

    \I__13727\ : Odrv4
    port map (
            O => \N__61160\,
            I => \c0.n18_adj_4228\
        );

    \I__13726\ : Odrv4
    port map (
            O => \N__61157\,
            I => \c0.n18_adj_4228\
        );

    \I__13725\ : CascadeMux
    port map (
            O => \N__61152\,
            I => \c0.n27_cascade_\
        );

    \I__13724\ : InMux
    port map (
            O => \N__61149\,
            I => \N__61146\
        );

    \I__13723\ : LocalMux
    port map (
            O => \N__61146\,
            I => \N__61143\
        );

    \I__13722\ : Span4Mux_h
    port map (
            O => \N__61143\,
            I => \N__61139\
        );

    \I__13721\ : InMux
    port map (
            O => \N__61142\,
            I => \N__61136\
        );

    \I__13720\ : Span4Mux_h
    port map (
            O => \N__61139\,
            I => \N__61133\
        );

    \I__13719\ : LocalMux
    port map (
            O => \N__61136\,
            I => \c0.n19\
        );

    \I__13718\ : Odrv4
    port map (
            O => \N__61133\,
            I => \c0.n19\
        );

    \I__13717\ : CascadeMux
    port map (
            O => \N__61128\,
            I => \c0.n23528_cascade_\
        );

    \I__13716\ : CascadeMux
    port map (
            O => \N__61125\,
            I => \c0.n34_adj_4278_cascade_\
        );

    \I__13715\ : InMux
    port map (
            O => \N__61122\,
            I => \N__61119\
        );

    \I__13714\ : LocalMux
    port map (
            O => \N__61119\,
            I => \N__61116\
        );

    \I__13713\ : Odrv4
    port map (
            O => \N__61116\,
            I => \c0.n36\
        );

    \I__13712\ : InMux
    port map (
            O => \N__61113\,
            I => \N__61104\
        );

    \I__13711\ : InMux
    port map (
            O => \N__61112\,
            I => \N__61104\
        );

    \I__13710\ : InMux
    port map (
            O => \N__61111\,
            I => \N__61104\
        );

    \I__13709\ : LocalMux
    port map (
            O => \N__61104\,
            I => \c0.n48_adj_4227\
        );

    \I__13708\ : InMux
    port map (
            O => \N__61101\,
            I => \N__61098\
        );

    \I__13707\ : LocalMux
    port map (
            O => \N__61098\,
            I => \N__61095\
        );

    \I__13706\ : Span4Mux_v
    port map (
            O => \N__61095\,
            I => \N__61091\
        );

    \I__13705\ : InMux
    port map (
            O => \N__61094\,
            I => \N__61088\
        );

    \I__13704\ : Odrv4
    port map (
            O => \N__61091\,
            I => \c0.n18_adj_4314\
        );

    \I__13703\ : LocalMux
    port map (
            O => \N__61088\,
            I => \c0.n18_adj_4314\
        );

    \I__13702\ : CascadeMux
    port map (
            O => \N__61083\,
            I => \N__61080\
        );

    \I__13701\ : InMux
    port map (
            O => \N__61080\,
            I => \N__61077\
        );

    \I__13700\ : LocalMux
    port map (
            O => \N__61077\,
            I => \N__61074\
        );

    \I__13699\ : Span4Mux_h
    port map (
            O => \N__61074\,
            I => \N__61071\
        );

    \I__13698\ : Odrv4
    port map (
            O => \N__61071\,
            I => \c0.n24_adj_4724\
        );

    \I__13697\ : InMux
    port map (
            O => \N__61068\,
            I => \N__61065\
        );

    \I__13696\ : LocalMux
    port map (
            O => \N__61065\,
            I => \N__61061\
        );

    \I__13695\ : CascadeMux
    port map (
            O => \N__61064\,
            I => \N__61058\
        );

    \I__13694\ : Span4Mux_v
    port map (
            O => \N__61061\,
            I => \N__61054\
        );

    \I__13693\ : InMux
    port map (
            O => \N__61058\,
            I => \N__61051\
        );

    \I__13692\ : InMux
    port map (
            O => \N__61057\,
            I => \N__61048\
        );

    \I__13691\ : Span4Mux_v
    port map (
            O => \N__61054\,
            I => \N__61045\
        );

    \I__13690\ : LocalMux
    port map (
            O => \N__61051\,
            I => \N__61040\
        );

    \I__13689\ : LocalMux
    port map (
            O => \N__61048\,
            I => \N__61037\
        );

    \I__13688\ : Span4Mux_v
    port map (
            O => \N__61045\,
            I => \N__61032\
        );

    \I__13687\ : InMux
    port map (
            O => \N__61044\,
            I => \N__61025\
        );

    \I__13686\ : InMux
    port map (
            O => \N__61043\,
            I => \N__61025\
        );

    \I__13685\ : Span4Mux_v
    port map (
            O => \N__61040\,
            I => \N__61020\
        );

    \I__13684\ : Span4Mux_v
    port map (
            O => \N__61037\,
            I => \N__61020\
        );

    \I__13683\ : InMux
    port map (
            O => \N__61036\,
            I => \N__61017\
        );

    \I__13682\ : InMux
    port map (
            O => \N__61035\,
            I => \N__61014\
        );

    \I__13681\ : Span4Mux_h
    port map (
            O => \N__61032\,
            I => \N__61011\
        );

    \I__13680\ : InMux
    port map (
            O => \N__61031\,
            I => \N__61008\
        );

    \I__13679\ : InMux
    port map (
            O => \N__61030\,
            I => \N__61005\
        );

    \I__13678\ : LocalMux
    port map (
            O => \N__61025\,
            I => \N__60998\
        );

    \I__13677\ : Sp12to4
    port map (
            O => \N__61020\,
            I => \N__60998\
        );

    \I__13676\ : LocalMux
    port map (
            O => \N__61017\,
            I => \N__60998\
        );

    \I__13675\ : LocalMux
    port map (
            O => \N__61014\,
            I => data_in_frame_1_0
        );

    \I__13674\ : Odrv4
    port map (
            O => \N__61011\,
            I => data_in_frame_1_0
        );

    \I__13673\ : LocalMux
    port map (
            O => \N__61008\,
            I => data_in_frame_1_0
        );

    \I__13672\ : LocalMux
    port map (
            O => \N__61005\,
            I => data_in_frame_1_0
        );

    \I__13671\ : Odrv12
    port map (
            O => \N__60998\,
            I => data_in_frame_1_0
        );

    \I__13670\ : InMux
    port map (
            O => \N__60987\,
            I => \N__60984\
        );

    \I__13669\ : LocalMux
    port map (
            O => \N__60984\,
            I => \c0.n5_adj_4711\
        );

    \I__13668\ : InMux
    port map (
            O => \N__60981\,
            I => \N__60978\
        );

    \I__13667\ : LocalMux
    port map (
            O => \N__60978\,
            I => \N__60975\
        );

    \I__13666\ : Span4Mux_v
    port map (
            O => \N__60975\,
            I => \N__60972\
        );

    \I__13665\ : Odrv4
    port map (
            O => \N__60972\,
            I => \c0.n16_adj_4716\
        );

    \I__13664\ : CascadeMux
    port map (
            O => \N__60969\,
            I => \c0.n28_adj_4718_cascade_\
        );

    \I__13663\ : InMux
    port map (
            O => \N__60966\,
            I => \N__60963\
        );

    \I__13662\ : LocalMux
    port map (
            O => \N__60963\,
            I => \N__60960\
        );

    \I__13661\ : Odrv4
    port map (
            O => \N__60960\,
            I => \c0.n24_adj_4717\
        );

    \I__13660\ : InMux
    port map (
            O => \N__60957\,
            I => \N__60954\
        );

    \I__13659\ : LocalMux
    port map (
            O => \N__60954\,
            I => \N__60949\
        );

    \I__13658\ : CascadeMux
    port map (
            O => \N__60953\,
            I => \N__60946\
        );

    \I__13657\ : CascadeMux
    port map (
            O => \N__60952\,
            I => \N__60943\
        );

    \I__13656\ : Span4Mux_h
    port map (
            O => \N__60949\,
            I => \N__60939\
        );

    \I__13655\ : InMux
    port map (
            O => \N__60946\,
            I => \N__60934\
        );

    \I__13654\ : InMux
    port map (
            O => \N__60943\,
            I => \N__60934\
        );

    \I__13653\ : InMux
    port map (
            O => \N__60942\,
            I => \N__60931\
        );

    \I__13652\ : Odrv4
    port map (
            O => \N__60939\,
            I => \c0.n23_adj_4599\
        );

    \I__13651\ : LocalMux
    port map (
            O => \N__60934\,
            I => \c0.n23_adj_4599\
        );

    \I__13650\ : LocalMux
    port map (
            O => \N__60931\,
            I => \c0.n23_adj_4599\
        );

    \I__13649\ : InMux
    port map (
            O => \N__60924\,
            I => \N__60921\
        );

    \I__13648\ : LocalMux
    port map (
            O => \N__60921\,
            I => \N__60918\
        );

    \I__13647\ : Odrv4
    port map (
            O => \N__60918\,
            I => \c0.n4_adj_4446\
        );

    \I__13646\ : CascadeMux
    port map (
            O => \N__60915\,
            I => \c0.n4_adj_4446_cascade_\
        );

    \I__13645\ : InMux
    port map (
            O => \N__60912\,
            I => \N__60909\
        );

    \I__13644\ : LocalMux
    port map (
            O => \N__60909\,
            I => \c0.n26_adj_4714\
        );

    \I__13643\ : InMux
    port map (
            O => \N__60906\,
            I => \N__60900\
        );

    \I__13642\ : InMux
    port map (
            O => \N__60905\,
            I => \N__60900\
        );

    \I__13641\ : LocalMux
    port map (
            O => \N__60900\,
            I => \N__60896\
        );

    \I__13640\ : CascadeMux
    port map (
            O => \N__60899\,
            I => \N__60892\
        );

    \I__13639\ : Span4Mux_v
    port map (
            O => \N__60896\,
            I => \N__60888\
        );

    \I__13638\ : CascadeMux
    port map (
            O => \N__60895\,
            I => \N__60885\
        );

    \I__13637\ : InMux
    port map (
            O => \N__60892\,
            I => \N__60877\
        );

    \I__13636\ : InMux
    port map (
            O => \N__60891\,
            I => \N__60877\
        );

    \I__13635\ : Span4Mux_h
    port map (
            O => \N__60888\,
            I => \N__60874\
        );

    \I__13634\ : InMux
    port map (
            O => \N__60885\,
            I => \N__60867\
        );

    \I__13633\ : InMux
    port map (
            O => \N__60884\,
            I => \N__60867\
        );

    \I__13632\ : InMux
    port map (
            O => \N__60883\,
            I => \N__60867\
        );

    \I__13631\ : InMux
    port map (
            O => \N__60882\,
            I => \N__60864\
        );

    \I__13630\ : LocalMux
    port map (
            O => \N__60877\,
            I => \c0.data_in_frame_4_0\
        );

    \I__13629\ : Odrv4
    port map (
            O => \N__60874\,
            I => \c0.data_in_frame_4_0\
        );

    \I__13628\ : LocalMux
    port map (
            O => \N__60867\,
            I => \c0.data_in_frame_4_0\
        );

    \I__13627\ : LocalMux
    port map (
            O => \N__60864\,
            I => \c0.data_in_frame_4_0\
        );

    \I__13626\ : InMux
    port map (
            O => \N__60855\,
            I => \N__60851\
        );

    \I__13625\ : InMux
    port map (
            O => \N__60854\,
            I => \N__60847\
        );

    \I__13624\ : LocalMux
    port map (
            O => \N__60851\,
            I => \N__60844\
        );

    \I__13623\ : InMux
    port map (
            O => \N__60850\,
            I => \N__60841\
        );

    \I__13622\ : LocalMux
    port map (
            O => \N__60847\,
            I => \N__60836\
        );

    \I__13621\ : Span4Mux_v
    port map (
            O => \N__60844\,
            I => \N__60836\
        );

    \I__13620\ : LocalMux
    port map (
            O => \N__60841\,
            I => \N__60829\
        );

    \I__13619\ : Span4Mux_h
    port map (
            O => \N__60836\,
            I => \N__60829\
        );

    \I__13618\ : InMux
    port map (
            O => \N__60835\,
            I => \N__60824\
        );

    \I__13617\ : InMux
    port map (
            O => \N__60834\,
            I => \N__60824\
        );

    \I__13616\ : Odrv4
    port map (
            O => \N__60829\,
            I => \c0.data_in_frame_3_6\
        );

    \I__13615\ : LocalMux
    port map (
            O => \N__60824\,
            I => \c0.data_in_frame_3_6\
        );

    \I__13614\ : InMux
    port map (
            O => \N__60819\,
            I => \N__60814\
        );

    \I__13613\ : InMux
    port map (
            O => \N__60818\,
            I => \N__60809\
        );

    \I__13612\ : InMux
    port map (
            O => \N__60817\,
            I => \N__60809\
        );

    \I__13611\ : LocalMux
    port map (
            O => \N__60814\,
            I => \N__60806\
        );

    \I__13610\ : LocalMux
    port map (
            O => \N__60809\,
            I => \N__60803\
        );

    \I__13609\ : Odrv4
    port map (
            O => \N__60806\,
            I => \c0.n23597\
        );

    \I__13608\ : Odrv4
    port map (
            O => \N__60803\,
            I => \c0.n23597\
        );

    \I__13607\ : CascadeMux
    port map (
            O => \N__60798\,
            I => \N__60793\
        );

    \I__13606\ : CascadeMux
    port map (
            O => \N__60797\,
            I => \N__60789\
        );

    \I__13605\ : CascadeMux
    port map (
            O => \N__60796\,
            I => \N__60786\
        );

    \I__13604\ : InMux
    port map (
            O => \N__60793\,
            I => \N__60783\
        );

    \I__13603\ : InMux
    port map (
            O => \N__60792\,
            I => \N__60780\
        );

    \I__13602\ : InMux
    port map (
            O => \N__60789\,
            I => \N__60775\
        );

    \I__13601\ : InMux
    port map (
            O => \N__60786\,
            I => \N__60775\
        );

    \I__13600\ : LocalMux
    port map (
            O => \N__60783\,
            I => \N__60770\
        );

    \I__13599\ : LocalMux
    port map (
            O => \N__60780\,
            I => \N__60765\
        );

    \I__13598\ : LocalMux
    port map (
            O => \N__60775\,
            I => \N__60765\
        );

    \I__13597\ : InMux
    port map (
            O => \N__60774\,
            I => \N__60760\
        );

    \I__13596\ : InMux
    port map (
            O => \N__60773\,
            I => \N__60760\
        );

    \I__13595\ : Odrv12
    port map (
            O => \N__60770\,
            I => \c0.data_in_frame_2_0\
        );

    \I__13594\ : Odrv4
    port map (
            O => \N__60765\,
            I => \c0.data_in_frame_2_0\
        );

    \I__13593\ : LocalMux
    port map (
            O => \N__60760\,
            I => \c0.data_in_frame_2_0\
        );

    \I__13592\ : CascadeMux
    port map (
            O => \N__60753\,
            I => \c0.n37_cascade_\
        );

    \I__13591\ : CascadeMux
    port map (
            O => \N__60750\,
            I => \c0.n22647_cascade_\
        );

    \I__13590\ : CascadeMux
    port map (
            O => \N__60747\,
            I => \N__60743\
        );

    \I__13589\ : CascadeMux
    port map (
            O => \N__60746\,
            I => \N__60738\
        );

    \I__13588\ : InMux
    port map (
            O => \N__60743\,
            I => \N__60734\
        );

    \I__13587\ : InMux
    port map (
            O => \N__60742\,
            I => \N__60731\
        );

    \I__13586\ : InMux
    port map (
            O => \N__60741\,
            I => \N__60728\
        );

    \I__13585\ : InMux
    port map (
            O => \N__60738\,
            I => \N__60723\
        );

    \I__13584\ : InMux
    port map (
            O => \N__60737\,
            I => \N__60723\
        );

    \I__13583\ : LocalMux
    port map (
            O => \N__60734\,
            I => \c0.data_in_frame_2_6\
        );

    \I__13582\ : LocalMux
    port map (
            O => \N__60731\,
            I => \c0.data_in_frame_2_6\
        );

    \I__13581\ : LocalMux
    port map (
            O => \N__60728\,
            I => \c0.data_in_frame_2_6\
        );

    \I__13580\ : LocalMux
    port map (
            O => \N__60723\,
            I => \c0.data_in_frame_2_6\
        );

    \I__13579\ : InMux
    port map (
            O => \N__60714\,
            I => \N__60711\
        );

    \I__13578\ : LocalMux
    port map (
            O => \N__60711\,
            I => \N__60708\
        );

    \I__13577\ : Span4Mux_h
    port map (
            O => \N__60708\,
            I => \N__60705\
        );

    \I__13576\ : Span4Mux_h
    port map (
            O => \N__60705\,
            I => \N__60702\
        );

    \I__13575\ : Odrv4
    port map (
            O => \N__60702\,
            I => \c0.n24747\
        );

    \I__13574\ : InMux
    port map (
            O => \N__60699\,
            I => \N__60696\
        );

    \I__13573\ : LocalMux
    port map (
            O => \N__60696\,
            I => \c0.n10_adj_4722\
        );

    \I__13572\ : CascadeMux
    port map (
            O => \N__60693\,
            I => \c0.n14_adj_4616_cascade_\
        );

    \I__13571\ : InMux
    port map (
            O => \N__60690\,
            I => \N__60687\
        );

    \I__13570\ : LocalMux
    port map (
            O => \N__60687\,
            I => \N__60683\
        );

    \I__13569\ : InMux
    port map (
            O => \N__60686\,
            I => \N__60680\
        );

    \I__13568\ : Span4Mux_v
    port map (
            O => \N__60683\,
            I => \N__60677\
        );

    \I__13567\ : LocalMux
    port map (
            O => \N__60680\,
            I => \N__60674\
        );

    \I__13566\ : Span4Mux_h
    port map (
            O => \N__60677\,
            I => \N__60671\
        );

    \I__13565\ : Odrv4
    port map (
            O => \N__60674\,
            I => \c0.n23666\
        );

    \I__13564\ : Odrv4
    port map (
            O => \N__60671\,
            I => \c0.n23666\
        );

    \I__13563\ : CascadeMux
    port map (
            O => \N__60666\,
            I => \N__60663\
        );

    \I__13562\ : InMux
    port map (
            O => \N__60663\,
            I => \N__60660\
        );

    \I__13561\ : LocalMux
    port map (
            O => \N__60660\,
            I => \N__60657\
        );

    \I__13560\ : Odrv4
    port map (
            O => \N__60657\,
            I => \c0.n37\
        );

    \I__13559\ : InMux
    port map (
            O => \N__60654\,
            I => \N__60651\
        );

    \I__13558\ : LocalMux
    port map (
            O => \N__60651\,
            I => \c0.n55\
        );

    \I__13557\ : CascadeMux
    port map (
            O => \N__60648\,
            I => \N__60645\
        );

    \I__13556\ : InMux
    port map (
            O => \N__60645\,
            I => \N__60641\
        );

    \I__13555\ : InMux
    port map (
            O => \N__60644\,
            I => \N__60638\
        );

    \I__13554\ : LocalMux
    port map (
            O => \N__60641\,
            I => \N__60628\
        );

    \I__13553\ : LocalMux
    port map (
            O => \N__60638\,
            I => \N__60625\
        );

    \I__13552\ : InMux
    port map (
            O => \N__60637\,
            I => \N__60620\
        );

    \I__13551\ : InMux
    port map (
            O => \N__60636\,
            I => \N__60620\
        );

    \I__13550\ : InMux
    port map (
            O => \N__60635\,
            I => \N__60617\
        );

    \I__13549\ : InMux
    port map (
            O => \N__60634\,
            I => \N__60610\
        );

    \I__13548\ : InMux
    port map (
            O => \N__60633\,
            I => \N__60610\
        );

    \I__13547\ : InMux
    port map (
            O => \N__60632\,
            I => \N__60610\
        );

    \I__13546\ : InMux
    port map (
            O => \N__60631\,
            I => \N__60607\
        );

    \I__13545\ : Odrv4
    port map (
            O => \N__60628\,
            I => \c0.data_in_frame_0_6\
        );

    \I__13544\ : Odrv4
    port map (
            O => \N__60625\,
            I => \c0.data_in_frame_0_6\
        );

    \I__13543\ : LocalMux
    port map (
            O => \N__60620\,
            I => \c0.data_in_frame_0_6\
        );

    \I__13542\ : LocalMux
    port map (
            O => \N__60617\,
            I => \c0.data_in_frame_0_6\
        );

    \I__13541\ : LocalMux
    port map (
            O => \N__60610\,
            I => \c0.data_in_frame_0_6\
        );

    \I__13540\ : LocalMux
    port map (
            O => \N__60607\,
            I => \c0.data_in_frame_0_6\
        );

    \I__13539\ : InMux
    port map (
            O => \N__60594\,
            I => \N__60591\
        );

    \I__13538\ : LocalMux
    port map (
            O => \N__60591\,
            I => \c0.n24016\
        );

    \I__13537\ : InMux
    port map (
            O => \N__60588\,
            I => \N__60585\
        );

    \I__13536\ : LocalMux
    port map (
            O => \N__60585\,
            I => \N__60582\
        );

    \I__13535\ : Span4Mux_h
    port map (
            O => \N__60582\,
            I => \N__60579\
        );

    \I__13534\ : Span4Mux_h
    port map (
            O => \N__60579\,
            I => \N__60576\
        );

    \I__13533\ : Odrv4
    port map (
            O => \N__60576\,
            I => \c0.n24749\
        );

    \I__13532\ : InMux
    port map (
            O => \N__60573\,
            I => \N__60570\
        );

    \I__13531\ : LocalMux
    port map (
            O => \N__60570\,
            I => \N__60567\
        );

    \I__13530\ : Span4Mux_v
    port map (
            O => \N__60567\,
            I => \N__60563\
        );

    \I__13529\ : InMux
    port map (
            O => \N__60566\,
            I => \N__60559\
        );

    \I__13528\ : Span4Mux_h
    port map (
            O => \N__60563\,
            I => \N__60554\
        );

    \I__13527\ : CascadeMux
    port map (
            O => \N__60562\,
            I => \N__60549\
        );

    \I__13526\ : LocalMux
    port map (
            O => \N__60559\,
            I => \N__60542\
        );

    \I__13525\ : InMux
    port map (
            O => \N__60558\,
            I => \N__60537\
        );

    \I__13524\ : InMux
    port map (
            O => \N__60557\,
            I => \N__60537\
        );

    \I__13523\ : Sp12to4
    port map (
            O => \N__60554\,
            I => \N__60530\
        );

    \I__13522\ : InMux
    port map (
            O => \N__60553\,
            I => \N__60527\
        );

    \I__13521\ : InMux
    port map (
            O => \N__60552\,
            I => \N__60524\
        );

    \I__13520\ : InMux
    port map (
            O => \N__60549\,
            I => \N__60521\
        );

    \I__13519\ : InMux
    port map (
            O => \N__60548\,
            I => \N__60518\
        );

    \I__13518\ : InMux
    port map (
            O => \N__60547\,
            I => \N__60515\
        );

    \I__13517\ : CascadeMux
    port map (
            O => \N__60546\,
            I => \N__60512\
        );

    \I__13516\ : CascadeMux
    port map (
            O => \N__60545\,
            I => \N__60508\
        );

    \I__13515\ : Span4Mux_v
    port map (
            O => \N__60542\,
            I => \N__60504\
        );

    \I__13514\ : LocalMux
    port map (
            O => \N__60537\,
            I => \N__60501\
        );

    \I__13513\ : InMux
    port map (
            O => \N__60536\,
            I => \N__60494\
        );

    \I__13512\ : InMux
    port map (
            O => \N__60535\,
            I => \N__60494\
        );

    \I__13511\ : InMux
    port map (
            O => \N__60534\,
            I => \N__60494\
        );

    \I__13510\ : CascadeMux
    port map (
            O => \N__60533\,
            I => \N__60491\
        );

    \I__13509\ : Span12Mux_h
    port map (
            O => \N__60530\,
            I => \N__60481\
        );

    \I__13508\ : LocalMux
    port map (
            O => \N__60527\,
            I => \N__60481\
        );

    \I__13507\ : LocalMux
    port map (
            O => \N__60524\,
            I => \N__60481\
        );

    \I__13506\ : LocalMux
    port map (
            O => \N__60521\,
            I => \N__60481\
        );

    \I__13505\ : LocalMux
    port map (
            O => \N__60518\,
            I => \N__60478\
        );

    \I__13504\ : LocalMux
    port map (
            O => \N__60515\,
            I => \N__60475\
        );

    \I__13503\ : InMux
    port map (
            O => \N__60512\,
            I => \N__60470\
        );

    \I__13502\ : InMux
    port map (
            O => \N__60511\,
            I => \N__60470\
        );

    \I__13501\ : InMux
    port map (
            O => \N__60508\,
            I => \N__60465\
        );

    \I__13500\ : InMux
    port map (
            O => \N__60507\,
            I => \N__60465\
        );

    \I__13499\ : Span4Mux_h
    port map (
            O => \N__60504\,
            I => \N__60458\
        );

    \I__13498\ : Span4Mux_h
    port map (
            O => \N__60501\,
            I => \N__60458\
        );

    \I__13497\ : LocalMux
    port map (
            O => \N__60494\,
            I => \N__60458\
        );

    \I__13496\ : InMux
    port map (
            O => \N__60491\,
            I => \N__60453\
        );

    \I__13495\ : InMux
    port map (
            O => \N__60490\,
            I => \N__60453\
        );

    \I__13494\ : Odrv12
    port map (
            O => \N__60481\,
            I => data_in_frame_1_4
        );

    \I__13493\ : Odrv4
    port map (
            O => \N__60478\,
            I => data_in_frame_1_4
        );

    \I__13492\ : Odrv4
    port map (
            O => \N__60475\,
            I => data_in_frame_1_4
        );

    \I__13491\ : LocalMux
    port map (
            O => \N__60470\,
            I => data_in_frame_1_4
        );

    \I__13490\ : LocalMux
    port map (
            O => \N__60465\,
            I => data_in_frame_1_4
        );

    \I__13489\ : Odrv4
    port map (
            O => \N__60458\,
            I => data_in_frame_1_4
        );

    \I__13488\ : LocalMux
    port map (
            O => \N__60453\,
            I => data_in_frame_1_4
        );

    \I__13487\ : InMux
    port map (
            O => \N__60438\,
            I => \N__60435\
        );

    \I__13486\ : LocalMux
    port map (
            O => \N__60435\,
            I => \N__60432\
        );

    \I__13485\ : Span4Mux_v
    port map (
            O => \N__60432\,
            I => \N__60428\
        );

    \I__13484\ : InMux
    port map (
            O => \N__60431\,
            I => \N__60424\
        );

    \I__13483\ : Span4Mux_h
    port map (
            O => \N__60428\,
            I => \N__60421\
        );

    \I__13482\ : CascadeMux
    port map (
            O => \N__60427\,
            I => \N__60418\
        );

    \I__13481\ : LocalMux
    port map (
            O => \N__60424\,
            I => \N__60410\
        );

    \I__13480\ : Span4Mux_v
    port map (
            O => \N__60421\,
            I => \N__60405\
        );

    \I__13479\ : InMux
    port map (
            O => \N__60418\,
            I => \N__60394\
        );

    \I__13478\ : InMux
    port map (
            O => \N__60417\,
            I => \N__60394\
        );

    \I__13477\ : InMux
    port map (
            O => \N__60416\,
            I => \N__60394\
        );

    \I__13476\ : InMux
    port map (
            O => \N__60415\,
            I => \N__60394\
        );

    \I__13475\ : InMux
    port map (
            O => \N__60414\,
            I => \N__60394\
        );

    \I__13474\ : InMux
    port map (
            O => \N__60413\,
            I => \N__60391\
        );

    \I__13473\ : Span4Mux_h
    port map (
            O => \N__60410\,
            I => \N__60388\
        );

    \I__13472\ : CascadeMux
    port map (
            O => \N__60409\,
            I => \N__60382\
        );

    \I__13471\ : CascadeMux
    port map (
            O => \N__60408\,
            I => \N__60379\
        );

    \I__13470\ : Span4Mux_v
    port map (
            O => \N__60405\,
            I => \N__60372\
        );

    \I__13469\ : LocalMux
    port map (
            O => \N__60394\,
            I => \N__60372\
        );

    \I__13468\ : LocalMux
    port map (
            O => \N__60391\,
            I => \N__60369\
        );

    \I__13467\ : Span4Mux_h
    port map (
            O => \N__60388\,
            I => \N__60366\
        );

    \I__13466\ : InMux
    port map (
            O => \N__60387\,
            I => \N__60363\
        );

    \I__13465\ : InMux
    port map (
            O => \N__60386\,
            I => \N__60360\
        );

    \I__13464\ : InMux
    port map (
            O => \N__60385\,
            I => \N__60357\
        );

    \I__13463\ : InMux
    port map (
            O => \N__60382\,
            I => \N__60354\
        );

    \I__13462\ : InMux
    port map (
            O => \N__60379\,
            I => \N__60347\
        );

    \I__13461\ : InMux
    port map (
            O => \N__60378\,
            I => \N__60347\
        );

    \I__13460\ : InMux
    port map (
            O => \N__60377\,
            I => \N__60347\
        );

    \I__13459\ : Span4Mux_v
    port map (
            O => \N__60372\,
            I => \N__60342\
        );

    \I__13458\ : Span4Mux_v
    port map (
            O => \N__60369\,
            I => \N__60342\
        );

    \I__13457\ : Odrv4
    port map (
            O => \N__60366\,
            I => data_in_frame_1_5
        );

    \I__13456\ : LocalMux
    port map (
            O => \N__60363\,
            I => data_in_frame_1_5
        );

    \I__13455\ : LocalMux
    port map (
            O => \N__60360\,
            I => data_in_frame_1_5
        );

    \I__13454\ : LocalMux
    port map (
            O => \N__60357\,
            I => data_in_frame_1_5
        );

    \I__13453\ : LocalMux
    port map (
            O => \N__60354\,
            I => data_in_frame_1_5
        );

    \I__13452\ : LocalMux
    port map (
            O => \N__60347\,
            I => data_in_frame_1_5
        );

    \I__13451\ : Odrv4
    port map (
            O => \N__60342\,
            I => data_in_frame_1_5
        );

    \I__13450\ : InMux
    port map (
            O => \N__60327\,
            I => \N__60324\
        );

    \I__13449\ : LocalMux
    port map (
            O => \N__60324\,
            I => \N__60321\
        );

    \I__13448\ : Span4Mux_h
    port map (
            O => \N__60321\,
            I => \N__60318\
        );

    \I__13447\ : Span4Mux_h
    port map (
            O => \N__60318\,
            I => \N__60315\
        );

    \I__13446\ : Odrv4
    port map (
            O => \N__60315\,
            I => \c0.n37_adj_4738\
        );

    \I__13445\ : CascadeMux
    port map (
            O => \N__60312\,
            I => \N__60309\
        );

    \I__13444\ : InMux
    port map (
            O => \N__60309\,
            I => \N__60306\
        );

    \I__13443\ : LocalMux
    port map (
            O => \N__60306\,
            I => \N__60298\
        );

    \I__13442\ : InMux
    port map (
            O => \N__60305\,
            I => \N__60292\
        );

    \I__13441\ : InMux
    port map (
            O => \N__60304\,
            I => \N__60289\
        );

    \I__13440\ : InMux
    port map (
            O => \N__60303\,
            I => \N__60284\
        );

    \I__13439\ : InMux
    port map (
            O => \N__60302\,
            I => \N__60284\
        );

    \I__13438\ : InMux
    port map (
            O => \N__60301\,
            I => \N__60280\
        );

    \I__13437\ : Span4Mux_v
    port map (
            O => \N__60298\,
            I => \N__60277\
        );

    \I__13436\ : InMux
    port map (
            O => \N__60297\,
            I => \N__60274\
        );

    \I__13435\ : InMux
    port map (
            O => \N__60296\,
            I => \N__60269\
        );

    \I__13434\ : InMux
    port map (
            O => \N__60295\,
            I => \N__60269\
        );

    \I__13433\ : LocalMux
    port map (
            O => \N__60292\,
            I => \N__60266\
        );

    \I__13432\ : LocalMux
    port map (
            O => \N__60289\,
            I => \N__60261\
        );

    \I__13431\ : LocalMux
    port map (
            O => \N__60284\,
            I => \N__60261\
        );

    \I__13430\ : InMux
    port map (
            O => \N__60283\,
            I => \N__60258\
        );

    \I__13429\ : LocalMux
    port map (
            O => \N__60280\,
            I => \c0.data_in_frame_0_5\
        );

    \I__13428\ : Odrv4
    port map (
            O => \N__60277\,
            I => \c0.data_in_frame_0_5\
        );

    \I__13427\ : LocalMux
    port map (
            O => \N__60274\,
            I => \c0.data_in_frame_0_5\
        );

    \I__13426\ : LocalMux
    port map (
            O => \N__60269\,
            I => \c0.data_in_frame_0_5\
        );

    \I__13425\ : Odrv12
    port map (
            O => \N__60266\,
            I => \c0.data_in_frame_0_5\
        );

    \I__13424\ : Odrv4
    port map (
            O => \N__60261\,
            I => \c0.data_in_frame_0_5\
        );

    \I__13423\ : LocalMux
    port map (
            O => \N__60258\,
            I => \c0.data_in_frame_0_5\
        );

    \I__13422\ : CascadeMux
    port map (
            O => \N__60243\,
            I => \N__60240\
        );

    \I__13421\ : InMux
    port map (
            O => \N__60240\,
            I => \N__60236\
        );

    \I__13420\ : CascadeMux
    port map (
            O => \N__60239\,
            I => \N__60231\
        );

    \I__13419\ : LocalMux
    port map (
            O => \N__60236\,
            I => \N__60224\
        );

    \I__13418\ : InMux
    port map (
            O => \N__60235\,
            I => \N__60219\
        );

    \I__13417\ : InMux
    port map (
            O => \N__60234\,
            I => \N__60219\
        );

    \I__13416\ : InMux
    port map (
            O => \N__60231\,
            I => \N__60212\
        );

    \I__13415\ : InMux
    port map (
            O => \N__60230\,
            I => \N__60212\
        );

    \I__13414\ : InMux
    port map (
            O => \N__60229\,
            I => \N__60212\
        );

    \I__13413\ : CascadeMux
    port map (
            O => \N__60228\,
            I => \N__60209\
        );

    \I__13412\ : CascadeMux
    port map (
            O => \N__60227\,
            I => \N__60205\
        );

    \I__13411\ : Span4Mux_v
    port map (
            O => \N__60224\,
            I => \N__60198\
        );

    \I__13410\ : LocalMux
    port map (
            O => \N__60219\,
            I => \N__60198\
        );

    \I__13409\ : LocalMux
    port map (
            O => \N__60212\,
            I => \N__60195\
        );

    \I__13408\ : InMux
    port map (
            O => \N__60209\,
            I => \N__60188\
        );

    \I__13407\ : InMux
    port map (
            O => \N__60208\,
            I => \N__60188\
        );

    \I__13406\ : InMux
    port map (
            O => \N__60205\,
            I => \N__60188\
        );

    \I__13405\ : InMux
    port map (
            O => \N__60204\,
            I => \N__60183\
        );

    \I__13404\ : InMux
    port map (
            O => \N__60203\,
            I => \N__60180\
        );

    \I__13403\ : Span4Mux_v
    port map (
            O => \N__60198\,
            I => \N__60173\
        );

    \I__13402\ : Span4Mux_h
    port map (
            O => \N__60195\,
            I => \N__60173\
        );

    \I__13401\ : LocalMux
    port map (
            O => \N__60188\,
            I => \N__60173\
        );

    \I__13400\ : InMux
    port map (
            O => \N__60187\,
            I => \N__60168\
        );

    \I__13399\ : InMux
    port map (
            O => \N__60186\,
            I => \N__60168\
        );

    \I__13398\ : LocalMux
    port map (
            O => \N__60183\,
            I => \c0.data_in_frame_0_7\
        );

    \I__13397\ : LocalMux
    port map (
            O => \N__60180\,
            I => \c0.data_in_frame_0_7\
        );

    \I__13396\ : Odrv4
    port map (
            O => \N__60173\,
            I => \c0.data_in_frame_0_7\
        );

    \I__13395\ : LocalMux
    port map (
            O => \N__60168\,
            I => \c0.data_in_frame_0_7\
        );

    \I__13394\ : InMux
    port map (
            O => \N__60159\,
            I => \N__60156\
        );

    \I__13393\ : LocalMux
    port map (
            O => \N__60156\,
            I => \N__60152\
        );

    \I__13392\ : InMux
    port map (
            O => \N__60155\,
            I => \N__60149\
        );

    \I__13391\ : Span4Mux_v
    port map (
            O => \N__60152\,
            I => \N__60143\
        );

    \I__13390\ : LocalMux
    port map (
            O => \N__60149\,
            I => \N__60143\
        );

    \I__13389\ : InMux
    port map (
            O => \N__60148\,
            I => \N__60140\
        );

    \I__13388\ : Odrv4
    port map (
            O => \N__60143\,
            I => \c0.n22316\
        );

    \I__13387\ : LocalMux
    port map (
            O => \N__60140\,
            I => \c0.n22316\
        );

    \I__13386\ : InMux
    port map (
            O => \N__60135\,
            I => \N__60132\
        );

    \I__13385\ : LocalMux
    port map (
            O => \N__60132\,
            I => \N__60128\
        );

    \I__13384\ : InMux
    port map (
            O => \N__60131\,
            I => \N__60125\
        );

    \I__13383\ : Odrv4
    port map (
            O => \N__60128\,
            I => \c0.n23554\
        );

    \I__13382\ : LocalMux
    port map (
            O => \N__60125\,
            I => \c0.n23554\
        );

    \I__13381\ : CascadeMux
    port map (
            O => \N__60120\,
            I => \c0.n34_cascade_\
        );

    \I__13380\ : InMux
    port map (
            O => \N__60117\,
            I => \N__60113\
        );

    \I__13379\ : InMux
    port map (
            O => \N__60116\,
            I => \N__60110\
        );

    \I__13378\ : LocalMux
    port map (
            O => \N__60113\,
            I => \N__60107\
        );

    \I__13377\ : LocalMux
    port map (
            O => \N__60110\,
            I => \N__60102\
        );

    \I__13376\ : Span4Mux_h
    port map (
            O => \N__60107\,
            I => \N__60102\
        );

    \I__13375\ : Odrv4
    port map (
            O => \N__60102\,
            I => \c0.n23655\
        );

    \I__13374\ : InMux
    port map (
            O => \N__60099\,
            I => \N__60096\
        );

    \I__13373\ : LocalMux
    port map (
            O => \N__60096\,
            I => \N__60093\
        );

    \I__13372\ : Span4Mux_h
    port map (
            O => \N__60093\,
            I => \N__60090\
        );

    \I__13371\ : Odrv4
    port map (
            O => \N__60090\,
            I => \c0.n53\
        );

    \I__13370\ : CascadeMux
    port map (
            O => \N__60087\,
            I => \c0.n54_cascade_\
        );

    \I__13369\ : InMux
    port map (
            O => \N__60084\,
            I => \N__60081\
        );

    \I__13368\ : LocalMux
    port map (
            O => \N__60081\,
            I => \N__60077\
        );

    \I__13367\ : InMux
    port map (
            O => \N__60080\,
            I => \N__60074\
        );

    \I__13366\ : Span4Mux_h
    port map (
            O => \N__60077\,
            I => \N__60071\
        );

    \I__13365\ : LocalMux
    port map (
            O => \N__60074\,
            I => \N__60068\
        );

    \I__13364\ : Odrv4
    port map (
            O => \N__60071\,
            I => \c0.n56\
        );

    \I__13363\ : Odrv4
    port map (
            O => \N__60068\,
            I => \c0.n56\
        );

    \I__13362\ : InMux
    port map (
            O => \N__60063\,
            I => \N__60057\
        );

    \I__13361\ : InMux
    port map (
            O => \N__60062\,
            I => \N__60054\
        );

    \I__13360\ : InMux
    port map (
            O => \N__60061\,
            I => \N__60049\
        );

    \I__13359\ : InMux
    port map (
            O => \N__60060\,
            I => \N__60049\
        );

    \I__13358\ : LocalMux
    port map (
            O => \N__60057\,
            I => \N__60045\
        );

    \I__13357\ : LocalMux
    port map (
            O => \N__60054\,
            I => \N__60040\
        );

    \I__13356\ : LocalMux
    port map (
            O => \N__60049\,
            I => \N__60040\
        );

    \I__13355\ : InMux
    port map (
            O => \N__60048\,
            I => \N__60037\
        );

    \I__13354\ : Span4Mux_h
    port map (
            O => \N__60045\,
            I => \N__60030\
        );

    \I__13353\ : Span4Mux_v
    port map (
            O => \N__60040\,
            I => \N__60030\
        );

    \I__13352\ : LocalMux
    port map (
            O => \N__60037\,
            I => \N__60030\
        );

    \I__13351\ : Span4Mux_v
    port map (
            O => \N__60030\,
            I => \N__60026\
        );

    \I__13350\ : InMux
    port map (
            O => \N__60029\,
            I => \N__60023\
        );

    \I__13349\ : Span4Mux_v
    port map (
            O => \N__60026\,
            I => \N__60020\
        );

    \I__13348\ : LocalMux
    port map (
            O => \N__60023\,
            I => \N__60017\
        );

    \I__13347\ : Odrv4
    port map (
            O => \N__60020\,
            I => \c0.n13821\
        );

    \I__13346\ : Odrv4
    port map (
            O => \N__60017\,
            I => \c0.n13821\
        );

    \I__13345\ : InMux
    port map (
            O => \N__60012\,
            I => \N__60009\
        );

    \I__13344\ : LocalMux
    port map (
            O => \N__60009\,
            I => \N__60006\
        );

    \I__13343\ : Odrv4
    port map (
            O => \N__60006\,
            I => \c0.n48\
        );

    \I__13342\ : CascadeMux
    port map (
            O => \N__60003\,
            I => \c0.n24441_cascade_\
        );

    \I__13341\ : InMux
    port map (
            O => \N__60000\,
            I => \N__59997\
        );

    \I__13340\ : LocalMux
    port map (
            O => \N__59997\,
            I => \N__59994\
        );

    \I__13339\ : Span4Mux_h
    port map (
            O => \N__59994\,
            I => \N__59991\
        );

    \I__13338\ : Span4Mux_h
    port map (
            O => \N__59991\,
            I => \N__59988\
        );

    \I__13337\ : Odrv4
    port map (
            O => \N__59988\,
            I => \c0.n30_adj_4545\
        );

    \I__13336\ : InMux
    port map (
            O => \N__59985\,
            I => \N__59982\
        );

    \I__13335\ : LocalMux
    port map (
            O => \N__59982\,
            I => \c0.n72\
        );

    \I__13334\ : InMux
    port map (
            O => \N__59979\,
            I => \N__59976\
        );

    \I__13333\ : LocalMux
    port map (
            O => \N__59976\,
            I => \N__59973\
        );

    \I__13332\ : Span4Mux_v
    port map (
            O => \N__59973\,
            I => \N__59970\
        );

    \I__13331\ : Odrv4
    port map (
            O => \N__59970\,
            I => \c0.n24559\
        );

    \I__13330\ : CascadeMux
    port map (
            O => \N__59967\,
            I => \N__59964\
        );

    \I__13329\ : InMux
    port map (
            O => \N__59964\,
            I => \N__59961\
        );

    \I__13328\ : LocalMux
    port map (
            O => \N__59961\,
            I => \N__59958\
        );

    \I__13327\ : Odrv4
    port map (
            O => \N__59958\,
            I => \c0.n42_adj_4510\
        );

    \I__13326\ : InMux
    port map (
            O => \N__59955\,
            I => \N__59952\
        );

    \I__13325\ : LocalMux
    port map (
            O => \N__59952\,
            I => \c0.n20_adj_4518\
        );

    \I__13324\ : CascadeMux
    port map (
            O => \N__59949\,
            I => \N__59946\
        );

    \I__13323\ : InMux
    port map (
            O => \N__59946\,
            I => \N__59943\
        );

    \I__13322\ : LocalMux
    port map (
            O => \N__59943\,
            I => \N__59940\
        );

    \I__13321\ : Span4Mux_h
    port map (
            O => \N__59940\,
            I => \N__59937\
        );

    \I__13320\ : Odrv4
    port map (
            O => \N__59937\,
            I => \c0.n24751\
        );

    \I__13319\ : CascadeMux
    port map (
            O => \N__59934\,
            I => \c0.n14_adj_4676_cascade_\
        );

    \I__13318\ : InMux
    port map (
            O => \N__59931\,
            I => \N__59928\
        );

    \I__13317\ : LocalMux
    port map (
            O => \N__59928\,
            I => \N__59925\
        );

    \I__13316\ : Span4Mux_h
    port map (
            O => \N__59925\,
            I => \N__59922\
        );

    \I__13315\ : Odrv4
    port map (
            O => \N__59922\,
            I => \c0.data_out_frame_0__7__N_2777\
        );

    \I__13314\ : InMux
    port map (
            O => \N__59919\,
            I => \N__59916\
        );

    \I__13313\ : LocalMux
    port map (
            O => \N__59916\,
            I => \N__59913\
        );

    \I__13312\ : Span4Mux_h
    port map (
            O => \N__59913\,
            I => \N__59909\
        );

    \I__13311\ : InMux
    port map (
            O => \N__59912\,
            I => \N__59906\
        );

    \I__13310\ : Odrv4
    port map (
            O => \N__59909\,
            I => \c0.n10_adj_4513\
        );

    \I__13309\ : LocalMux
    port map (
            O => \N__59906\,
            I => \c0.n10_adj_4513\
        );

    \I__13308\ : InMux
    port map (
            O => \N__59901\,
            I => \N__59898\
        );

    \I__13307\ : LocalMux
    port map (
            O => \N__59898\,
            I => \N__59893\
        );

    \I__13306\ : InMux
    port map (
            O => \N__59897\,
            I => \N__59890\
        );

    \I__13305\ : InMux
    port map (
            O => \N__59896\,
            I => \N__59887\
        );

    \I__13304\ : Odrv4
    port map (
            O => \N__59893\,
            I => \c0.n15_adj_4497\
        );

    \I__13303\ : LocalMux
    port map (
            O => \N__59890\,
            I => \c0.n15_adj_4497\
        );

    \I__13302\ : LocalMux
    port map (
            O => \N__59887\,
            I => \c0.n15_adj_4497\
        );

    \I__13301\ : CascadeMux
    port map (
            O => \N__59880\,
            I => \N__59877\
        );

    \I__13300\ : InMux
    port map (
            O => \N__59877\,
            I => \N__59872\
        );

    \I__13299\ : InMux
    port map (
            O => \N__59876\,
            I => \N__59869\
        );

    \I__13298\ : CascadeMux
    port map (
            O => \N__59875\,
            I => \N__59864\
        );

    \I__13297\ : LocalMux
    port map (
            O => \N__59872\,
            I => \N__59861\
        );

    \I__13296\ : LocalMux
    port map (
            O => \N__59869\,
            I => \N__59858\
        );

    \I__13295\ : InMux
    port map (
            O => \N__59868\,
            I => \N__59853\
        );

    \I__13294\ : InMux
    port map (
            O => \N__59867\,
            I => \N__59853\
        );

    \I__13293\ : InMux
    port map (
            O => \N__59864\,
            I => \N__59850\
        );

    \I__13292\ : Span4Mux_h
    port map (
            O => \N__59861\,
            I => \N__59845\
        );

    \I__13291\ : Span4Mux_h
    port map (
            O => \N__59858\,
            I => \N__59845\
        );

    \I__13290\ : LocalMux
    port map (
            O => \N__59853\,
            I => \c0.data_in_frame_25_4\
        );

    \I__13289\ : LocalMux
    port map (
            O => \N__59850\,
            I => \c0.data_in_frame_25_4\
        );

    \I__13288\ : Odrv4
    port map (
            O => \N__59845\,
            I => \c0.data_in_frame_25_4\
        );

    \I__13287\ : InMux
    port map (
            O => \N__59838\,
            I => \N__59835\
        );

    \I__13286\ : LocalMux
    port map (
            O => \N__59835\,
            I => \N__59832\
        );

    \I__13285\ : Span4Mux_v
    port map (
            O => \N__59832\,
            I => \N__59829\
        );

    \I__13284\ : Odrv4
    port map (
            O => \N__59829\,
            I => \c0.n23_adj_4551\
        );

    \I__13283\ : InMux
    port map (
            O => \N__59826\,
            I => \N__59823\
        );

    \I__13282\ : LocalMux
    port map (
            O => \N__59823\,
            I => \c0.n26_adj_4548\
        );

    \I__13281\ : CascadeMux
    port map (
            O => \N__59820\,
            I => \c0.n24_adj_4550_cascade_\
        );

    \I__13280\ : CascadeMux
    port map (
            O => \N__59817\,
            I => \c0.n21010_cascade_\
        );

    \I__13279\ : InMux
    port map (
            O => \N__59814\,
            I => \N__59811\
        );

    \I__13278\ : LocalMux
    port map (
            O => \N__59811\,
            I => \c0.n53_adj_4538\
        );

    \I__13277\ : InMux
    port map (
            O => \N__59808\,
            I => \N__59805\
        );

    \I__13276\ : LocalMux
    port map (
            O => \N__59805\,
            I => \c0.n61_adj_4543\
        );

    \I__13275\ : InMux
    port map (
            O => \N__59802\,
            I => \N__59799\
        );

    \I__13274\ : LocalMux
    port map (
            O => \N__59799\,
            I => \c0.n42_adj_4540\
        );

    \I__13273\ : CascadeMux
    port map (
            O => \N__59796\,
            I => \N__59793\
        );

    \I__13272\ : InMux
    port map (
            O => \N__59793\,
            I => \N__59790\
        );

    \I__13271\ : LocalMux
    port map (
            O => \N__59790\,
            I => \c0.n62_adj_4541\
        );

    \I__13270\ : CascadeMux
    port map (
            O => \N__59787\,
            I => \N__59783\
        );

    \I__13269\ : InMux
    port map (
            O => \N__59786\,
            I => \N__59777\
        );

    \I__13268\ : InMux
    port map (
            O => \N__59783\,
            I => \N__59777\
        );

    \I__13267\ : InMux
    port map (
            O => \N__59782\,
            I => \N__59774\
        );

    \I__13266\ : LocalMux
    port map (
            O => \N__59777\,
            I => \N__59771\
        );

    \I__13265\ : LocalMux
    port map (
            O => \N__59774\,
            I => \N__59768\
        );

    \I__13264\ : Odrv4
    port map (
            O => \N__59771\,
            I => \c0.n13_adj_4492\
        );

    \I__13263\ : Odrv12
    port map (
            O => \N__59768\,
            I => \c0.n13_adj_4492\
        );

    \I__13262\ : InMux
    port map (
            O => \N__59763\,
            I => \N__59760\
        );

    \I__13261\ : LocalMux
    port map (
            O => \N__59760\,
            I => \N__59757\
        );

    \I__13260\ : Odrv4
    port map (
            O => \N__59757\,
            I => \c0.n18_adj_4493\
        );

    \I__13259\ : InMux
    port map (
            O => \N__59754\,
            I => \N__59751\
        );

    \I__13258\ : LocalMux
    port map (
            O => \N__59751\,
            I => \N__59748\
        );

    \I__13257\ : Odrv4
    port map (
            O => \N__59748\,
            I => \c0.n22_adj_4498\
        );

    \I__13256\ : CascadeMux
    port map (
            O => \N__59745\,
            I => \c0.n26_adj_4499_cascade_\
        );

    \I__13255\ : InMux
    port map (
            O => \N__59742\,
            I => \N__59739\
        );

    \I__13254\ : LocalMux
    port map (
            O => \N__59739\,
            I => \N__59735\
        );

    \I__13253\ : InMux
    port map (
            O => \N__59738\,
            I => \N__59732\
        );

    \I__13252\ : Span4Mux_v
    port map (
            O => \N__59735\,
            I => \N__59725\
        );

    \I__13251\ : LocalMux
    port map (
            O => \N__59732\,
            I => \N__59725\
        );

    \I__13250\ : CascadeMux
    port map (
            O => \N__59731\,
            I => \N__59721\
        );

    \I__13249\ : InMux
    port map (
            O => \N__59730\,
            I => \N__59717\
        );

    \I__13248\ : Span4Mux_h
    port map (
            O => \N__59725\,
            I => \N__59714\
        );

    \I__13247\ : InMux
    port map (
            O => \N__59724\,
            I => \N__59711\
        );

    \I__13246\ : InMux
    port map (
            O => \N__59721\,
            I => \N__59706\
        );

    \I__13245\ : InMux
    port map (
            O => \N__59720\,
            I => \N__59706\
        );

    \I__13244\ : LocalMux
    port map (
            O => \N__59717\,
            I => \N__59703\
        );

    \I__13243\ : Span4Mux_v
    port map (
            O => \N__59714\,
            I => \N__59699\
        );

    \I__13242\ : LocalMux
    port map (
            O => \N__59711\,
            I => \N__59692\
        );

    \I__13241\ : LocalMux
    port map (
            O => \N__59706\,
            I => \N__59692\
        );

    \I__13240\ : Sp12to4
    port map (
            O => \N__59703\,
            I => \N__59692\
        );

    \I__13239\ : InMux
    port map (
            O => \N__59702\,
            I => \N__59689\
        );

    \I__13238\ : Span4Mux_v
    port map (
            O => \N__59699\,
            I => \N__59686\
        );

    \I__13237\ : Span12Mux_v
    port map (
            O => \N__59692\,
            I => \N__59683\
        );

    \I__13236\ : LocalMux
    port map (
            O => \N__59689\,
            I => \c0.data_in_frame_20_4\
        );

    \I__13235\ : Odrv4
    port map (
            O => \N__59686\,
            I => \c0.data_in_frame_20_4\
        );

    \I__13234\ : Odrv12
    port map (
            O => \N__59683\,
            I => \c0.data_in_frame_20_4\
        );

    \I__13233\ : InMux
    port map (
            O => \N__59676\,
            I => \N__59673\
        );

    \I__13232\ : LocalMux
    port map (
            O => \N__59673\,
            I => \c0.n30_adj_4357\
        );

    \I__13231\ : CascadeMux
    port map (
            O => \N__59670\,
            I => \N__59667\
        );

    \I__13230\ : InMux
    port map (
            O => \N__59667\,
            I => \N__59664\
        );

    \I__13229\ : LocalMux
    port map (
            O => \N__59664\,
            I => \N__59660\
        );

    \I__13228\ : InMux
    port map (
            O => \N__59663\,
            I => \N__59657\
        );

    \I__13227\ : Span4Mux_h
    port map (
            O => \N__59660\,
            I => \N__59654\
        );

    \I__13226\ : LocalMux
    port map (
            O => \N__59657\,
            I => \N__59651\
        );

    \I__13225\ : Span4Mux_v
    port map (
            O => \N__59654\,
            I => \N__59648\
        );

    \I__13224\ : Span4Mux_h
    port map (
            O => \N__59651\,
            I => \N__59645\
        );

    \I__13223\ : Odrv4
    port map (
            O => \N__59648\,
            I => \c0.n22334\
        );

    \I__13222\ : Odrv4
    port map (
            O => \N__59645\,
            I => \c0.n22334\
        );

    \I__13221\ : CascadeMux
    port map (
            O => \N__59640\,
            I => \N__59637\
        );

    \I__13220\ : InMux
    port map (
            O => \N__59637\,
            I => \N__59633\
        );

    \I__13219\ : CascadeMux
    port map (
            O => \N__59636\,
            I => \N__59630\
        );

    \I__13218\ : LocalMux
    port map (
            O => \N__59633\,
            I => \N__59625\
        );

    \I__13217\ : InMux
    port map (
            O => \N__59630\,
            I => \N__59622\
        );

    \I__13216\ : CascadeMux
    port map (
            O => \N__59629\,
            I => \N__59619\
        );

    \I__13215\ : CascadeMux
    port map (
            O => \N__59628\,
            I => \N__59616\
        );

    \I__13214\ : Span4Mux_v
    port map (
            O => \N__59625\,
            I => \N__59613\
        );

    \I__13213\ : LocalMux
    port map (
            O => \N__59622\,
            I => \N__59610\
        );

    \I__13212\ : InMux
    port map (
            O => \N__59619\,
            I => \N__59607\
        );

    \I__13211\ : InMux
    port map (
            O => \N__59616\,
            I => \N__59604\
        );

    \I__13210\ : Span4Mux_h
    port map (
            O => \N__59613\,
            I => \N__59601\
        );

    \I__13209\ : Span4Mux_v
    port map (
            O => \N__59610\,
            I => \N__59598\
        );

    \I__13208\ : LocalMux
    port map (
            O => \N__59607\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13207\ : LocalMux
    port map (
            O => \N__59604\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13206\ : Odrv4
    port map (
            O => \N__59601\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13205\ : Odrv4
    port map (
            O => \N__59598\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13204\ : InMux
    port map (
            O => \N__59589\,
            I => \N__59582\
        );

    \I__13203\ : InMux
    port map (
            O => \N__59588\,
            I => \N__59582\
        );

    \I__13202\ : CascadeMux
    port map (
            O => \N__59587\,
            I => \N__59579\
        );

    \I__13201\ : LocalMux
    port map (
            O => \N__59582\,
            I => \N__59575\
        );

    \I__13200\ : InMux
    port map (
            O => \N__59579\,
            I => \N__59570\
        );

    \I__13199\ : InMux
    port map (
            O => \N__59578\,
            I => \N__59570\
        );

    \I__13198\ : Span4Mux_h
    port map (
            O => \N__59575\,
            I => \N__59567\
        );

    \I__13197\ : LocalMux
    port map (
            O => \N__59570\,
            I => \c0.data_in_frame_24_3\
        );

    \I__13196\ : Odrv4
    port map (
            O => \N__59567\,
            I => \c0.data_in_frame_24_3\
        );

    \I__13195\ : InMux
    port map (
            O => \N__59562\,
            I => \N__59558\
        );

    \I__13194\ : InMux
    port map (
            O => \N__59561\,
            I => \N__59553\
        );

    \I__13193\ : LocalMux
    port map (
            O => \N__59558\,
            I => \N__59550\
        );

    \I__13192\ : InMux
    port map (
            O => \N__59557\,
            I => \N__59545\
        );

    \I__13191\ : InMux
    port map (
            O => \N__59556\,
            I => \N__59545\
        );

    \I__13190\ : LocalMux
    port map (
            O => \N__59553\,
            I => \N__59542\
        );

    \I__13189\ : Span4Mux_h
    port map (
            O => \N__59550\,
            I => \N__59539\
        );

    \I__13188\ : LocalMux
    port map (
            O => \N__59545\,
            I => \c0.n24547\
        );

    \I__13187\ : Odrv4
    port map (
            O => \N__59542\,
            I => \c0.n24547\
        );

    \I__13186\ : Odrv4
    port map (
            O => \N__59539\,
            I => \c0.n24547\
        );

    \I__13185\ : CascadeMux
    port map (
            O => \N__59532\,
            I => \N__59529\
        );

    \I__13184\ : InMux
    port map (
            O => \N__59529\,
            I => \N__59526\
        );

    \I__13183\ : LocalMux
    port map (
            O => \N__59526\,
            I => \N__59521\
        );

    \I__13182\ : InMux
    port map (
            O => \N__59525\,
            I => \N__59516\
        );

    \I__13181\ : InMux
    port map (
            O => \N__59524\,
            I => \N__59516\
        );

    \I__13180\ : Span4Mux_v
    port map (
            O => \N__59521\,
            I => \N__59513\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__59516\,
            I => \c0.n21353\
        );

    \I__13178\ : Odrv4
    port map (
            O => \N__59513\,
            I => \c0.n21353\
        );

    \I__13177\ : CascadeMux
    port map (
            O => \N__59508\,
            I => \c0.n66_cascade_\
        );

    \I__13176\ : InMux
    port map (
            O => \N__59505\,
            I => \N__59502\
        );

    \I__13175\ : LocalMux
    port map (
            O => \N__59502\,
            I => \c0.n75\
        );

    \I__13174\ : InMux
    port map (
            O => \N__59499\,
            I => \N__59496\
        );

    \I__13173\ : LocalMux
    port map (
            O => \N__59496\,
            I => \c0.n46_adj_4461\
        );

    \I__13172\ : InMux
    port map (
            O => \N__59493\,
            I => \N__59490\
        );

    \I__13171\ : LocalMux
    port map (
            O => \N__59490\,
            I => \N__59487\
        );

    \I__13170\ : Odrv12
    port map (
            O => \N__59487\,
            I => \c0.n4_adj_4347\
        );

    \I__13169\ : InMux
    port map (
            O => \N__59484\,
            I => \N__59481\
        );

    \I__13168\ : LocalMux
    port map (
            O => \N__59481\,
            I => \N__59476\
        );

    \I__13167\ : InMux
    port map (
            O => \N__59480\,
            I => \N__59471\
        );

    \I__13166\ : InMux
    port map (
            O => \N__59479\,
            I => \N__59471\
        );

    \I__13165\ : Span4Mux_h
    port map (
            O => \N__59476\,
            I => \N__59468\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__59471\,
            I => \c0.data_in_frame_23_4\
        );

    \I__13163\ : Odrv4
    port map (
            O => \N__59468\,
            I => \c0.data_in_frame_23_4\
        );

    \I__13162\ : CascadeMux
    port map (
            O => \N__59463\,
            I => \c0.n4_adj_4347_cascade_\
        );

    \I__13161\ : CascadeMux
    port map (
            O => \N__59460\,
            I => \N__59457\
        );

    \I__13160\ : InMux
    port map (
            O => \N__59457\,
            I => \N__59453\
        );

    \I__13159\ : InMux
    port map (
            O => \N__59456\,
            I => \N__59450\
        );

    \I__13158\ : LocalMux
    port map (
            O => \N__59453\,
            I => \c0.data_in_frame_23_1\
        );

    \I__13157\ : LocalMux
    port map (
            O => \N__59450\,
            I => \c0.data_in_frame_23_1\
        );

    \I__13156\ : CascadeMux
    port map (
            O => \N__59445\,
            I => \c0.n30_adj_4357_cascade_\
        );

    \I__13155\ : InMux
    port map (
            O => \N__59442\,
            I => \N__59435\
        );

    \I__13154\ : InMux
    port map (
            O => \N__59441\,
            I => \N__59435\
        );

    \I__13153\ : InMux
    port map (
            O => \N__59440\,
            I => \N__59430\
        );

    \I__13152\ : LocalMux
    port map (
            O => \N__59435\,
            I => \N__59427\
        );

    \I__13151\ : InMux
    port map (
            O => \N__59434\,
            I => \N__59424\
        );

    \I__13150\ : InMux
    port map (
            O => \N__59433\,
            I => \N__59421\
        );

    \I__13149\ : LocalMux
    port map (
            O => \N__59430\,
            I => \N__59418\
        );

    \I__13148\ : Span4Mux_h
    port map (
            O => \N__59427\,
            I => \N__59415\
        );

    \I__13147\ : LocalMux
    port map (
            O => \N__59424\,
            I => \N__59412\
        );

    \I__13146\ : LocalMux
    port map (
            O => \N__59421\,
            I => \c0.n14_adj_4356\
        );

    \I__13145\ : Odrv4
    port map (
            O => \N__59418\,
            I => \c0.n14_adj_4356\
        );

    \I__13144\ : Odrv4
    port map (
            O => \N__59415\,
            I => \c0.n14_adj_4356\
        );

    \I__13143\ : Odrv4
    port map (
            O => \N__59412\,
            I => \c0.n14_adj_4356\
        );

    \I__13142\ : InMux
    port map (
            O => \N__59403\,
            I => \N__59400\
        );

    \I__13141\ : LocalMux
    port map (
            O => \N__59400\,
            I => \c0.n40_adj_4359\
        );

    \I__13140\ : CascadeMux
    port map (
            O => \N__59397\,
            I => \c0.n42_adj_4358_cascade_\
        );

    \I__13139\ : InMux
    port map (
            O => \N__59394\,
            I => \N__59391\
        );

    \I__13138\ : LocalMux
    port map (
            O => \N__59391\,
            I => \N__59388\
        );

    \I__13137\ : Odrv12
    port map (
            O => \N__59388\,
            I => \c0.n41_adj_4360\
        );

    \I__13136\ : InMux
    port map (
            O => \N__59385\,
            I => \N__59382\
        );

    \I__13135\ : LocalMux
    port map (
            O => \N__59382\,
            I => \c0.n37_adj_4458\
        );

    \I__13134\ : CascadeMux
    port map (
            O => \N__59379\,
            I => \c0.n34_adj_4361_cascade_\
        );

    \I__13133\ : InMux
    port map (
            O => \N__59376\,
            I => \N__59373\
        );

    \I__13132\ : LocalMux
    port map (
            O => \N__59373\,
            I => \c0.n14148\
        );

    \I__13131\ : InMux
    port map (
            O => \N__59370\,
            I => \N__59367\
        );

    \I__13130\ : LocalMux
    port map (
            O => \N__59367\,
            I => \N__59363\
        );

    \I__13129\ : InMux
    port map (
            O => \N__59366\,
            I => \N__59360\
        );

    \I__13128\ : Odrv12
    port map (
            O => \N__59363\,
            I => \c0.n9_adj_4208\
        );

    \I__13127\ : LocalMux
    port map (
            O => \N__59360\,
            I => \c0.n9_adj_4208\
        );

    \I__13126\ : CascadeMux
    port map (
            O => \N__59355\,
            I => \c0.n6_adj_4587_cascade_\
        );

    \I__13125\ : InMux
    port map (
            O => \N__59352\,
            I => \N__59349\
        );

    \I__13124\ : LocalMux
    port map (
            O => \N__59349\,
            I => \N__59345\
        );

    \I__13123\ : InMux
    port map (
            O => \N__59348\,
            I => \N__59342\
        );

    \I__13122\ : Span4Mux_h
    port map (
            O => \N__59345\,
            I => \N__59339\
        );

    \I__13121\ : LocalMux
    port map (
            O => \N__59342\,
            I => \c0.n13461\
        );

    \I__13120\ : Odrv4
    port map (
            O => \N__59339\,
            I => \c0.n13461\
        );

    \I__13119\ : CascadeMux
    port map (
            O => \N__59334\,
            I => \N__59330\
        );

    \I__13118\ : InMux
    port map (
            O => \N__59333\,
            I => \N__59326\
        );

    \I__13117\ : InMux
    port map (
            O => \N__59330\,
            I => \N__59321\
        );

    \I__13116\ : InMux
    port map (
            O => \N__59329\,
            I => \N__59321\
        );

    \I__13115\ : LocalMux
    port map (
            O => \N__59326\,
            I => \N__59316\
        );

    \I__13114\ : LocalMux
    port map (
            O => \N__59321\,
            I => \N__59316\
        );

    \I__13113\ : Sp12to4
    port map (
            O => \N__59316\,
            I => \N__59313\
        );

    \I__13112\ : Odrv12
    port map (
            O => \N__59313\,
            I => \c0.n13756\
        );

    \I__13111\ : CascadeMux
    port map (
            O => \N__59310\,
            I => \c0.n13461_cascade_\
        );

    \I__13110\ : CascadeMux
    port map (
            O => \N__59307\,
            I => \c0.n6227_cascade_\
        );

    \I__13109\ : InMux
    port map (
            O => \N__59304\,
            I => \N__59301\
        );

    \I__13108\ : LocalMux
    port map (
            O => \N__59301\,
            I => \N__59297\
        );

    \I__13107\ : InMux
    port map (
            O => \N__59300\,
            I => \N__59294\
        );

    \I__13106\ : Span4Mux_v
    port map (
            O => \N__59297\,
            I => \N__59289\
        );

    \I__13105\ : LocalMux
    port map (
            O => \N__59294\,
            I => \N__59289\
        );

    \I__13104\ : Odrv4
    port map (
            O => \N__59289\,
            I => \c0.n22173\
        );

    \I__13103\ : InMux
    port map (
            O => \N__59286\,
            I => \N__59283\
        );

    \I__13102\ : LocalMux
    port map (
            O => \N__59283\,
            I => \N__59277\
        );

    \I__13101\ : InMux
    port map (
            O => \N__59282\,
            I => \N__59270\
        );

    \I__13100\ : InMux
    port map (
            O => \N__59281\,
            I => \N__59270\
        );

    \I__13099\ : InMux
    port map (
            O => \N__59280\,
            I => \N__59270\
        );

    \I__13098\ : Odrv12
    port map (
            O => \N__59277\,
            I => \c0.n19_adj_4291\
        );

    \I__13097\ : LocalMux
    port map (
            O => \N__59270\,
            I => \c0.n19_adj_4291\
        );

    \I__13096\ : CascadeMux
    port map (
            O => \N__59265\,
            I => \N__59262\
        );

    \I__13095\ : InMux
    port map (
            O => \N__59262\,
            I => \N__59256\
        );

    \I__13094\ : InMux
    port map (
            O => \N__59261\,
            I => \N__59253\
        );

    \I__13093\ : InMux
    port map (
            O => \N__59260\,
            I => \N__59250\
        );

    \I__13092\ : InMux
    port map (
            O => \N__59259\,
            I => \N__59247\
        );

    \I__13091\ : LocalMux
    port map (
            O => \N__59256\,
            I => \N__59244\
        );

    \I__13090\ : LocalMux
    port map (
            O => \N__59253\,
            I => \N__59240\
        );

    \I__13089\ : LocalMux
    port map (
            O => \N__59250\,
            I => \N__59237\
        );

    \I__13088\ : LocalMux
    port map (
            O => \N__59247\,
            I => \N__59232\
        );

    \I__13087\ : Span4Mux_h
    port map (
            O => \N__59244\,
            I => \N__59232\
        );

    \I__13086\ : CascadeMux
    port map (
            O => \N__59243\,
            I => \N__59228\
        );

    \I__13085\ : Span4Mux_v
    port map (
            O => \N__59240\,
            I => \N__59225\
        );

    \I__13084\ : Span4Mux_h
    port map (
            O => \N__59237\,
            I => \N__59220\
        );

    \I__13083\ : Span4Mux_v
    port map (
            O => \N__59232\,
            I => \N__59220\
        );

    \I__13082\ : InMux
    port map (
            O => \N__59231\,
            I => \N__59215\
        );

    \I__13081\ : InMux
    port map (
            O => \N__59228\,
            I => \N__59215\
        );

    \I__13080\ : Odrv4
    port map (
            O => \N__59225\,
            I => data_in_frame_14_6
        );

    \I__13079\ : Odrv4
    port map (
            O => \N__59220\,
            I => data_in_frame_14_6
        );

    \I__13078\ : LocalMux
    port map (
            O => \N__59215\,
            I => data_in_frame_14_6
        );

    \I__13077\ : InMux
    port map (
            O => \N__59208\,
            I => \N__59202\
        );

    \I__13076\ : InMux
    port map (
            O => \N__59207\,
            I => \N__59199\
        );

    \I__13075\ : InMux
    port map (
            O => \N__59206\,
            I => \N__59194\
        );

    \I__13074\ : InMux
    port map (
            O => \N__59205\,
            I => \N__59191\
        );

    \I__13073\ : LocalMux
    port map (
            O => \N__59202\,
            I => \N__59187\
        );

    \I__13072\ : LocalMux
    port map (
            O => \N__59199\,
            I => \N__59184\
        );

    \I__13071\ : InMux
    port map (
            O => \N__59198\,
            I => \N__59179\
        );

    \I__13070\ : InMux
    port map (
            O => \N__59197\,
            I => \N__59179\
        );

    \I__13069\ : LocalMux
    port map (
            O => \N__59194\,
            I => \N__59176\
        );

    \I__13068\ : LocalMux
    port map (
            O => \N__59191\,
            I => \N__59173\
        );

    \I__13067\ : InMux
    port map (
            O => \N__59190\,
            I => \N__59170\
        );

    \I__13066\ : Span4Mux_v
    port map (
            O => \N__59187\,
            I => \N__59165\
        );

    \I__13065\ : Span4Mux_h
    port map (
            O => \N__59184\,
            I => \N__59165\
        );

    \I__13064\ : LocalMux
    port map (
            O => \N__59179\,
            I => \N__59162\
        );

    \I__13063\ : Span4Mux_h
    port map (
            O => \N__59176\,
            I => \N__59157\
        );

    \I__13062\ : Span4Mux_h
    port map (
            O => \N__59173\,
            I => \N__59157\
        );

    \I__13061\ : LocalMux
    port map (
            O => \N__59170\,
            I => \N__59154\
        );

    \I__13060\ : Span4Mux_v
    port map (
            O => \N__59165\,
            I => \N__59149\
        );

    \I__13059\ : Span4Mux_h
    port map (
            O => \N__59162\,
            I => \N__59149\
        );

    \I__13058\ : Span4Mux_v
    port map (
            O => \N__59157\,
            I => \N__59143\
        );

    \I__13057\ : Span4Mux_h
    port map (
            O => \N__59154\,
            I => \N__59143\
        );

    \I__13056\ : Span4Mux_v
    port map (
            O => \N__59149\,
            I => \N__59140\
        );

    \I__13055\ : InMux
    port map (
            O => \N__59148\,
            I => \N__59137\
        );

    \I__13054\ : Odrv4
    port map (
            O => \N__59143\,
            I => n22118
        );

    \I__13053\ : Odrv4
    port map (
            O => \N__59140\,
            I => n22118
        );

    \I__13052\ : LocalMux
    port map (
            O => \N__59137\,
            I => n22118
        );

    \I__13051\ : InMux
    port map (
            O => \N__59130\,
            I => \N__59126\
        );

    \I__13050\ : InMux
    port map (
            O => \N__59129\,
            I => \N__59122\
        );

    \I__13049\ : LocalMux
    port map (
            O => \N__59126\,
            I => \N__59119\
        );

    \I__13048\ : InMux
    port map (
            O => \N__59125\,
            I => \N__59116\
        );

    \I__13047\ : LocalMux
    port map (
            O => \N__59122\,
            I => \c0.data_in_frame_19_3\
        );

    \I__13046\ : Odrv4
    port map (
            O => \N__59119\,
            I => \c0.data_in_frame_19_3\
        );

    \I__13045\ : LocalMux
    port map (
            O => \N__59116\,
            I => \c0.data_in_frame_19_3\
        );

    \I__13044\ : InMux
    port map (
            O => \N__59109\,
            I => \N__59106\
        );

    \I__13043\ : LocalMux
    port map (
            O => \N__59106\,
            I => \N__59102\
        );

    \I__13042\ : InMux
    port map (
            O => \N__59105\,
            I => \N__59099\
        );

    \I__13041\ : Span4Mux_v
    port map (
            O => \N__59102\,
            I => \N__59096\
        );

    \I__13040\ : LocalMux
    port map (
            O => \N__59099\,
            I => \N__59093\
        );

    \I__13039\ : Odrv4
    port map (
            O => \N__59096\,
            I => \c0.n14088\
        );

    \I__13038\ : Odrv12
    port map (
            O => \N__59093\,
            I => \c0.n14088\
        );

    \I__13037\ : InMux
    port map (
            O => \N__59088\,
            I => \N__59085\
        );

    \I__13036\ : LocalMux
    port map (
            O => \N__59085\,
            I => \c0.n23300\
        );

    \I__13035\ : InMux
    port map (
            O => \N__59082\,
            I => \N__59078\
        );

    \I__13034\ : InMux
    port map (
            O => \N__59081\,
            I => \N__59075\
        );

    \I__13033\ : LocalMux
    port map (
            O => \N__59078\,
            I => \N__59072\
        );

    \I__13032\ : LocalMux
    port map (
            O => \N__59075\,
            I => \N__59069\
        );

    \I__13031\ : Span4Mux_v
    port map (
            O => \N__59072\,
            I => \N__59064\
        );

    \I__13030\ : Span4Mux_v
    port map (
            O => \N__59069\,
            I => \N__59064\
        );

    \I__13029\ : Span4Mux_h
    port map (
            O => \N__59064\,
            I => \N__59061\
        );

    \I__13028\ : Odrv4
    port map (
            O => \N__59061\,
            I => \c0.n6_adj_4577\
        );

    \I__13027\ : CascadeMux
    port map (
            O => \N__59058\,
            I => \N__59054\
        );

    \I__13026\ : InMux
    port map (
            O => \N__59057\,
            I => \N__59050\
        );

    \I__13025\ : InMux
    port map (
            O => \N__59054\,
            I => \N__59047\
        );

    \I__13024\ : InMux
    port map (
            O => \N__59053\,
            I => \N__59044\
        );

    \I__13023\ : LocalMux
    port map (
            O => \N__59050\,
            I => \N__59039\
        );

    \I__13022\ : LocalMux
    port map (
            O => \N__59047\,
            I => \N__59039\
        );

    \I__13021\ : LocalMux
    port map (
            O => \N__59044\,
            I => \c0.n22662\
        );

    \I__13020\ : Odrv12
    port map (
            O => \N__59039\,
            I => \c0.n22662\
        );

    \I__13019\ : CascadeMux
    port map (
            O => \N__59034\,
            I => \c0.n23300_cascade_\
        );

    \I__13018\ : InMux
    port map (
            O => \N__59031\,
            I => \N__59028\
        );

    \I__13017\ : LocalMux
    port map (
            O => \N__59028\,
            I => \c0.n21_adj_4594\
        );

    \I__13016\ : InMux
    port map (
            O => \N__59025\,
            I => \N__59022\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__59022\,
            I => \N__59019\
        );

    \I__13014\ : Span4Mux_v
    port map (
            O => \N__59019\,
            I => \N__59015\
        );

    \I__13013\ : InMux
    port map (
            O => \N__59018\,
            I => \N__59012\
        );

    \I__13012\ : Span4Mux_h
    port map (
            O => \N__59015\,
            I => \N__59005\
        );

    \I__13011\ : LocalMux
    port map (
            O => \N__59012\,
            I => \N__59005\
        );

    \I__13010\ : CascadeMux
    port map (
            O => \N__59011\,
            I => \N__59002\
        );

    \I__13009\ : InMux
    port map (
            O => \N__59010\,
            I => \N__58998\
        );

    \I__13008\ : Span4Mux_v
    port map (
            O => \N__59005\,
            I => \N__58995\
        );

    \I__13007\ : InMux
    port map (
            O => \N__59002\,
            I => \N__58990\
        );

    \I__13006\ : InMux
    port map (
            O => \N__59001\,
            I => \N__58990\
        );

    \I__13005\ : LocalMux
    port map (
            O => \N__58998\,
            I => \c0.data_in_frame_12_4\
        );

    \I__13004\ : Odrv4
    port map (
            O => \N__58995\,
            I => \c0.data_in_frame_12_4\
        );

    \I__13003\ : LocalMux
    port map (
            O => \N__58990\,
            I => \c0.data_in_frame_12_4\
        );

    \I__13002\ : CascadeMux
    port map (
            O => \N__58983\,
            I => \c0.n4_adj_4658_cascade_\
        );

    \I__13001\ : InMux
    port map (
            O => \N__58980\,
            I => \N__58974\
        );

    \I__13000\ : InMux
    port map (
            O => \N__58979\,
            I => \N__58974\
        );

    \I__12999\ : LocalMux
    port map (
            O => \N__58974\,
            I => \N__58971\
        );

    \I__12998\ : Span4Mux_v
    port map (
            O => \N__58971\,
            I => \N__58968\
        );

    \I__12997\ : Span4Mux_h
    port map (
            O => \N__58968\,
            I => \N__58963\
        );

    \I__12996\ : InMux
    port map (
            O => \N__58967\,
            I => \N__58960\
        );

    \I__12995\ : InMux
    port map (
            O => \N__58966\,
            I => \N__58957\
        );

    \I__12994\ : Span4Mux_v
    port map (
            O => \N__58963\,
            I => \N__58952\
        );

    \I__12993\ : LocalMux
    port map (
            O => \N__58960\,
            I => \N__58952\
        );

    \I__12992\ : LocalMux
    port map (
            O => \N__58957\,
            I => \N__58949\
        );

    \I__12991\ : Span4Mux_v
    port map (
            O => \N__58952\,
            I => \N__58946\
        );

    \I__12990\ : Span12Mux_h
    port map (
            O => \N__58949\,
            I => \N__58943\
        );

    \I__12989\ : Odrv4
    port map (
            O => \N__58946\,
            I => \c0.n24433\
        );

    \I__12988\ : Odrv12
    port map (
            O => \N__58943\,
            I => \c0.n24433\
        );

    \I__12987\ : InMux
    port map (
            O => \N__58938\,
            I => \N__58934\
        );

    \I__12986\ : CascadeMux
    port map (
            O => \N__58937\,
            I => \N__58931\
        );

    \I__12985\ : LocalMux
    port map (
            O => \N__58934\,
            I => \N__58927\
        );

    \I__12984\ : InMux
    port map (
            O => \N__58931\,
            I => \N__58924\
        );

    \I__12983\ : CascadeMux
    port map (
            O => \N__58930\,
            I => \N__58921\
        );

    \I__12982\ : Span4Mux_h
    port map (
            O => \N__58927\,
            I => \N__58918\
        );

    \I__12981\ : LocalMux
    port map (
            O => \N__58924\,
            I => \N__58915\
        );

    \I__12980\ : InMux
    port map (
            O => \N__58921\,
            I => \N__58912\
        );

    \I__12979\ : Span4Mux_h
    port map (
            O => \N__58918\,
            I => \N__58907\
        );

    \I__12978\ : Span4Mux_v
    port map (
            O => \N__58915\,
            I => \N__58907\
        );

    \I__12977\ : LocalMux
    port map (
            O => \N__58912\,
            I => \c0.data_in_frame_16_6\
        );

    \I__12976\ : Odrv4
    port map (
            O => \N__58907\,
            I => \c0.data_in_frame_16_6\
        );

    \I__12975\ : CascadeMux
    port map (
            O => \N__58902\,
            I => \c0.n12_adj_4682_cascade_\
        );

    \I__12974\ : InMux
    port map (
            O => \N__58899\,
            I => \N__58896\
        );

    \I__12973\ : LocalMux
    port map (
            O => \N__58896\,
            I => \N__58893\
        );

    \I__12972\ : Span4Mux_h
    port map (
            O => \N__58893\,
            I => \N__58887\
        );

    \I__12971\ : InMux
    port map (
            O => \N__58892\,
            I => \N__58884\
        );

    \I__12970\ : InMux
    port map (
            O => \N__58891\,
            I => \N__58879\
        );

    \I__12969\ : InMux
    port map (
            O => \N__58890\,
            I => \N__58879\
        );

    \I__12968\ : Odrv4
    port map (
            O => \N__58887\,
            I => \c0.n23390\
        );

    \I__12967\ : LocalMux
    port map (
            O => \N__58884\,
            I => \c0.n23390\
        );

    \I__12966\ : LocalMux
    port map (
            O => \N__58879\,
            I => \c0.n23390\
        );

    \I__12965\ : InMux
    port map (
            O => \N__58872\,
            I => \N__58868\
        );

    \I__12964\ : InMux
    port map (
            O => \N__58871\,
            I => \N__58865\
        );

    \I__12963\ : LocalMux
    port map (
            O => \N__58868\,
            I => \N__58862\
        );

    \I__12962\ : LocalMux
    port map (
            O => \N__58865\,
            I => \N__58859\
        );

    \I__12961\ : Odrv12
    port map (
            O => \N__58862\,
            I => \c0.n22249\
        );

    \I__12960\ : Odrv12
    port map (
            O => \N__58859\,
            I => \c0.n22249\
        );

    \I__12959\ : InMux
    port map (
            O => \N__58854\,
            I => \N__58851\
        );

    \I__12958\ : LocalMux
    port map (
            O => \N__58851\,
            I => \c0.n10_adj_4315\
        );

    \I__12957\ : CascadeMux
    port map (
            O => \N__58848\,
            I => \N__58844\
        );

    \I__12956\ : InMux
    port map (
            O => \N__58847\,
            I => \N__58836\
        );

    \I__12955\ : InMux
    port map (
            O => \N__58844\,
            I => \N__58836\
        );

    \I__12954\ : InMux
    port map (
            O => \N__58843\,
            I => \N__58836\
        );

    \I__12953\ : LocalMux
    port map (
            O => \N__58836\,
            I => \c0.n24534\
        );

    \I__12952\ : InMux
    port map (
            O => \N__58833\,
            I => \N__58830\
        );

    \I__12951\ : LocalMux
    port map (
            O => \N__58830\,
            I => \N__58825\
        );

    \I__12950\ : CascadeMux
    port map (
            O => \N__58829\,
            I => \N__58822\
        );

    \I__12949\ : InMux
    port map (
            O => \N__58828\,
            I => \N__58818\
        );

    \I__12948\ : Span4Mux_h
    port map (
            O => \N__58825\,
            I => \N__58815\
        );

    \I__12947\ : InMux
    port map (
            O => \N__58822\,
            I => \N__58810\
        );

    \I__12946\ : InMux
    port map (
            O => \N__58821\,
            I => \N__58810\
        );

    \I__12945\ : LocalMux
    port map (
            O => \N__58818\,
            I => \c0.data_in_frame_17_3\
        );

    \I__12944\ : Odrv4
    port map (
            O => \N__58815\,
            I => \c0.data_in_frame_17_3\
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__58810\,
            I => \c0.data_in_frame_17_3\
        );

    \I__12942\ : InMux
    port map (
            O => \N__58803\,
            I => \N__58800\
        );

    \I__12941\ : LocalMux
    port map (
            O => \N__58800\,
            I => \c0.n4_adj_4345\
        );

    \I__12940\ : CascadeMux
    port map (
            O => \N__58797\,
            I => \c0.n24534_cascade_\
        );

    \I__12939\ : InMux
    port map (
            O => \N__58794\,
            I => \N__58791\
        );

    \I__12938\ : LocalMux
    port map (
            O => \N__58791\,
            I => \N__58788\
        );

    \I__12937\ : Span4Mux_h
    port map (
            O => \N__58788\,
            I => \N__58785\
        );

    \I__12936\ : Odrv4
    port map (
            O => \N__58785\,
            I => \c0.n12_adj_4346\
        );

    \I__12935\ : CascadeMux
    port map (
            O => \N__58782\,
            I => \N__58779\
        );

    \I__12934\ : InMux
    port map (
            O => \N__58779\,
            I => \N__58768\
        );

    \I__12933\ : InMux
    port map (
            O => \N__58778\,
            I => \N__58768\
        );

    \I__12932\ : InMux
    port map (
            O => \N__58777\,
            I => \N__58768\
        );

    \I__12931\ : InMux
    port map (
            O => \N__58776\,
            I => \N__58764\
        );

    \I__12930\ : InMux
    port map (
            O => \N__58775\,
            I => \N__58761\
        );

    \I__12929\ : LocalMux
    port map (
            O => \N__58768\,
            I => \N__58758\
        );

    \I__12928\ : InMux
    port map (
            O => \N__58767\,
            I => \N__58755\
        );

    \I__12927\ : LocalMux
    port map (
            O => \N__58764\,
            I => \N__58752\
        );

    \I__12926\ : LocalMux
    port map (
            O => \N__58761\,
            I => \N__58748\
        );

    \I__12925\ : Span4Mux_v
    port map (
            O => \N__58758\,
            I => \N__58743\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__58755\,
            I => \N__58743\
        );

    \I__12923\ : Span4Mux_v
    port map (
            O => \N__58752\,
            I => \N__58740\
        );

    \I__12922\ : InMux
    port map (
            O => \N__58751\,
            I => \N__58737\
        );

    \I__12921\ : Span4Mux_v
    port map (
            O => \N__58748\,
            I => \N__58732\
        );

    \I__12920\ : Span4Mux_h
    port map (
            O => \N__58743\,
            I => \N__58732\
        );

    \I__12919\ : Odrv4
    port map (
            O => \N__58740\,
            I => \c0.n13329\
        );

    \I__12918\ : LocalMux
    port map (
            O => \N__58737\,
            I => \c0.n13329\
        );

    \I__12917\ : Odrv4
    port map (
            O => \N__58732\,
            I => \c0.n13329\
        );

    \I__12916\ : InMux
    port map (
            O => \N__58725\,
            I => \N__58722\
        );

    \I__12915\ : LocalMux
    port map (
            O => \N__58722\,
            I => \c0.n4_adj_4621\
        );

    \I__12914\ : InMux
    port map (
            O => \N__58719\,
            I => \N__58716\
        );

    \I__12913\ : LocalMux
    port map (
            O => \N__58716\,
            I => \N__58712\
        );

    \I__12912\ : InMux
    port map (
            O => \N__58715\,
            I => \N__58709\
        );

    \I__12911\ : Odrv4
    port map (
            O => \N__58712\,
            I => \c0.n12_adj_4500\
        );

    \I__12910\ : LocalMux
    port map (
            O => \N__58709\,
            I => \c0.n12_adj_4500\
        );

    \I__12909\ : CascadeMux
    port map (
            O => \N__58704\,
            I => \c0.n22514_cascade_\
        );

    \I__12908\ : InMux
    port map (
            O => \N__58701\,
            I => \N__58697\
        );

    \I__12907\ : InMux
    port map (
            O => \N__58700\,
            I => \N__58694\
        );

    \I__12906\ : LocalMux
    port map (
            O => \N__58697\,
            I => \c0.data_in_frame_16_1\
        );

    \I__12905\ : LocalMux
    port map (
            O => \N__58694\,
            I => \c0.data_in_frame_16_1\
        );

    \I__12904\ : InMux
    port map (
            O => \N__58689\,
            I => \N__58686\
        );

    \I__12903\ : LocalMux
    port map (
            O => \N__58686\,
            I => \N__58683\
        );

    \I__12902\ : Span4Mux_v
    port map (
            O => \N__58683\,
            I => \N__58680\
        );

    \I__12901\ : Span4Mux_h
    port map (
            O => \N__58680\,
            I => \N__58677\
        );

    \I__12900\ : Odrv4
    port map (
            O => \N__58677\,
            I => \c0.n14_adj_4566\
        );

    \I__12899\ : CascadeMux
    port map (
            O => \N__58674\,
            I => \c0.n14165_cascade_\
        );

    \I__12898\ : CascadeMux
    port map (
            O => \N__58671\,
            I => \N__58666\
        );

    \I__12897\ : CascadeMux
    port map (
            O => \N__58670\,
            I => \N__58663\
        );

    \I__12896\ : InMux
    port map (
            O => \N__58669\,
            I => \N__58659\
        );

    \I__12895\ : InMux
    port map (
            O => \N__58666\,
            I => \N__58656\
        );

    \I__12894\ : InMux
    port map (
            O => \N__58663\,
            I => \N__58651\
        );

    \I__12893\ : InMux
    port map (
            O => \N__58662\,
            I => \N__58651\
        );

    \I__12892\ : LocalMux
    port map (
            O => \N__58659\,
            I => \N__58646\
        );

    \I__12891\ : LocalMux
    port map (
            O => \N__58656\,
            I => \N__58646\
        );

    \I__12890\ : LocalMux
    port map (
            O => \N__58651\,
            I => \N__58643\
        );

    \I__12889\ : Odrv12
    port map (
            O => \N__58646\,
            I => \c0.data_in_frame_17_2\
        );

    \I__12888\ : Odrv4
    port map (
            O => \N__58643\,
            I => \c0.data_in_frame_17_2\
        );

    \I__12887\ : CascadeMux
    port map (
            O => \N__58638\,
            I => \N__58635\
        );

    \I__12886\ : InMux
    port map (
            O => \N__58635\,
            I => \N__58632\
        );

    \I__12885\ : LocalMux
    port map (
            O => \N__58632\,
            I => \N__58629\
        );

    \I__12884\ : Span4Mux_v
    port map (
            O => \N__58629\,
            I => \N__58626\
        );

    \I__12883\ : Odrv4
    port map (
            O => \N__58626\,
            I => \c0.n22_adj_4622\
        );

    \I__12882\ : CascadeMux
    port map (
            O => \N__58623\,
            I => \c0.n22825_cascade_\
        );

    \I__12881\ : InMux
    port map (
            O => \N__58620\,
            I => \N__58615\
        );

    \I__12880\ : InMux
    port map (
            O => \N__58619\,
            I => \N__58611\
        );

    \I__12879\ : InMux
    port map (
            O => \N__58618\,
            I => \N__58608\
        );

    \I__12878\ : LocalMux
    port map (
            O => \N__58615\,
            I => \N__58605\
        );

    \I__12877\ : InMux
    port map (
            O => \N__58614\,
            I => \N__58602\
        );

    \I__12876\ : LocalMux
    port map (
            O => \N__58611\,
            I => \N__58599\
        );

    \I__12875\ : LocalMux
    port map (
            O => \N__58608\,
            I => \N__58594\
        );

    \I__12874\ : Span4Mux_h
    port map (
            O => \N__58605\,
            I => \N__58594\
        );

    \I__12873\ : LocalMux
    port map (
            O => \N__58602\,
            I => data_in_frame_14_0
        );

    \I__12872\ : Odrv12
    port map (
            O => \N__58599\,
            I => data_in_frame_14_0
        );

    \I__12871\ : Odrv4
    port map (
            O => \N__58594\,
            I => data_in_frame_14_0
        );

    \I__12870\ : InMux
    port map (
            O => \N__58587\,
            I => \N__58584\
        );

    \I__12869\ : LocalMux
    port map (
            O => \N__58584\,
            I => \N__58581\
        );

    \I__12868\ : Span4Mux_h
    port map (
            O => \N__58581\,
            I => \N__58578\
        );

    \I__12867\ : Span4Mux_h
    port map (
            O => \N__58578\,
            I => \N__58575\
        );

    \I__12866\ : Odrv4
    port map (
            O => \N__58575\,
            I => \c0.n136\
        );

    \I__12865\ : CascadeMux
    port map (
            O => \N__58572\,
            I => \c0.n22751_cascade_\
        );

    \I__12864\ : InMux
    port map (
            O => \N__58569\,
            I => \N__58566\
        );

    \I__12863\ : LocalMux
    port map (
            O => \N__58566\,
            I => \N__58563\
        );

    \I__12862\ : Odrv4
    port map (
            O => \N__58563\,
            I => \c0.n107\
        );

    \I__12861\ : InMux
    port map (
            O => \N__58560\,
            I => \N__58557\
        );

    \I__12860\ : LocalMux
    port map (
            O => \N__58557\,
            I => \c0.n149\
        );

    \I__12859\ : InMux
    port map (
            O => \N__58554\,
            I => \N__58551\
        );

    \I__12858\ : LocalMux
    port map (
            O => \N__58551\,
            I => \c0.n140\
        );

    \I__12857\ : InMux
    port map (
            O => \N__58548\,
            I => \N__58545\
        );

    \I__12856\ : LocalMux
    port map (
            O => \N__58545\,
            I => \N__58541\
        );

    \I__12855\ : InMux
    port map (
            O => \N__58544\,
            I => \N__58538\
        );

    \I__12854\ : Span12Mux_h
    port map (
            O => \N__58541\,
            I => \N__58535\
        );

    \I__12853\ : LocalMux
    port map (
            O => \N__58538\,
            I => \N__58532\
        );

    \I__12852\ : Odrv12
    port map (
            O => \N__58535\,
            I => \c0.n22843\
        );

    \I__12851\ : Odrv4
    port map (
            O => \N__58532\,
            I => \c0.n22843\
        );

    \I__12850\ : InMux
    port map (
            O => \N__58527\,
            I => \N__58524\
        );

    \I__12849\ : LocalMux
    port map (
            O => \N__58524\,
            I => \N__58520\
        );

    \I__12848\ : InMux
    port map (
            O => \N__58523\,
            I => \N__58517\
        );

    \I__12847\ : Span4Mux_v
    port map (
            O => \N__58520\,
            I => \N__58514\
        );

    \I__12846\ : LocalMux
    port map (
            O => \N__58517\,
            I => \N__58511\
        );

    \I__12845\ : Span4Mux_h
    port map (
            O => \N__58514\,
            I => \N__58506\
        );

    \I__12844\ : Span4Mux_v
    port map (
            O => \N__58511\,
            I => \N__58506\
        );

    \I__12843\ : Odrv4
    port map (
            O => \N__58506\,
            I => \c0.n22_adj_4245\
        );

    \I__12842\ : CascadeMux
    port map (
            O => \N__58503\,
            I => \c0.n23598_cascade_\
        );

    \I__12841\ : InMux
    port map (
            O => \N__58500\,
            I => \N__58497\
        );

    \I__12840\ : LocalMux
    port map (
            O => \N__58497\,
            I => \N__58493\
        );

    \I__12839\ : InMux
    port map (
            O => \N__58496\,
            I => \N__58490\
        );

    \I__12838\ : Odrv12
    port map (
            O => \N__58493\,
            I => \c0.n23611\
        );

    \I__12837\ : LocalMux
    port map (
            O => \N__58490\,
            I => \c0.n23611\
        );

    \I__12836\ : CascadeMux
    port map (
            O => \N__58485\,
            I => \c0.n9_adj_4208_cascade_\
        );

    \I__12835\ : InMux
    port map (
            O => \N__58482\,
            I => \N__58479\
        );

    \I__12834\ : LocalMux
    port map (
            O => \N__58479\,
            I => \N__58476\
        );

    \I__12833\ : Span4Mux_v
    port map (
            O => \N__58476\,
            I => \N__58473\
        );

    \I__12832\ : Span4Mux_h
    port map (
            O => \N__58473\,
            I => \N__58469\
        );

    \I__12831\ : InMux
    port map (
            O => \N__58472\,
            I => \N__58466\
        );

    \I__12830\ : Odrv4
    port map (
            O => \N__58469\,
            I => \c0.n22304\
        );

    \I__12829\ : LocalMux
    port map (
            O => \N__58466\,
            I => \c0.n22304\
        );

    \I__12828\ : CascadeMux
    port map (
            O => \N__58461\,
            I => \c0.n13892_cascade_\
        );

    \I__12827\ : CascadeMux
    port map (
            O => \N__58458\,
            I => \N__58455\
        );

    \I__12826\ : InMux
    port map (
            O => \N__58455\,
            I => \N__58452\
        );

    \I__12825\ : LocalMux
    port map (
            O => \N__58452\,
            I => \N__58448\
        );

    \I__12824\ : CascadeMux
    port map (
            O => \N__58451\,
            I => \N__58444\
        );

    \I__12823\ : Span4Mux_v
    port map (
            O => \N__58448\,
            I => \N__58441\
        );

    \I__12822\ : InMux
    port map (
            O => \N__58447\,
            I => \N__58438\
        );

    \I__12821\ : InMux
    port map (
            O => \N__58444\,
            I => \N__58435\
        );

    \I__12820\ : Span4Mux_h
    port map (
            O => \N__58441\,
            I => \N__58430\
        );

    \I__12819\ : LocalMux
    port map (
            O => \N__58438\,
            I => \N__58430\
        );

    \I__12818\ : LocalMux
    port map (
            O => \N__58435\,
            I => \c0.data_in_frame_11_6\
        );

    \I__12817\ : Odrv4
    port map (
            O => \N__58430\,
            I => \c0.data_in_frame_11_6\
        );

    \I__12816\ : InMux
    port map (
            O => \N__58425\,
            I => \N__58422\
        );

    \I__12815\ : LocalMux
    port map (
            O => \N__58422\,
            I => \c0.n13892\
        );

    \I__12814\ : InMux
    port map (
            O => \N__58419\,
            I => \N__58416\
        );

    \I__12813\ : LocalMux
    port map (
            O => \N__58416\,
            I => \N__58413\
        );

    \I__12812\ : Odrv12
    port map (
            O => \N__58413\,
            I => \c0.n31\
        );

    \I__12811\ : CascadeMux
    port map (
            O => \N__58410\,
            I => \c0.n31_cascade_\
        );

    \I__12810\ : InMux
    port map (
            O => \N__58407\,
            I => \N__58404\
        );

    \I__12809\ : LocalMux
    port map (
            O => \N__58404\,
            I => \N__58400\
        );

    \I__12808\ : CascadeMux
    port map (
            O => \N__58403\,
            I => \N__58396\
        );

    \I__12807\ : Span4Mux_v
    port map (
            O => \N__58400\,
            I => \N__58392\
        );

    \I__12806\ : InMux
    port map (
            O => \N__58399\,
            I => \N__58387\
        );

    \I__12805\ : InMux
    port map (
            O => \N__58396\,
            I => \N__58387\
        );

    \I__12804\ : InMux
    port map (
            O => \N__58395\,
            I => \N__58384\
        );

    \I__12803\ : Odrv4
    port map (
            O => \N__58392\,
            I => \c0.data_in_frame_10_0\
        );

    \I__12802\ : LocalMux
    port map (
            O => \N__58387\,
            I => \c0.data_in_frame_10_0\
        );

    \I__12801\ : LocalMux
    port map (
            O => \N__58384\,
            I => \c0.data_in_frame_10_0\
        );

    \I__12800\ : InMux
    port map (
            O => \N__58377\,
            I => \N__58374\
        );

    \I__12799\ : LocalMux
    port map (
            O => \N__58374\,
            I => \N__58369\
        );

    \I__12798\ : InMux
    port map (
            O => \N__58373\,
            I => \N__58366\
        );

    \I__12797\ : InMux
    port map (
            O => \N__58372\,
            I => \N__58363\
        );

    \I__12796\ : Span4Mux_v
    port map (
            O => \N__58369\,
            I => \N__58360\
        );

    \I__12795\ : LocalMux
    port map (
            O => \N__58366\,
            I => \N__58355\
        );

    \I__12794\ : LocalMux
    port map (
            O => \N__58363\,
            I => \N__58355\
        );

    \I__12793\ : Odrv4
    port map (
            O => \N__58360\,
            I => \c0.n28\
        );

    \I__12792\ : Odrv12
    port map (
            O => \N__58355\,
            I => \c0.n28\
        );

    \I__12791\ : CascadeMux
    port map (
            O => \N__58350\,
            I => \N__58347\
        );

    \I__12790\ : InMux
    port map (
            O => \N__58347\,
            I => \N__58344\
        );

    \I__12789\ : LocalMux
    port map (
            O => \N__58344\,
            I => \c0.n24\
        );

    \I__12788\ : InMux
    port map (
            O => \N__58341\,
            I => \N__58338\
        );

    \I__12787\ : LocalMux
    port map (
            O => \N__58338\,
            I => \N__58335\
        );

    \I__12786\ : Odrv4
    port map (
            O => \N__58335\,
            I => \c0.n16\
        );

    \I__12785\ : InMux
    port map (
            O => \N__58332\,
            I => \N__58326\
        );

    \I__12784\ : InMux
    port map (
            O => \N__58331\,
            I => \N__58326\
        );

    \I__12783\ : LocalMux
    port map (
            O => \N__58326\,
            I => data_in_frame_14_2
        );

    \I__12782\ : CascadeMux
    port map (
            O => \N__58323\,
            I => \N__58320\
        );

    \I__12781\ : InMux
    port map (
            O => \N__58320\,
            I => \N__58317\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__58317\,
            I => \c0.n8_adj_4673\
        );

    \I__12779\ : InMux
    port map (
            O => \N__58314\,
            I => \N__58308\
        );

    \I__12778\ : InMux
    port map (
            O => \N__58313\,
            I => \N__58308\
        );

    \I__12777\ : LocalMux
    port map (
            O => \N__58308\,
            I => data_in_frame_6_2
        );

    \I__12776\ : InMux
    port map (
            O => \N__58305\,
            I => \N__58301\
        );

    \I__12775\ : CascadeMux
    port map (
            O => \N__58304\,
            I => \N__58298\
        );

    \I__12774\ : LocalMux
    port map (
            O => \N__58301\,
            I => \N__58295\
        );

    \I__12773\ : InMux
    port map (
            O => \N__58298\,
            I => \N__58292\
        );

    \I__12772\ : Span4Mux_v
    port map (
            O => \N__58295\,
            I => \N__58289\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__58292\,
            I => \c0.data_in_frame_13_0\
        );

    \I__12770\ : Odrv4
    port map (
            O => \N__58289\,
            I => \c0.data_in_frame_13_0\
        );

    \I__12769\ : CascadeMux
    port map (
            O => \N__58284\,
            I => \c0.n22205_cascade_\
        );

    \I__12768\ : InMux
    port map (
            O => \N__58281\,
            I => \N__58274\
        );

    \I__12767\ : InMux
    port map (
            O => \N__58280\,
            I => \N__58274\
        );

    \I__12766\ : InMux
    port map (
            O => \N__58279\,
            I => \N__58271\
        );

    \I__12765\ : LocalMux
    port map (
            O => \N__58274\,
            I => \N__58268\
        );

    \I__12764\ : LocalMux
    port map (
            O => \N__58271\,
            I => \c0.n23491\
        );

    \I__12763\ : Odrv4
    port map (
            O => \N__58268\,
            I => \c0.n23491\
        );

    \I__12762\ : InMux
    port map (
            O => \N__58263\,
            I => \N__58260\
        );

    \I__12761\ : LocalMux
    port map (
            O => \N__58260\,
            I => \N__58257\
        );

    \I__12760\ : Span4Mux_h
    port map (
            O => \N__58257\,
            I => \N__58254\
        );

    \I__12759\ : Span4Mux_v
    port map (
            O => \N__58254\,
            I => \N__58250\
        );

    \I__12758\ : InMux
    port map (
            O => \N__58253\,
            I => \N__58247\
        );

    \I__12757\ : Odrv4
    port map (
            O => \N__58250\,
            I => \c0.n17_adj_4224\
        );

    \I__12756\ : LocalMux
    port map (
            O => \N__58247\,
            I => \c0.n17_adj_4224\
        );

    \I__12755\ : InMux
    port map (
            O => \N__58242\,
            I => \N__58239\
        );

    \I__12754\ : LocalMux
    port map (
            O => \N__58239\,
            I => \N__58236\
        );

    \I__12753\ : Span4Mux_v
    port map (
            O => \N__58236\,
            I => \N__58233\
        );

    \I__12752\ : Odrv4
    port map (
            O => \N__58233\,
            I => \c0.n130\
        );

    \I__12751\ : InMux
    port map (
            O => \N__58230\,
            I => \N__58227\
        );

    \I__12750\ : LocalMux
    port map (
            O => \N__58227\,
            I => \N__58224\
        );

    \I__12749\ : Span4Mux_v
    port map (
            O => \N__58224\,
            I => \N__58221\
        );

    \I__12748\ : Span4Mux_h
    port map (
            O => \N__58221\,
            I => \N__58218\
        );

    \I__12747\ : Sp12to4
    port map (
            O => \N__58218\,
            I => \N__58215\
        );

    \I__12746\ : Odrv12
    port map (
            O => \N__58215\,
            I => \c0.n14_adj_4707\
        );

    \I__12745\ : InMux
    port map (
            O => \N__58212\,
            I => \N__58209\
        );

    \I__12744\ : LocalMux
    port map (
            O => \N__58209\,
            I => \N__58206\
        );

    \I__12743\ : Span4Mux_h
    port map (
            O => \N__58206\,
            I => \N__58203\
        );

    \I__12742\ : Odrv4
    port map (
            O => \N__58203\,
            I => \c0.n15_adj_4710\
        );

    \I__12741\ : CascadeMux
    port map (
            O => \N__58200\,
            I => \N__58196\
        );

    \I__12740\ : InMux
    port map (
            O => \N__58199\,
            I => \N__58193\
        );

    \I__12739\ : InMux
    port map (
            O => \N__58196\,
            I => \N__58190\
        );

    \I__12738\ : LocalMux
    port map (
            O => \N__58193\,
            I => \N__58187\
        );

    \I__12737\ : LocalMux
    port map (
            O => \N__58190\,
            I => \N__58184\
        );

    \I__12736\ : Span4Mux_v
    port map (
            O => \N__58187\,
            I => \N__58181\
        );

    \I__12735\ : Span12Mux_v
    port map (
            O => \N__58184\,
            I => \N__58178\
        );

    \I__12734\ : Odrv4
    port map (
            O => \N__58181\,
            I => \c0.n22511\
        );

    \I__12733\ : Odrv12
    port map (
            O => \N__58178\,
            I => \c0.n22511\
        );

    \I__12732\ : CascadeMux
    port map (
            O => \N__58173\,
            I => \N__58170\
        );

    \I__12731\ : InMux
    port map (
            O => \N__58170\,
            I => \N__58166\
        );

    \I__12730\ : InMux
    port map (
            O => \N__58169\,
            I => \N__58163\
        );

    \I__12729\ : LocalMux
    port map (
            O => \N__58166\,
            I => \N__58159\
        );

    \I__12728\ : LocalMux
    port map (
            O => \N__58163\,
            I => \N__58156\
        );

    \I__12727\ : InMux
    port map (
            O => \N__58162\,
            I => \N__58152\
        );

    \I__12726\ : Span4Mux_v
    port map (
            O => \N__58159\,
            I => \N__58147\
        );

    \I__12725\ : Span4Mux_v
    port map (
            O => \N__58156\,
            I => \N__58147\
        );

    \I__12724\ : InMux
    port map (
            O => \N__58155\,
            I => \N__58144\
        );

    \I__12723\ : LocalMux
    port map (
            O => \N__58152\,
            I => \c0.n22_adj_4259\
        );

    \I__12722\ : Odrv4
    port map (
            O => \N__58147\,
            I => \c0.n22_adj_4259\
        );

    \I__12721\ : LocalMux
    port map (
            O => \N__58144\,
            I => \c0.n22_adj_4259\
        );

    \I__12720\ : InMux
    port map (
            O => \N__58137\,
            I => \N__58133\
        );

    \I__12719\ : InMux
    port map (
            O => \N__58136\,
            I => \N__58129\
        );

    \I__12718\ : LocalMux
    port map (
            O => \N__58133\,
            I => \N__58125\
        );

    \I__12717\ : InMux
    port map (
            O => \N__58132\,
            I => \N__58122\
        );

    \I__12716\ : LocalMux
    port map (
            O => \N__58129\,
            I => \N__58119\
        );

    \I__12715\ : InMux
    port map (
            O => \N__58128\,
            I => \N__58116\
        );

    \I__12714\ : Span4Mux_v
    port map (
            O => \N__58125\,
            I => \N__58113\
        );

    \I__12713\ : LocalMux
    port map (
            O => \N__58122\,
            I => \N__58108\
        );

    \I__12712\ : Span4Mux_v
    port map (
            O => \N__58119\,
            I => \N__58108\
        );

    \I__12711\ : LocalMux
    port map (
            O => \N__58116\,
            I => data_in_frame_6_1
        );

    \I__12710\ : Odrv4
    port map (
            O => \N__58113\,
            I => data_in_frame_6_1
        );

    \I__12709\ : Odrv4
    port map (
            O => \N__58108\,
            I => data_in_frame_6_1
        );

    \I__12708\ : CascadeMux
    port map (
            O => \N__58101\,
            I => \c0.n18_adj_4314_cascade_\
        );

    \I__12707\ : InMux
    port map (
            O => \N__58098\,
            I => \N__58094\
        );

    \I__12706\ : InMux
    port map (
            O => \N__58097\,
            I => \N__58091\
        );

    \I__12705\ : LocalMux
    port map (
            O => \N__58094\,
            I => \N__58087\
        );

    \I__12704\ : LocalMux
    port map (
            O => \N__58091\,
            I => \N__58084\
        );

    \I__12703\ : CascadeMux
    port map (
            O => \N__58090\,
            I => \N__58081\
        );

    \I__12702\ : Span4Mux_h
    port map (
            O => \N__58087\,
            I => \N__58075\
        );

    \I__12701\ : Span4Mux_v
    port map (
            O => \N__58084\,
            I => \N__58072\
        );

    \I__12700\ : InMux
    port map (
            O => \N__58081\,
            I => \N__58063\
        );

    \I__12699\ : InMux
    port map (
            O => \N__58080\,
            I => \N__58063\
        );

    \I__12698\ : InMux
    port map (
            O => \N__58079\,
            I => \N__58063\
        );

    \I__12697\ : InMux
    port map (
            O => \N__58078\,
            I => \N__58063\
        );

    \I__12696\ : Odrv4
    port map (
            O => \N__58075\,
            I => \c0.data_in_frame_3_7\
        );

    \I__12695\ : Odrv4
    port map (
            O => \N__58072\,
            I => \c0.data_in_frame_3_7\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__58063\,
            I => \c0.data_in_frame_3_7\
        );

    \I__12693\ : InMux
    port map (
            O => \N__58056\,
            I => \N__58044\
        );

    \I__12692\ : CascadeMux
    port map (
            O => \N__58055\,
            I => \N__58040\
        );

    \I__12691\ : InMux
    port map (
            O => \N__58054\,
            I => \N__58037\
        );

    \I__12690\ : InMux
    port map (
            O => \N__58053\,
            I => \N__58026\
        );

    \I__12689\ : InMux
    port map (
            O => \N__58052\,
            I => \N__58026\
        );

    \I__12688\ : InMux
    port map (
            O => \N__58051\,
            I => \N__58026\
        );

    \I__12687\ : InMux
    port map (
            O => \N__58050\,
            I => \N__58026\
        );

    \I__12686\ : InMux
    port map (
            O => \N__58049\,
            I => \N__58026\
        );

    \I__12685\ : InMux
    port map (
            O => \N__58048\,
            I => \N__58021\
        );

    \I__12684\ : InMux
    port map (
            O => \N__58047\,
            I => \N__58021\
        );

    \I__12683\ : LocalMux
    port map (
            O => \N__58044\,
            I => \N__58018\
        );

    \I__12682\ : InMux
    port map (
            O => \N__58043\,
            I => \N__58015\
        );

    \I__12681\ : InMux
    port map (
            O => \N__58040\,
            I => \N__58009\
        );

    \I__12680\ : LocalMux
    port map (
            O => \N__58037\,
            I => \N__58002\
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__58026\,
            I => \N__58002\
        );

    \I__12678\ : LocalMux
    port map (
            O => \N__58021\,
            I => \N__58002\
        );

    \I__12677\ : Span12Mux_h
    port map (
            O => \N__58018\,
            I => \N__57999\
        );

    \I__12676\ : LocalMux
    port map (
            O => \N__58015\,
            I => \N__57996\
        );

    \I__12675\ : InMux
    port map (
            O => \N__58014\,
            I => \N__57993\
        );

    \I__12674\ : InMux
    port map (
            O => \N__58013\,
            I => \N__57988\
        );

    \I__12673\ : InMux
    port map (
            O => \N__58012\,
            I => \N__57988\
        );

    \I__12672\ : LocalMux
    port map (
            O => \N__58009\,
            I => \N__57983\
        );

    \I__12671\ : Span4Mux_v
    port map (
            O => \N__58002\,
            I => \N__57983\
        );

    \I__12670\ : Odrv12
    port map (
            O => \N__57999\,
            I => data_in_frame_1_6
        );

    \I__12669\ : Odrv4
    port map (
            O => \N__57996\,
            I => data_in_frame_1_6
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__57993\,
            I => data_in_frame_1_6
        );

    \I__12667\ : LocalMux
    port map (
            O => \N__57988\,
            I => data_in_frame_1_6
        );

    \I__12666\ : Odrv4
    port map (
            O => \N__57983\,
            I => data_in_frame_1_6
        );

    \I__12665\ : InMux
    port map (
            O => \N__57972\,
            I => \N__57969\
        );

    \I__12664\ : LocalMux
    port map (
            O => \N__57969\,
            I => \c0.n38_adj_4448\
        );

    \I__12663\ : InMux
    port map (
            O => \N__57966\,
            I => \N__57963\
        );

    \I__12662\ : LocalMux
    port map (
            O => \N__57963\,
            I => \c0.n42_adj_4449\
        );

    \I__12661\ : InMux
    port map (
            O => \N__57960\,
            I => \N__57952\
        );

    \I__12660\ : InMux
    port map (
            O => \N__57959\,
            I => \N__57952\
        );

    \I__12659\ : InMux
    port map (
            O => \N__57958\,
            I => \N__57946\
        );

    \I__12658\ : InMux
    port map (
            O => \N__57957\,
            I => \N__57943\
        );

    \I__12657\ : LocalMux
    port map (
            O => \N__57952\,
            I => \N__57939\
        );

    \I__12656\ : InMux
    port map (
            O => \N__57951\,
            I => \N__57934\
        );

    \I__12655\ : InMux
    port map (
            O => \N__57950\,
            I => \N__57934\
        );

    \I__12654\ : CascadeMux
    port map (
            O => \N__57949\,
            I => \N__57931\
        );

    \I__12653\ : LocalMux
    port map (
            O => \N__57946\,
            I => \N__57925\
        );

    \I__12652\ : LocalMux
    port map (
            O => \N__57943\,
            I => \N__57925\
        );

    \I__12651\ : InMux
    port map (
            O => \N__57942\,
            I => \N__57922\
        );

    \I__12650\ : Span4Mux_v
    port map (
            O => \N__57939\,
            I => \N__57917\
        );

    \I__12649\ : LocalMux
    port map (
            O => \N__57934\,
            I => \N__57917\
        );

    \I__12648\ : InMux
    port map (
            O => \N__57931\,
            I => \N__57912\
        );

    \I__12647\ : InMux
    port map (
            O => \N__57930\,
            I => \N__57912\
        );

    \I__12646\ : Span4Mux_h
    port map (
            O => \N__57925\,
            I => \N__57909\
        );

    \I__12645\ : LocalMux
    port map (
            O => \N__57922\,
            I => \c0.data_in_frame_3_3\
        );

    \I__12644\ : Odrv4
    port map (
            O => \N__57917\,
            I => \c0.data_in_frame_3_3\
        );

    \I__12643\ : LocalMux
    port map (
            O => \N__57912\,
            I => \c0.data_in_frame_3_3\
        );

    \I__12642\ : Odrv4
    port map (
            O => \N__57909\,
            I => \c0.data_in_frame_3_3\
        );

    \I__12641\ : InMux
    port map (
            O => \N__57900\,
            I => \N__57897\
        );

    \I__12640\ : LocalMux
    port map (
            O => \N__57897\,
            I => \N__57894\
        );

    \I__12639\ : Span4Mux_h
    port map (
            O => \N__57894\,
            I => \N__57891\
        );

    \I__12638\ : Odrv4
    port map (
            O => \N__57891\,
            I => \c0.n24_adj_4689\
        );

    \I__12637\ : InMux
    port map (
            O => \N__57888\,
            I => \N__57883\
        );

    \I__12636\ : InMux
    port map (
            O => \N__57887\,
            I => \N__57878\
        );

    \I__12635\ : InMux
    port map (
            O => \N__57886\,
            I => \N__57878\
        );

    \I__12634\ : LocalMux
    port map (
            O => \N__57883\,
            I => \N__57875\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__57878\,
            I => \N__57872\
        );

    \I__12632\ : Span4Mux_h
    port map (
            O => \N__57875\,
            I => \N__57869\
        );

    \I__12631\ : Odrv4
    port map (
            O => \N__57872\,
            I => \c0.n13_adj_4281\
        );

    \I__12630\ : Odrv4
    port map (
            O => \N__57869\,
            I => \c0.n13_adj_4281\
        );

    \I__12629\ : InMux
    port map (
            O => \N__57864\,
            I => \N__57861\
        );

    \I__12628\ : LocalMux
    port map (
            O => \N__57861\,
            I => \N__57858\
        );

    \I__12627\ : Odrv4
    port map (
            O => \N__57858\,
            I => \c0.n102_adj_4445\
        );

    \I__12626\ : InMux
    port map (
            O => \N__57855\,
            I => \N__57852\
        );

    \I__12625\ : LocalMux
    port map (
            O => \N__57852\,
            I => \c0.n101\
        );

    \I__12624\ : InMux
    port map (
            O => \N__57849\,
            I => \N__57846\
        );

    \I__12623\ : LocalMux
    port map (
            O => \N__57846\,
            I => \c0.n103\
        );

    \I__12622\ : InMux
    port map (
            O => \N__57843\,
            I => \N__57840\
        );

    \I__12621\ : LocalMux
    port map (
            O => \N__57840\,
            I => \c0.n98\
        );

    \I__12620\ : InMux
    port map (
            O => \N__57837\,
            I => \N__57834\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__57834\,
            I => \N__57831\
        );

    \I__12618\ : Span4Mux_v
    port map (
            O => \N__57831\,
            I => \N__57828\
        );

    \I__12617\ : Odrv4
    port map (
            O => \N__57828\,
            I => \c0.n97\
        );

    \I__12616\ : CascadeMux
    port map (
            O => \N__57825\,
            I => \c0.n110_cascade_\
        );

    \I__12615\ : InMux
    port map (
            O => \N__57822\,
            I => \N__57819\
        );

    \I__12614\ : LocalMux
    port map (
            O => \N__57819\,
            I => \c0.n24465\
        );

    \I__12613\ : InMux
    port map (
            O => \N__57816\,
            I => \N__57813\
        );

    \I__12612\ : LocalMux
    port map (
            O => \N__57813\,
            I => \N__57810\
        );

    \I__12611\ : Span4Mux_v
    port map (
            O => \N__57810\,
            I => \N__57807\
        );

    \I__12610\ : Span4Mux_h
    port map (
            O => \N__57807\,
            I => \N__57804\
        );

    \I__12609\ : Odrv4
    port map (
            O => \N__57804\,
            I => \c0.data_out_frame_0__7__N_2579\
        );

    \I__12608\ : InMux
    port map (
            O => \N__57801\,
            I => \N__57797\
        );

    \I__12607\ : CascadeMux
    port map (
            O => \N__57800\,
            I => \N__57794\
        );

    \I__12606\ : LocalMux
    port map (
            O => \N__57797\,
            I => \N__57791\
        );

    \I__12605\ : InMux
    port map (
            O => \N__57794\,
            I => \N__57788\
        );

    \I__12604\ : Odrv4
    port map (
            O => \N__57791\,
            I => \c0.n15_adj_4450\
        );

    \I__12603\ : LocalMux
    port map (
            O => \N__57788\,
            I => \c0.n15_adj_4450\
        );

    \I__12602\ : CascadeMux
    port map (
            O => \N__57783\,
            I => \N__57779\
        );

    \I__12601\ : InMux
    port map (
            O => \N__57782\,
            I => \N__57776\
        );

    \I__12600\ : InMux
    port map (
            O => \N__57779\,
            I => \N__57773\
        );

    \I__12599\ : LocalMux
    port map (
            O => \N__57776\,
            I => \N__57768\
        );

    \I__12598\ : LocalMux
    port map (
            O => \N__57773\,
            I => \N__57768\
        );

    \I__12597\ : Odrv12
    port map (
            O => \N__57768\,
            I => \c0.n87\
        );

    \I__12596\ : InMux
    port map (
            O => \N__57765\,
            I => \N__57762\
        );

    \I__12595\ : LocalMux
    port map (
            O => \N__57762\,
            I => \N__57759\
        );

    \I__12594\ : Span4Mux_v
    port map (
            O => \N__57759\,
            I => \N__57756\
        );

    \I__12593\ : Odrv4
    port map (
            O => \N__57756\,
            I => \c0.n85\
        );

    \I__12592\ : InMux
    port map (
            O => \N__57753\,
            I => \N__57750\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__57750\,
            I => \N__57747\
        );

    \I__12590\ : Span4Mux_h
    port map (
            O => \N__57747\,
            I => \N__57744\
        );

    \I__12589\ : Odrv4
    port map (
            O => \N__57744\,
            I => \c0.n88\
        );

    \I__12588\ : CascadeMux
    port map (
            O => \N__57741\,
            I => \c0.n87_cascade_\
        );

    \I__12587\ : InMux
    port map (
            O => \N__57738\,
            I => \N__57735\
        );

    \I__12586\ : LocalMux
    port map (
            O => \N__57735\,
            I => \c0.n106\
        );

    \I__12585\ : InMux
    port map (
            O => \N__57732\,
            I => \N__57725\
        );

    \I__12584\ : InMux
    port map (
            O => \N__57731\,
            I => \N__57722\
        );

    \I__12583\ : InMux
    port map (
            O => \N__57730\,
            I => \N__57714\
        );

    \I__12582\ : InMux
    port map (
            O => \N__57729\,
            I => \N__57714\
        );

    \I__12581\ : InMux
    port map (
            O => \N__57728\,
            I => \N__57714\
        );

    \I__12580\ : LocalMux
    port map (
            O => \N__57725\,
            I => \N__57711\
        );

    \I__12579\ : LocalMux
    port map (
            O => \N__57722\,
            I => \N__57708\
        );

    \I__12578\ : InMux
    port map (
            O => \N__57721\,
            I => \N__57705\
        );

    \I__12577\ : LocalMux
    port map (
            O => \N__57714\,
            I => \N__57702\
        );

    \I__12576\ : Span4Mux_v
    port map (
            O => \N__57711\,
            I => \N__57699\
        );

    \I__12575\ : Span4Mux_v
    port map (
            O => \N__57708\,
            I => \N__57694\
        );

    \I__12574\ : LocalMux
    port map (
            O => \N__57705\,
            I => \N__57694\
        );

    \I__12573\ : Span4Mux_h
    port map (
            O => \N__57702\,
            I => \N__57691\
        );

    \I__12572\ : Odrv4
    port map (
            O => \N__57699\,
            I => \c0.n22160\
        );

    \I__12571\ : Odrv4
    port map (
            O => \N__57694\,
            I => \c0.n22160\
        );

    \I__12570\ : Odrv4
    port map (
            O => \N__57691\,
            I => \c0.n22160\
        );

    \I__12569\ : InMux
    port map (
            O => \N__57684\,
            I => \N__57678\
        );

    \I__12568\ : InMux
    port map (
            O => \N__57683\,
            I => \N__57678\
        );

    \I__12567\ : LocalMux
    port map (
            O => \N__57678\,
            I => \c0.n7_adj_4304\
        );

    \I__12566\ : CascadeMux
    port map (
            O => \N__57675\,
            I => \c0.n7_adj_4304_cascade_\
        );

    \I__12565\ : CascadeMux
    port map (
            O => \N__57672\,
            I => \N__57668\
        );

    \I__12564\ : CascadeMux
    port map (
            O => \N__57671\,
            I => \N__57664\
        );

    \I__12563\ : InMux
    port map (
            O => \N__57668\,
            I => \N__57658\
        );

    \I__12562\ : InMux
    port map (
            O => \N__57667\,
            I => \N__57655\
        );

    \I__12561\ : InMux
    port map (
            O => \N__57664\,
            I => \N__57650\
        );

    \I__12560\ : InMux
    port map (
            O => \N__57663\,
            I => \N__57650\
        );

    \I__12559\ : InMux
    port map (
            O => \N__57662\,
            I => \N__57647\
        );

    \I__12558\ : InMux
    port map (
            O => \N__57661\,
            I => \N__57644\
        );

    \I__12557\ : LocalMux
    port map (
            O => \N__57658\,
            I => \N__57639\
        );

    \I__12556\ : LocalMux
    port map (
            O => \N__57655\,
            I => \N__57639\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__57650\,
            I => \N__57633\
        );

    \I__12554\ : LocalMux
    port map (
            O => \N__57647\,
            I => \N__57628\
        );

    \I__12553\ : LocalMux
    port map (
            O => \N__57644\,
            I => \N__57628\
        );

    \I__12552\ : Span4Mux_h
    port map (
            O => \N__57639\,
            I => \N__57625\
        );

    \I__12551\ : InMux
    port map (
            O => \N__57638\,
            I => \N__57620\
        );

    \I__12550\ : InMux
    port map (
            O => \N__57637\,
            I => \N__57620\
        );

    \I__12549\ : InMux
    port map (
            O => \N__57636\,
            I => \N__57617\
        );

    \I__12548\ : Odrv12
    port map (
            O => \N__57633\,
            I => data_in_frame_5_7
        );

    \I__12547\ : Odrv12
    port map (
            O => \N__57628\,
            I => data_in_frame_5_7
        );

    \I__12546\ : Odrv4
    port map (
            O => \N__57625\,
            I => data_in_frame_5_7
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__57620\,
            I => data_in_frame_5_7
        );

    \I__12544\ : LocalMux
    port map (
            O => \N__57617\,
            I => data_in_frame_5_7
        );

    \I__12543\ : InMux
    port map (
            O => \N__57606\,
            I => \N__57603\
        );

    \I__12542\ : LocalMux
    port map (
            O => \N__57603\,
            I => \N__57600\
        );

    \I__12541\ : Span4Mux_h
    port map (
            O => \N__57600\,
            I => \N__57597\
        );

    \I__12540\ : Sp12to4
    port map (
            O => \N__57597\,
            I => \N__57594\
        );

    \I__12539\ : Span12Mux_v
    port map (
            O => \N__57594\,
            I => \N__57589\
        );

    \I__12538\ : InMux
    port map (
            O => \N__57593\,
            I => \N__57584\
        );

    \I__12537\ : InMux
    port map (
            O => \N__57592\,
            I => \N__57584\
        );

    \I__12536\ : Odrv12
    port map (
            O => \N__57589\,
            I => data_in_frame_6_0
        );

    \I__12535\ : LocalMux
    port map (
            O => \N__57584\,
            I => data_in_frame_6_0
        );

    \I__12534\ : InMux
    port map (
            O => \N__57579\,
            I => \N__57576\
        );

    \I__12533\ : LocalMux
    port map (
            O => \N__57576\,
            I => \N__57573\
        );

    \I__12532\ : Span4Mux_v
    port map (
            O => \N__57573\,
            I => \N__57570\
        );

    \I__12531\ : Span4Mux_h
    port map (
            O => \N__57570\,
            I => \N__57567\
        );

    \I__12530\ : Odrv4
    port map (
            O => \N__57567\,
            I => \c0.n27_adj_4725\
        );

    \I__12529\ : InMux
    port map (
            O => \N__57564\,
            I => \N__57559\
        );

    \I__12528\ : InMux
    port map (
            O => \N__57563\,
            I => \N__57554\
        );

    \I__12527\ : InMux
    port map (
            O => \N__57562\,
            I => \N__57554\
        );

    \I__12526\ : LocalMux
    port map (
            O => \N__57559\,
            I => \N__57551\
        );

    \I__12525\ : LocalMux
    port map (
            O => \N__57554\,
            I => \N__57548\
        );

    \I__12524\ : Span4Mux_h
    port map (
            O => \N__57551\,
            I => \N__57545\
        );

    \I__12523\ : Span4Mux_v
    port map (
            O => \N__57548\,
            I => \N__57542\
        );

    \I__12522\ : Odrv4
    port map (
            O => \N__57545\,
            I => \c0.n13453\
        );

    \I__12521\ : Odrv4
    port map (
            O => \N__57542\,
            I => \c0.n13453\
        );

    \I__12520\ : InMux
    port map (
            O => \N__57537\,
            I => \N__57532\
        );

    \I__12519\ : InMux
    port map (
            O => \N__57536\,
            I => \N__57529\
        );

    \I__12518\ : CascadeMux
    port map (
            O => \N__57535\,
            I => \N__57526\
        );

    \I__12517\ : LocalMux
    port map (
            O => \N__57532\,
            I => \N__57523\
        );

    \I__12516\ : LocalMux
    port map (
            O => \N__57529\,
            I => \N__57520\
        );

    \I__12515\ : InMux
    port map (
            O => \N__57526\,
            I => \N__57517\
        );

    \I__12514\ : Odrv4
    port map (
            O => \N__57523\,
            I => \c0.n13_adj_4584\
        );

    \I__12513\ : Odrv12
    port map (
            O => \N__57520\,
            I => \c0.n13_adj_4584\
        );

    \I__12512\ : LocalMux
    port map (
            O => \N__57517\,
            I => \c0.n13_adj_4584\
        );

    \I__12511\ : CascadeMux
    port map (
            O => \N__57510\,
            I => \c0.n15_adj_4444_cascade_\
        );

    \I__12510\ : InMux
    port map (
            O => \N__57507\,
            I => \N__57504\
        );

    \I__12509\ : LocalMux
    port map (
            O => \N__57504\,
            I => \N__57501\
        );

    \I__12508\ : Span4Mux_h
    port map (
            O => \N__57501\,
            I => \N__57498\
        );

    \I__12507\ : Odrv4
    port map (
            O => \N__57498\,
            I => \c0.n11_adj_4656\
        );

    \I__12506\ : InMux
    port map (
            O => \N__57495\,
            I => \N__57489\
        );

    \I__12505\ : InMux
    port map (
            O => \N__57494\,
            I => \N__57489\
        );

    \I__12504\ : LocalMux
    port map (
            O => \N__57489\,
            I => \N__57485\
        );

    \I__12503\ : CascadeMux
    port map (
            O => \N__57488\,
            I => \N__57480\
        );

    \I__12502\ : Span4Mux_h
    port map (
            O => \N__57485\,
            I => \N__57477\
        );

    \I__12501\ : InMux
    port map (
            O => \N__57484\,
            I => \N__57474\
        );

    \I__12500\ : InMux
    port map (
            O => \N__57483\,
            I => \N__57469\
        );

    \I__12499\ : InMux
    port map (
            O => \N__57480\,
            I => \N__57469\
        );

    \I__12498\ : Odrv4
    port map (
            O => \N__57477\,
            I => \c0.data_in_frame_3_2\
        );

    \I__12497\ : LocalMux
    port map (
            O => \N__57474\,
            I => \c0.data_in_frame_3_2\
        );

    \I__12496\ : LocalMux
    port map (
            O => \N__57469\,
            I => \c0.data_in_frame_3_2\
        );

    \I__12495\ : CascadeMux
    port map (
            O => \N__57462\,
            I => \N__57457\
        );

    \I__12494\ : InMux
    port map (
            O => \N__57461\,
            I => \N__57450\
        );

    \I__12493\ : InMux
    port map (
            O => \N__57460\,
            I => \N__57450\
        );

    \I__12492\ : InMux
    port map (
            O => \N__57457\,
            I => \N__57450\
        );

    \I__12491\ : LocalMux
    port map (
            O => \N__57450\,
            I => data_in_frame_5_4
        );

    \I__12490\ : CascadeMux
    port map (
            O => \N__57447\,
            I => \N__57444\
        );

    \I__12489\ : InMux
    port map (
            O => \N__57444\,
            I => \N__57441\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__57441\,
            I => \c0.n6_adj_4611\
        );

    \I__12487\ : CascadeMux
    port map (
            O => \N__57438\,
            I => \c0.n6_adj_4611_cascade_\
        );

    \I__12486\ : InMux
    port map (
            O => \N__57435\,
            I => \N__57432\
        );

    \I__12485\ : LocalMux
    port map (
            O => \N__57432\,
            I => \N__57429\
        );

    \I__12484\ : Span4Mux_v
    port map (
            O => \N__57429\,
            I => \N__57425\
        );

    \I__12483\ : InMux
    port map (
            O => \N__57428\,
            I => \N__57422\
        );

    \I__12482\ : Odrv4
    port map (
            O => \N__57425\,
            I => \c0.n91\
        );

    \I__12481\ : LocalMux
    port map (
            O => \N__57422\,
            I => \c0.n91\
        );

    \I__12480\ : CascadeMux
    port map (
            O => \N__57417\,
            I => \N__57413\
        );

    \I__12479\ : InMux
    port map (
            O => \N__57416\,
            I => \N__57410\
        );

    \I__12478\ : InMux
    port map (
            O => \N__57413\,
            I => \N__57406\
        );

    \I__12477\ : LocalMux
    port map (
            O => \N__57410\,
            I => \N__57403\
        );

    \I__12476\ : CascadeMux
    port map (
            O => \N__57409\,
            I => \N__57400\
        );

    \I__12475\ : LocalMux
    port map (
            O => \N__57406\,
            I => \N__57396\
        );

    \I__12474\ : Span4Mux_v
    port map (
            O => \N__57403\,
            I => \N__57393\
        );

    \I__12473\ : InMux
    port map (
            O => \N__57400\,
            I => \N__57388\
        );

    \I__12472\ : InMux
    port map (
            O => \N__57399\,
            I => \N__57388\
        );

    \I__12471\ : Odrv4
    port map (
            O => \N__57396\,
            I => \c0.data_in_frame_9_6\
        );

    \I__12470\ : Odrv4
    port map (
            O => \N__57393\,
            I => \c0.data_in_frame_9_6\
        );

    \I__12469\ : LocalMux
    port map (
            O => \N__57388\,
            I => \c0.data_in_frame_9_6\
        );

    \I__12468\ : InMux
    port map (
            O => \N__57381\,
            I => \N__57378\
        );

    \I__12467\ : LocalMux
    port map (
            O => \N__57378\,
            I => \N__57373\
        );

    \I__12466\ : InMux
    port map (
            O => \N__57377\,
            I => \N__57370\
        );

    \I__12465\ : CascadeMux
    port map (
            O => \N__57376\,
            I => \N__57367\
        );

    \I__12464\ : Span4Mux_h
    port map (
            O => \N__57373\,
            I => \N__57362\
        );

    \I__12463\ : LocalMux
    port map (
            O => \N__57370\,
            I => \N__57359\
        );

    \I__12462\ : InMux
    port map (
            O => \N__57367\,
            I => \N__57356\
        );

    \I__12461\ : InMux
    port map (
            O => \N__57366\,
            I => \N__57352\
        );

    \I__12460\ : InMux
    port map (
            O => \N__57365\,
            I => \N__57349\
        );

    \I__12459\ : Span4Mux_v
    port map (
            O => \N__57362\,
            I => \N__57346\
        );

    \I__12458\ : Span4Mux_v
    port map (
            O => \N__57359\,
            I => \N__57343\
        );

    \I__12457\ : LocalMux
    port map (
            O => \N__57356\,
            I => \N__57340\
        );

    \I__12456\ : InMux
    port map (
            O => \N__57355\,
            I => \N__57337\
        );

    \I__12455\ : LocalMux
    port map (
            O => \N__57352\,
            I => data_in_frame_5_3
        );

    \I__12454\ : LocalMux
    port map (
            O => \N__57349\,
            I => data_in_frame_5_3
        );

    \I__12453\ : Odrv4
    port map (
            O => \N__57346\,
            I => data_in_frame_5_3
        );

    \I__12452\ : Odrv4
    port map (
            O => \N__57343\,
            I => data_in_frame_5_3
        );

    \I__12451\ : Odrv12
    port map (
            O => \N__57340\,
            I => data_in_frame_5_3
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__57337\,
            I => data_in_frame_5_3
        );

    \I__12449\ : InMux
    port map (
            O => \N__57324\,
            I => \N__57319\
        );

    \I__12448\ : InMux
    port map (
            O => \N__57323\,
            I => \N__57314\
        );

    \I__12447\ : InMux
    port map (
            O => \N__57322\,
            I => \N__57314\
        );

    \I__12446\ : LocalMux
    port map (
            O => \N__57319\,
            I => data_in_frame_5_2
        );

    \I__12445\ : LocalMux
    port map (
            O => \N__57314\,
            I => data_in_frame_5_2
        );

    \I__12444\ : CascadeMux
    port map (
            O => \N__57309\,
            I => \N__57305\
        );

    \I__12443\ : CascadeMux
    port map (
            O => \N__57308\,
            I => \N__57302\
        );

    \I__12442\ : InMux
    port map (
            O => \N__57305\,
            I => \N__57299\
        );

    \I__12441\ : InMux
    port map (
            O => \N__57302\,
            I => \N__57294\
        );

    \I__12440\ : LocalMux
    port map (
            O => \N__57299\,
            I => \N__57291\
        );

    \I__12439\ : InMux
    port map (
            O => \N__57298\,
            I => \N__57286\
        );

    \I__12438\ : InMux
    port map (
            O => \N__57297\,
            I => \N__57286\
        );

    \I__12437\ : LocalMux
    port map (
            O => \N__57294\,
            I => \N__57283\
        );

    \I__12436\ : Span4Mux_h
    port map (
            O => \N__57291\,
            I => \N__57280\
        );

    \I__12435\ : LocalMux
    port map (
            O => \N__57286\,
            I => \N__57277\
        );

    \I__12434\ : Odrv4
    port map (
            O => \N__57283\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12433\ : Odrv4
    port map (
            O => \N__57280\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12432\ : Odrv12
    port map (
            O => \N__57277\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12431\ : InMux
    port map (
            O => \N__57270\,
            I => \N__57267\
        );

    \I__12430\ : LocalMux
    port map (
            O => \N__57267\,
            I => \N__57264\
        );

    \I__12429\ : Span4Mux_v
    port map (
            O => \N__57264\,
            I => \N__57260\
        );

    \I__12428\ : CascadeMux
    port map (
            O => \N__57263\,
            I => \N__57257\
        );

    \I__12427\ : Span4Mux_h
    port map (
            O => \N__57260\,
            I => \N__57254\
        );

    \I__12426\ : InMux
    port map (
            O => \N__57257\,
            I => \N__57251\
        );

    \I__12425\ : Span4Mux_v
    port map (
            O => \N__57254\,
            I => \N__57246\
        );

    \I__12424\ : LocalMux
    port map (
            O => \N__57251\,
            I => \N__57246\
        );

    \I__12423\ : Span4Mux_v
    port map (
            O => \N__57246\,
            I => \N__57240\
        );

    \I__12422\ : InMux
    port map (
            O => \N__57245\,
            I => \N__57237\
        );

    \I__12421\ : CascadeMux
    port map (
            O => \N__57244\,
            I => \N__57229\
        );

    \I__12420\ : InMux
    port map (
            O => \N__57243\,
            I => \N__57225\
        );

    \I__12419\ : Sp12to4
    port map (
            O => \N__57240\,
            I => \N__57220\
        );

    \I__12418\ : LocalMux
    port map (
            O => \N__57237\,
            I => \N__57220\
        );

    \I__12417\ : InMux
    port map (
            O => \N__57236\,
            I => \N__57213\
        );

    \I__12416\ : InMux
    port map (
            O => \N__57235\,
            I => \N__57213\
        );

    \I__12415\ : InMux
    port map (
            O => \N__57234\,
            I => \N__57213\
        );

    \I__12414\ : InMux
    port map (
            O => \N__57233\,
            I => \N__57208\
        );

    \I__12413\ : InMux
    port map (
            O => \N__57232\,
            I => \N__57208\
        );

    \I__12412\ : InMux
    port map (
            O => \N__57229\,
            I => \N__57203\
        );

    \I__12411\ : InMux
    port map (
            O => \N__57228\,
            I => \N__57203\
        );

    \I__12410\ : LocalMux
    port map (
            O => \N__57225\,
            I => data_in_frame_1_2
        );

    \I__12409\ : Odrv12
    port map (
            O => \N__57220\,
            I => data_in_frame_1_2
        );

    \I__12408\ : LocalMux
    port map (
            O => \N__57213\,
            I => data_in_frame_1_2
        );

    \I__12407\ : LocalMux
    port map (
            O => \N__57208\,
            I => data_in_frame_1_2
        );

    \I__12406\ : LocalMux
    port map (
            O => \N__57203\,
            I => data_in_frame_1_2
        );

    \I__12405\ : InMux
    port map (
            O => \N__57192\,
            I => \N__57189\
        );

    \I__12404\ : LocalMux
    port map (
            O => \N__57189\,
            I => \c0.n12_adj_4612\
        );

    \I__12403\ : InMux
    port map (
            O => \N__57186\,
            I => \N__57183\
        );

    \I__12402\ : LocalMux
    port map (
            O => \N__57183\,
            I => \N__57180\
        );

    \I__12401\ : Span4Mux_h
    port map (
            O => \N__57180\,
            I => \N__57177\
        );

    \I__12400\ : Odrv4
    port map (
            O => \N__57177\,
            I => \c0.n15_adj_4444\
        );

    \I__12399\ : InMux
    port map (
            O => \N__57174\,
            I => \N__57171\
        );

    \I__12398\ : LocalMux
    port map (
            O => \N__57171\,
            I => \N__57168\
        );

    \I__12397\ : Span4Mux_h
    port map (
            O => \N__57168\,
            I => \N__57165\
        );

    \I__12396\ : Odrv4
    port map (
            O => \N__57165\,
            I => \c0.n70_adj_4514\
        );

    \I__12395\ : CascadeMux
    port map (
            O => \N__57162\,
            I => \c0.n71_cascade_\
        );

    \I__12394\ : CascadeMux
    port map (
            O => \N__57159\,
            I => \N__57156\
        );

    \I__12393\ : InMux
    port map (
            O => \N__57156\,
            I => \N__57152\
        );

    \I__12392\ : InMux
    port map (
            O => \N__57155\,
            I => \N__57149\
        );

    \I__12391\ : LocalMux
    port map (
            O => \N__57152\,
            I => \N__57146\
        );

    \I__12390\ : LocalMux
    port map (
            O => \N__57149\,
            I => \N__57143\
        );

    \I__12389\ : Span4Mux_h
    port map (
            O => \N__57146\,
            I => \N__57140\
        );

    \I__12388\ : Span12Mux_v
    port map (
            O => \N__57143\,
            I => \N__57137\
        );

    \I__12387\ : Span4Mux_h
    port map (
            O => \N__57140\,
            I => \N__57134\
        );

    \I__12386\ : Odrv12
    port map (
            O => \N__57137\,
            I => \c0.n17537\
        );

    \I__12385\ : Odrv4
    port map (
            O => \N__57134\,
            I => \c0.n17537\
        );

    \I__12384\ : CascadeMux
    port map (
            O => \N__57129\,
            I => \c0.n81_cascade_\
        );

    \I__12383\ : InMux
    port map (
            O => \N__57126\,
            I => \N__57123\
        );

    \I__12382\ : LocalMux
    port map (
            O => \N__57123\,
            I => \c0.n82_adj_4517\
        );

    \I__12381\ : InMux
    port map (
            O => \N__57120\,
            I => \N__57117\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__57117\,
            I => \c0.n28_adj_4523\
        );

    \I__12379\ : InMux
    port map (
            O => \N__57114\,
            I => \N__57109\
        );

    \I__12378\ : InMux
    port map (
            O => \N__57113\,
            I => \N__57106\
        );

    \I__12377\ : CascadeMux
    port map (
            O => \N__57112\,
            I => \N__57103\
        );

    \I__12376\ : LocalMux
    port map (
            O => \N__57109\,
            I => \N__57099\
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__57106\,
            I => \N__57096\
        );

    \I__12374\ : InMux
    port map (
            O => \N__57103\,
            I => \N__57091\
        );

    \I__12373\ : InMux
    port map (
            O => \N__57102\,
            I => \N__57091\
        );

    \I__12372\ : Span4Mux_h
    port map (
            O => \N__57099\,
            I => \N__57088\
        );

    \I__12371\ : Odrv12
    port map (
            O => \N__57096\,
            I => \c0.data_in_frame_27_3\
        );

    \I__12370\ : LocalMux
    port map (
            O => \N__57091\,
            I => \c0.data_in_frame_27_3\
        );

    \I__12369\ : Odrv4
    port map (
            O => \N__57088\,
            I => \c0.data_in_frame_27_3\
        );

    \I__12368\ : CascadeMux
    port map (
            O => \N__57081\,
            I => \N__57077\
        );

    \I__12367\ : InMux
    port map (
            O => \N__57080\,
            I => \N__57073\
        );

    \I__12366\ : InMux
    port map (
            O => \N__57077\,
            I => \N__57069\
        );

    \I__12365\ : InMux
    port map (
            O => \N__57076\,
            I => \N__57066\
        );

    \I__12364\ : LocalMux
    port map (
            O => \N__57073\,
            I => \N__57063\
        );

    \I__12363\ : InMux
    port map (
            O => \N__57072\,
            I => \N__57060\
        );

    \I__12362\ : LocalMux
    port map (
            O => \N__57069\,
            I => \N__57053\
        );

    \I__12361\ : LocalMux
    port map (
            O => \N__57066\,
            I => \N__57053\
        );

    \I__12360\ : Span4Mux_v
    port map (
            O => \N__57063\,
            I => \N__57053\
        );

    \I__12359\ : LocalMux
    port map (
            O => \N__57060\,
            I => \c0.data_in_frame_27_4\
        );

    \I__12358\ : Odrv4
    port map (
            O => \N__57053\,
            I => \c0.data_in_frame_27_4\
        );

    \I__12357\ : CascadeMux
    port map (
            O => \N__57048\,
            I => \c0.n23_adj_4532_cascade_\
        );

    \I__12356\ : InMux
    port map (
            O => \N__57045\,
            I => \N__57042\
        );

    \I__12355\ : LocalMux
    port map (
            O => \N__57042\,
            I => \c0.n31_adj_4542\
        );

    \I__12354\ : CascadeMux
    port map (
            O => \N__57039\,
            I => \c0.n38_adj_4535_cascade_\
        );

    \I__12353\ : InMux
    port map (
            O => \N__57036\,
            I => \N__57033\
        );

    \I__12352\ : LocalMux
    port map (
            O => \N__57033\,
            I => \c0.n32_adj_4534\
        );

    \I__12351\ : InMux
    port map (
            O => \N__57030\,
            I => \N__57027\
        );

    \I__12350\ : LocalMux
    port map (
            O => \N__57027\,
            I => \N__57024\
        );

    \I__12349\ : Odrv4
    port map (
            O => \N__57024\,
            I => \c0.n8_adj_4677\
        );

    \I__12348\ : CascadeMux
    port map (
            O => \N__57021\,
            I => \N__57018\
        );

    \I__12347\ : InMux
    port map (
            O => \N__57018\,
            I => \N__57011\
        );

    \I__12346\ : InMux
    port map (
            O => \N__57017\,
            I => \N__57002\
        );

    \I__12345\ : InMux
    port map (
            O => \N__57016\,
            I => \N__57002\
        );

    \I__12344\ : InMux
    port map (
            O => \N__57015\,
            I => \N__57002\
        );

    \I__12343\ : InMux
    port map (
            O => \N__57014\,
            I => \N__57002\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__57011\,
            I => \N__56998\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__57002\,
            I => \N__56995\
        );

    \I__12340\ : CascadeMux
    port map (
            O => \N__57001\,
            I => \N__56991\
        );

    \I__12339\ : Span4Mux_v
    port map (
            O => \N__56998\,
            I => \N__56988\
        );

    \I__12338\ : Span4Mux_v
    port map (
            O => \N__56995\,
            I => \N__56985\
        );

    \I__12337\ : InMux
    port map (
            O => \N__56994\,
            I => \N__56980\
        );

    \I__12336\ : InMux
    port map (
            O => \N__56991\,
            I => \N__56980\
        );

    \I__12335\ : Odrv4
    port map (
            O => \N__56988\,
            I => \c0.data_in_frame_25_0\
        );

    \I__12334\ : Odrv4
    port map (
            O => \N__56985\,
            I => \c0.data_in_frame_25_0\
        );

    \I__12333\ : LocalMux
    port map (
            O => \N__56980\,
            I => \c0.data_in_frame_25_0\
        );

    \I__12332\ : InMux
    port map (
            O => \N__56973\,
            I => \N__56970\
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__56970\,
            I => \N__56967\
        );

    \I__12330\ : Odrv4
    port map (
            O => \N__56967\,
            I => \c0.n64_adj_4539\
        );

    \I__12329\ : InMux
    port map (
            O => \N__56964\,
            I => \N__56961\
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__56961\,
            I => \N__56958\
        );

    \I__12327\ : Odrv4
    port map (
            O => \N__56958\,
            I => \c0.n10_adj_4544\
        );

    \I__12326\ : InMux
    port map (
            O => \N__56955\,
            I => \N__56952\
        );

    \I__12325\ : LocalMux
    port map (
            O => \N__56952\,
            I => \c0.n13911\
        );

    \I__12324\ : CascadeMux
    port map (
            O => \N__56949\,
            I => \c0.n23921_cascade_\
        );

    \I__12323\ : InMux
    port map (
            O => \N__56946\,
            I => \N__56943\
        );

    \I__12322\ : LocalMux
    port map (
            O => \N__56943\,
            I => \N__56940\
        );

    \I__12321\ : Span4Mux_h
    port map (
            O => \N__56940\,
            I => \N__56937\
        );

    \I__12320\ : Odrv4
    port map (
            O => \N__56937\,
            I => \c0.n21_adj_4547\
        );

    \I__12319\ : InMux
    port map (
            O => \N__56934\,
            I => \N__56931\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__56931\,
            I => \N__56928\
        );

    \I__12317\ : Odrv12
    port map (
            O => \N__56928\,
            I => \c0.n23975\
        );

    \I__12316\ : CascadeMux
    port map (
            O => \N__56925\,
            I => \N__56922\
        );

    \I__12315\ : InMux
    port map (
            O => \N__56922\,
            I => \N__56919\
        );

    \I__12314\ : LocalMux
    port map (
            O => \N__56919\,
            I => \N__56916\
        );

    \I__12313\ : Span4Mux_h
    port map (
            O => \N__56916\,
            I => \N__56913\
        );

    \I__12312\ : Odrv4
    port map (
            O => \N__56913\,
            I => \c0.n32_adj_4533\
        );

    \I__12311\ : InMux
    port map (
            O => \N__56910\,
            I => \N__56907\
        );

    \I__12310\ : LocalMux
    port map (
            O => \N__56907\,
            I => \c0.n74\
        );

    \I__12309\ : InMux
    port map (
            O => \N__56904\,
            I => \N__56898\
        );

    \I__12308\ : InMux
    port map (
            O => \N__56903\,
            I => \N__56898\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__56898\,
            I => \c0.data_in_frame_29_7\
        );

    \I__12306\ : InMux
    port map (
            O => \N__56895\,
            I => \N__56890\
        );

    \I__12305\ : InMux
    port map (
            O => \N__56894\,
            I => \N__56887\
        );

    \I__12304\ : InMux
    port map (
            O => \N__56893\,
            I => \N__56883\
        );

    \I__12303\ : LocalMux
    port map (
            O => \N__56890\,
            I => \N__56878\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__56887\,
            I => \N__56878\
        );

    \I__12301\ : InMux
    port map (
            O => \N__56886\,
            I => \N__56875\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__56883\,
            I => \N__56872\
        );

    \I__12299\ : Span4Mux_v
    port map (
            O => \N__56878\,
            I => \N__56869\
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__56875\,
            I => \c0.data_in_frame_27_5\
        );

    \I__12297\ : Odrv4
    port map (
            O => \N__56872\,
            I => \c0.data_in_frame_27_5\
        );

    \I__12296\ : Odrv4
    port map (
            O => \N__56869\,
            I => \c0.data_in_frame_27_5\
        );

    \I__12295\ : InMux
    port map (
            O => \N__56862\,
            I => \N__56859\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__56859\,
            I => \N__56855\
        );

    \I__12293\ : InMux
    port map (
            O => \N__56858\,
            I => \N__56850\
        );

    \I__12292\ : Span4Mux_v
    port map (
            O => \N__56855\,
            I => \N__56847\
        );

    \I__12291\ : InMux
    port map (
            O => \N__56854\,
            I => \N__56844\
        );

    \I__12290\ : CascadeMux
    port map (
            O => \N__56853\,
            I => \N__56841\
        );

    \I__12289\ : LocalMux
    port map (
            O => \N__56850\,
            I => \N__56836\
        );

    \I__12288\ : Span4Mux_h
    port map (
            O => \N__56847\,
            I => \N__56836\
        );

    \I__12287\ : LocalMux
    port map (
            O => \N__56844\,
            I => \N__56833\
        );

    \I__12286\ : InMux
    port map (
            O => \N__56841\,
            I => \N__56830\
        );

    \I__12285\ : Span4Mux_h
    port map (
            O => \N__56836\,
            I => \N__56827\
        );

    \I__12284\ : Span4Mux_v
    port map (
            O => \N__56833\,
            I => \N__56824\
        );

    \I__12283\ : LocalMux
    port map (
            O => \N__56830\,
            I => \c0.data_in_frame_27_6\
        );

    \I__12282\ : Odrv4
    port map (
            O => \N__56827\,
            I => \c0.data_in_frame_27_6\
        );

    \I__12281\ : Odrv4
    port map (
            O => \N__56824\,
            I => \c0.data_in_frame_27_6\
        );

    \I__12280\ : InMux
    port map (
            O => \N__56817\,
            I => \N__56811\
        );

    \I__12279\ : CascadeMux
    port map (
            O => \N__56816\,
            I => \N__56808\
        );

    \I__12278\ : InMux
    port map (
            O => \N__56815\,
            I => \N__56805\
        );

    \I__12277\ : InMux
    port map (
            O => \N__56814\,
            I => \N__56802\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__56811\,
            I => \N__56799\
        );

    \I__12275\ : InMux
    port map (
            O => \N__56808\,
            I => \N__56794\
        );

    \I__12274\ : LocalMux
    port map (
            O => \N__56805\,
            I => \N__56791\
        );

    \I__12273\ : LocalMux
    port map (
            O => \N__56802\,
            I => \N__56788\
        );

    \I__12272\ : Span4Mux_v
    port map (
            O => \N__56799\,
            I => \N__56785\
        );

    \I__12271\ : InMux
    port map (
            O => \N__56798\,
            I => \N__56780\
        );

    \I__12270\ : InMux
    port map (
            O => \N__56797\,
            I => \N__56780\
        );

    \I__12269\ : LocalMux
    port map (
            O => \N__56794\,
            I => \N__56773\
        );

    \I__12268\ : Span4Mux_v
    port map (
            O => \N__56791\,
            I => \N__56773\
        );

    \I__12267\ : Span4Mux_h
    port map (
            O => \N__56788\,
            I => \N__56773\
        );

    \I__12266\ : Odrv4
    port map (
            O => \N__56785\,
            I => \c0.data_in_frame_25_5\
        );

    \I__12265\ : LocalMux
    port map (
            O => \N__56780\,
            I => \c0.data_in_frame_25_5\
        );

    \I__12264\ : Odrv4
    port map (
            O => \N__56773\,
            I => \c0.data_in_frame_25_5\
        );

    \I__12263\ : InMux
    port map (
            O => \N__56766\,
            I => \N__56763\
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__56763\,
            I => \c0.n12_adj_4466\
        );

    \I__12261\ : CascadeMux
    port map (
            O => \N__56760\,
            I => \c0.n11_adj_4474_cascade_\
        );

    \I__12260\ : InMux
    port map (
            O => \N__56757\,
            I => \N__56754\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__56754\,
            I => \N__56748\
        );

    \I__12258\ : InMux
    port map (
            O => \N__56753\,
            I => \N__56745\
        );

    \I__12257\ : InMux
    port map (
            O => \N__56752\,
            I => \N__56742\
        );

    \I__12256\ : InMux
    port map (
            O => \N__56751\,
            I => \N__56739\
        );

    \I__12255\ : Span4Mux_h
    port map (
            O => \N__56748\,
            I => \N__56733\
        );

    \I__12254\ : LocalMux
    port map (
            O => \N__56745\,
            I => \N__56726\
        );

    \I__12253\ : LocalMux
    port map (
            O => \N__56742\,
            I => \N__56726\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__56739\,
            I => \N__56726\
        );

    \I__12251\ : InMux
    port map (
            O => \N__56738\,
            I => \N__56719\
        );

    \I__12250\ : InMux
    port map (
            O => \N__56737\,
            I => \N__56719\
        );

    \I__12249\ : InMux
    port map (
            O => \N__56736\,
            I => \N__56719\
        );

    \I__12248\ : Odrv4
    port map (
            O => \N__56733\,
            I => \c0.n21280\
        );

    \I__12247\ : Odrv4
    port map (
            O => \N__56726\,
            I => \c0.n21280\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__56719\,
            I => \c0.n21280\
        );

    \I__12245\ : CascadeMux
    port map (
            O => \N__56712\,
            I => \N__56709\
        );

    \I__12244\ : InMux
    port map (
            O => \N__56709\,
            I => \N__56706\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__56706\,
            I => \N__56702\
        );

    \I__12242\ : InMux
    port map (
            O => \N__56705\,
            I => \N__56699\
        );

    \I__12241\ : Span4Mux_v
    port map (
            O => \N__56702\,
            I => \N__56696\
        );

    \I__12240\ : LocalMux
    port map (
            O => \N__56699\,
            I => \c0.data_in_frame_29_2\
        );

    \I__12239\ : Odrv4
    port map (
            O => \N__56696\,
            I => \c0.data_in_frame_29_2\
        );

    \I__12238\ : InMux
    port map (
            O => \N__56691\,
            I => \N__56688\
        );

    \I__12237\ : LocalMux
    port map (
            O => \N__56688\,
            I => \c0.n25446\
        );

    \I__12236\ : CascadeMux
    port map (
            O => \N__56685\,
            I => \N__56681\
        );

    \I__12235\ : InMux
    port map (
            O => \N__56684\,
            I => \N__56678\
        );

    \I__12234\ : InMux
    port map (
            O => \N__56681\,
            I => \N__56675\
        );

    \I__12233\ : LocalMux
    port map (
            O => \N__56678\,
            I => \c0.data_in_frame_29_0\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__56675\,
            I => \c0.data_in_frame_29_0\
        );

    \I__12231\ : InMux
    port map (
            O => \N__56670\,
            I => \N__56666\
        );

    \I__12230\ : InMux
    port map (
            O => \N__56669\,
            I => \N__56663\
        );

    \I__12229\ : LocalMux
    port map (
            O => \N__56666\,
            I => \N__56658\
        );

    \I__12228\ : LocalMux
    port map (
            O => \N__56663\,
            I => \N__56658\
        );

    \I__12227\ : Odrv4
    port map (
            O => \N__56658\,
            I => \c0.n10874\
        );

    \I__12226\ : CascadeMux
    port map (
            O => \N__56655\,
            I => \c0.n43_adj_4463_cascade_\
        );

    \I__12225\ : InMux
    port map (
            O => \N__56652\,
            I => \N__56642\
        );

    \I__12224\ : InMux
    port map (
            O => \N__56651\,
            I => \N__56642\
        );

    \I__12223\ : InMux
    port map (
            O => \N__56650\,
            I => \N__56642\
        );

    \I__12222\ : CascadeMux
    port map (
            O => \N__56649\,
            I => \N__56639\
        );

    \I__12221\ : LocalMux
    port map (
            O => \N__56642\,
            I => \N__56636\
        );

    \I__12220\ : InMux
    port map (
            O => \N__56639\,
            I => \N__56633\
        );

    \I__12219\ : Span4Mux_v
    port map (
            O => \N__56636\,
            I => \N__56629\
        );

    \I__12218\ : LocalMux
    port map (
            O => \N__56633\,
            I => \N__56626\
        );

    \I__12217\ : InMux
    port map (
            O => \N__56632\,
            I => \N__56623\
        );

    \I__12216\ : Span4Mux_h
    port map (
            O => \N__56629\,
            I => \N__56620\
        );

    \I__12215\ : Span4Mux_v
    port map (
            O => \N__56626\,
            I => \N__56617\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__56623\,
            I => \c0.n21389\
        );

    \I__12213\ : Odrv4
    port map (
            O => \N__56620\,
            I => \c0.n21389\
        );

    \I__12212\ : Odrv4
    port map (
            O => \N__56617\,
            I => \c0.n21389\
        );

    \I__12211\ : InMux
    port map (
            O => \N__56610\,
            I => \N__56607\
        );

    \I__12210\ : LocalMux
    port map (
            O => \N__56607\,
            I => \c0.n9_adj_4521\
        );

    \I__12209\ : InMux
    port map (
            O => \N__56604\,
            I => \N__56601\
        );

    \I__12208\ : LocalMux
    port map (
            O => \N__56601\,
            I => \c0.n20_adj_4596\
        );

    \I__12207\ : CascadeMux
    port map (
            O => \N__56598\,
            I => \c0.n23733_cascade_\
        );

    \I__12206\ : InMux
    port map (
            O => \N__56595\,
            I => \N__56589\
        );

    \I__12205\ : InMux
    port map (
            O => \N__56594\,
            I => \N__56589\
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__56589\,
            I => \N__56585\
        );

    \I__12203\ : InMux
    port map (
            O => \N__56588\,
            I => \N__56582\
        );

    \I__12202\ : Span4Mux_v
    port map (
            O => \N__56585\,
            I => \N__56579\
        );

    \I__12201\ : LocalMux
    port map (
            O => \N__56582\,
            I => \c0.data_in_frame_26_0\
        );

    \I__12200\ : Odrv4
    port map (
            O => \N__56579\,
            I => \c0.data_in_frame_26_0\
        );

    \I__12199\ : CascadeMux
    port map (
            O => \N__56574\,
            I => \N__56569\
        );

    \I__12198\ : InMux
    port map (
            O => \N__56573\,
            I => \N__56564\
        );

    \I__12197\ : InMux
    port map (
            O => \N__56572\,
            I => \N__56564\
        );

    \I__12196\ : InMux
    port map (
            O => \N__56569\,
            I => \N__56561\
        );

    \I__12195\ : LocalMux
    port map (
            O => \N__56564\,
            I => \N__56557\
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__56561\,
            I => \N__56554\
        );

    \I__12193\ : CascadeMux
    port map (
            O => \N__56560\,
            I => \N__56551\
        );

    \I__12192\ : Span4Mux_v
    port map (
            O => \N__56557\,
            I => \N__56548\
        );

    \I__12191\ : Span4Mux_h
    port map (
            O => \N__56554\,
            I => \N__56545\
        );

    \I__12190\ : InMux
    port map (
            O => \N__56551\,
            I => \N__56542\
        );

    \I__12189\ : Span4Mux_h
    port map (
            O => \N__56548\,
            I => \N__56539\
        );

    \I__12188\ : Span4Mux_v
    port map (
            O => \N__56545\,
            I => \N__56536\
        );

    \I__12187\ : LocalMux
    port map (
            O => \N__56542\,
            I => \c0.data_in_frame_27_7\
        );

    \I__12186\ : Odrv4
    port map (
            O => \N__56539\,
            I => \c0.data_in_frame_27_7\
        );

    \I__12185\ : Odrv4
    port map (
            O => \N__56536\,
            I => \c0.data_in_frame_27_7\
        );

    \I__12184\ : CascadeMux
    port map (
            O => \N__56529\,
            I => \c0.n20314_cascade_\
        );

    \I__12183\ : InMux
    port map (
            O => \N__56526\,
            I => \N__56523\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__56523\,
            I => \N__56519\
        );

    \I__12181\ : InMux
    port map (
            O => \N__56522\,
            I => \N__56516\
        );

    \I__12180\ : Span4Mux_v
    port map (
            O => \N__56519\,
            I => \N__56512\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__56516\,
            I => \N__56509\
        );

    \I__12178\ : InMux
    port map (
            O => \N__56515\,
            I => \N__56506\
        );

    \I__12177\ : Odrv4
    port map (
            O => \N__56512\,
            I => \c0.n21325\
        );

    \I__12176\ : Odrv12
    port map (
            O => \N__56509\,
            I => \c0.n21325\
        );

    \I__12175\ : LocalMux
    port map (
            O => \N__56506\,
            I => \c0.n21325\
        );

    \I__12174\ : InMux
    port map (
            O => \N__56499\,
            I => \N__56496\
        );

    \I__12173\ : LocalMux
    port map (
            O => \N__56496\,
            I => \c0.n20314\
        );

    \I__12172\ : InMux
    port map (
            O => \N__56493\,
            I => \N__56490\
        );

    \I__12171\ : LocalMux
    port map (
            O => \N__56490\,
            I => \c0.n22_adj_4597\
        );

    \I__12170\ : InMux
    port map (
            O => \N__56487\,
            I => \N__56484\
        );

    \I__12169\ : LocalMux
    port map (
            O => \N__56484\,
            I => \N__56476\
        );

    \I__12168\ : InMux
    port map (
            O => \N__56483\,
            I => \N__56471\
        );

    \I__12167\ : InMux
    port map (
            O => \N__56482\,
            I => \N__56471\
        );

    \I__12166\ : InMux
    port map (
            O => \N__56481\,
            I => \N__56468\
        );

    \I__12165\ : InMux
    port map (
            O => \N__56480\,
            I => \N__56465\
        );

    \I__12164\ : CascadeMux
    port map (
            O => \N__56479\,
            I => \N__56462\
        );

    \I__12163\ : Span4Mux_h
    port map (
            O => \N__56476\,
            I => \N__56456\
        );

    \I__12162\ : LocalMux
    port map (
            O => \N__56471\,
            I => \N__56456\
        );

    \I__12161\ : LocalMux
    port map (
            O => \N__56468\,
            I => \N__56453\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__56465\,
            I => \N__56450\
        );

    \I__12159\ : InMux
    port map (
            O => \N__56462\,
            I => \N__56445\
        );

    \I__12158\ : InMux
    port map (
            O => \N__56461\,
            I => \N__56445\
        );

    \I__12157\ : Span4Mux_h
    port map (
            O => \N__56456\,
            I => \N__56438\
        );

    \I__12156\ : Span4Mux_v
    port map (
            O => \N__56453\,
            I => \N__56438\
        );

    \I__12155\ : Span4Mux_v
    port map (
            O => \N__56450\,
            I => \N__56438\
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__56445\,
            I => \N__56435\
        );

    \I__12153\ : Span4Mux_h
    port map (
            O => \N__56438\,
            I => \N__56432\
        );

    \I__12152\ : Odrv4
    port map (
            O => \N__56435\,
            I => \c0.n12_adj_4671\
        );

    \I__12151\ : Odrv4
    port map (
            O => \N__56432\,
            I => \c0.n12_adj_4671\
        );

    \I__12150\ : InMux
    port map (
            O => \N__56427\,
            I => \N__56424\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__56424\,
            I => \N__56421\
        );

    \I__12148\ : Odrv12
    port map (
            O => \N__56421\,
            I => \c0.n22_adj_4350\
        );

    \I__12147\ : CascadeMux
    port map (
            O => \N__56418\,
            I => \c0.n22_adj_4350_cascade_\
        );

    \I__12146\ : InMux
    port map (
            O => \N__56415\,
            I => \N__56412\
        );

    \I__12145\ : LocalMux
    port map (
            O => \N__56412\,
            I => \N__56408\
        );

    \I__12144\ : CascadeMux
    port map (
            O => \N__56411\,
            I => \N__56403\
        );

    \I__12143\ : Span4Mux_h
    port map (
            O => \N__56408\,
            I => \N__56400\
        );

    \I__12142\ : CascadeMux
    port map (
            O => \N__56407\,
            I => \N__56397\
        );

    \I__12141\ : InMux
    port map (
            O => \N__56406\,
            I => \N__56393\
        );

    \I__12140\ : InMux
    port map (
            O => \N__56403\,
            I => \N__56390\
        );

    \I__12139\ : Span4Mux_v
    port map (
            O => \N__56400\,
            I => \N__56387\
        );

    \I__12138\ : InMux
    port map (
            O => \N__56397\,
            I => \N__56382\
        );

    \I__12137\ : InMux
    port map (
            O => \N__56396\,
            I => \N__56382\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__56393\,
            I => \c0.data_in_frame_20_6\
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__56390\,
            I => \c0.data_in_frame_20_6\
        );

    \I__12134\ : Odrv4
    port map (
            O => \N__56387\,
            I => \c0.data_in_frame_20_6\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__56382\,
            I => \c0.data_in_frame_20_6\
        );

    \I__12132\ : InMux
    port map (
            O => \N__56373\,
            I => \N__56366\
        );

    \I__12131\ : InMux
    port map (
            O => \N__56372\,
            I => \N__56361\
        );

    \I__12130\ : InMux
    port map (
            O => \N__56371\,
            I => \N__56361\
        );

    \I__12129\ : CascadeMux
    port map (
            O => \N__56370\,
            I => \N__56358\
        );

    \I__12128\ : InMux
    port map (
            O => \N__56369\,
            I => \N__56355\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__56366\,
            I => \N__56351\
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__56361\,
            I => \N__56348\
        );

    \I__12125\ : InMux
    port map (
            O => \N__56358\,
            I => \N__56345\
        );

    \I__12124\ : LocalMux
    port map (
            O => \N__56355\,
            I => \N__56342\
        );

    \I__12123\ : InMux
    port map (
            O => \N__56354\,
            I => \N__56339\
        );

    \I__12122\ : Span4Mux_h
    port map (
            O => \N__56351\,
            I => \N__56334\
        );

    \I__12121\ : Span4Mux_v
    port map (
            O => \N__56348\,
            I => \N__56334\
        );

    \I__12120\ : LocalMux
    port map (
            O => \N__56345\,
            I => \c0.data_in_frame_20_7\
        );

    \I__12119\ : Odrv12
    port map (
            O => \N__56342\,
            I => \c0.data_in_frame_20_7\
        );

    \I__12118\ : LocalMux
    port map (
            O => \N__56339\,
            I => \c0.data_in_frame_20_7\
        );

    \I__12117\ : Odrv4
    port map (
            O => \N__56334\,
            I => \c0.data_in_frame_20_7\
        );

    \I__12116\ : InMux
    port map (
            O => \N__56325\,
            I => \N__56317\
        );

    \I__12115\ : InMux
    port map (
            O => \N__56324\,
            I => \N__56317\
        );

    \I__12114\ : InMux
    port map (
            O => \N__56323\,
            I => \N__56312\
        );

    \I__12113\ : InMux
    port map (
            O => \N__56322\,
            I => \N__56312\
        );

    \I__12112\ : LocalMux
    port map (
            O => \N__56317\,
            I => \N__56309\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__56312\,
            I => \N__56306\
        );

    \I__12110\ : Span4Mux_v
    port map (
            O => \N__56309\,
            I => \N__56303\
        );

    \I__12109\ : Odrv4
    port map (
            O => \N__56306\,
            I => \c0.n21_adj_4225\
        );

    \I__12108\ : Odrv4
    port map (
            O => \N__56303\,
            I => \c0.n21_adj_4225\
        );

    \I__12107\ : CascadeMux
    port map (
            O => \N__56298\,
            I => \N__56295\
        );

    \I__12106\ : InMux
    port map (
            O => \N__56295\,
            I => \N__56292\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__56292\,
            I => \N__56289\
        );

    \I__12104\ : Span4Mux_h
    port map (
            O => \N__56289\,
            I => \N__56286\
        );

    \I__12103\ : Span4Mux_h
    port map (
            O => \N__56286\,
            I => \N__56283\
        );

    \I__12102\ : Odrv4
    port map (
            O => \N__56283\,
            I => \c0.n22227\
        );

    \I__12101\ : InMux
    port map (
            O => \N__56280\,
            I => \N__56277\
        );

    \I__12100\ : LocalMux
    port map (
            O => \N__56277\,
            I => \N__56273\
        );

    \I__12099\ : InMux
    port map (
            O => \N__56276\,
            I => \N__56269\
        );

    \I__12098\ : Span4Mux_h
    port map (
            O => \N__56273\,
            I => \N__56265\
        );

    \I__12097\ : InMux
    port map (
            O => \N__56272\,
            I => \N__56262\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__56269\,
            I => \N__56259\
        );

    \I__12095\ : InMux
    port map (
            O => \N__56268\,
            I => \N__56256\
        );

    \I__12094\ : Odrv4
    port map (
            O => \N__56265\,
            I => \c0.n23863\
        );

    \I__12093\ : LocalMux
    port map (
            O => \N__56262\,
            I => \c0.n23863\
        );

    \I__12092\ : Odrv4
    port map (
            O => \N__56259\,
            I => \c0.n23863\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__56256\,
            I => \c0.n23863\
        );

    \I__12090\ : InMux
    port map (
            O => \N__56247\,
            I => \N__56244\
        );

    \I__12089\ : LocalMux
    port map (
            O => \N__56244\,
            I => \c0.n160\
        );

    \I__12088\ : InMux
    port map (
            O => \N__56241\,
            I => \N__56236\
        );

    \I__12087\ : InMux
    port map (
            O => \N__56240\,
            I => \N__56233\
        );

    \I__12086\ : InMux
    port map (
            O => \N__56239\,
            I => \N__56230\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__56236\,
            I => \N__56227\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__56233\,
            I => \N__56224\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__56230\,
            I => \N__56220\
        );

    \I__12082\ : Span4Mux_h
    port map (
            O => \N__56227\,
            I => \N__56217\
        );

    \I__12081\ : Span4Mux_h
    port map (
            O => \N__56224\,
            I => \N__56214\
        );

    \I__12080\ : InMux
    port map (
            O => \N__56223\,
            I => \N__56211\
        );

    \I__12079\ : Span4Mux_v
    port map (
            O => \N__56220\,
            I => \N__56208\
        );

    \I__12078\ : Span4Mux_v
    port map (
            O => \N__56217\,
            I => \N__56203\
        );

    \I__12077\ : Span4Mux_v
    port map (
            O => \N__56214\,
            I => \N__56203\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__56211\,
            I => \c0.n12989\
        );

    \I__12075\ : Odrv4
    port map (
            O => \N__56208\,
            I => \c0.n12989\
        );

    \I__12074\ : Odrv4
    port map (
            O => \N__56203\,
            I => \c0.n12989\
        );

    \I__12073\ : CascadeMux
    port map (
            O => \N__56196\,
            I => \c0.n22104_cascade_\
        );

    \I__12072\ : InMux
    port map (
            O => \N__56193\,
            I => \N__56189\
        );

    \I__12071\ : InMux
    port map (
            O => \N__56192\,
            I => \N__56186\
        );

    \I__12070\ : LocalMux
    port map (
            O => \N__56189\,
            I => \N__56182\
        );

    \I__12069\ : LocalMux
    port map (
            O => \N__56186\,
            I => \N__56179\
        );

    \I__12068\ : InMux
    port map (
            O => \N__56185\,
            I => \N__56176\
        );

    \I__12067\ : Span4Mux_v
    port map (
            O => \N__56182\,
            I => \N__56171\
        );

    \I__12066\ : Span4Mux_h
    port map (
            O => \N__56179\,
            I => \N__56171\
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__56176\,
            I => \c0.data_in_frame_19_4\
        );

    \I__12064\ : Odrv4
    port map (
            O => \N__56171\,
            I => \c0.data_in_frame_19_4\
        );

    \I__12063\ : CascadeMux
    port map (
            O => \N__56166\,
            I => \c0.n22347_cascade_\
        );

    \I__12062\ : InMux
    port map (
            O => \N__56163\,
            I => \N__56160\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__56160\,
            I => \N__56156\
        );

    \I__12060\ : InMux
    port map (
            O => \N__56159\,
            I => \N__56153\
        );

    \I__12059\ : Odrv4
    port map (
            O => \N__56156\,
            I => \c0.n24520\
        );

    \I__12058\ : LocalMux
    port map (
            O => \N__56153\,
            I => \c0.n24520\
        );

    \I__12057\ : InMux
    port map (
            O => \N__56148\,
            I => \N__56144\
        );

    \I__12056\ : InMux
    port map (
            O => \N__56147\,
            I => \N__56140\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__56144\,
            I => \N__56136\
        );

    \I__12054\ : InMux
    port map (
            O => \N__56143\,
            I => \N__56133\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__56140\,
            I => \N__56130\
        );

    \I__12052\ : InMux
    port map (
            O => \N__56139\,
            I => \N__56127\
        );

    \I__12051\ : Span4Mux_v
    port map (
            O => \N__56136\,
            I => \N__56124\
        );

    \I__12050\ : LocalMux
    port map (
            O => \N__56133\,
            I => \N__56119\
        );

    \I__12049\ : Span4Mux_v
    port map (
            O => \N__56130\,
            I => \N__56119\
        );

    \I__12048\ : LocalMux
    port map (
            O => \N__56127\,
            I => \c0.data_in_frame_20_5\
        );

    \I__12047\ : Odrv4
    port map (
            O => \N__56124\,
            I => \c0.data_in_frame_20_5\
        );

    \I__12046\ : Odrv4
    port map (
            O => \N__56119\,
            I => \c0.data_in_frame_20_5\
        );

    \I__12045\ : InMux
    port map (
            O => \N__56112\,
            I => \N__56109\
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__56109\,
            I => \N__56106\
        );

    \I__12043\ : Odrv4
    port map (
            O => \N__56106\,
            I => \c0.n33\
        );

    \I__12042\ : CascadeMux
    port map (
            O => \N__56103\,
            I => \c0.n34_adj_4600_cascade_\
        );

    \I__12041\ : InMux
    port map (
            O => \N__56100\,
            I => \N__56097\
        );

    \I__12040\ : LocalMux
    port map (
            O => \N__56097\,
            I => \N__56094\
        );

    \I__12039\ : Span4Mux_v
    port map (
            O => \N__56094\,
            I => \N__56091\
        );

    \I__12038\ : Odrv4
    port map (
            O => \N__56091\,
            I => \c0.n38_adj_4573\
        );

    \I__12037\ : CascadeMux
    port map (
            O => \N__56088\,
            I => \c0.n24333_cascade_\
        );

    \I__12036\ : InMux
    port map (
            O => \N__56085\,
            I => \N__56079\
        );

    \I__12035\ : InMux
    port map (
            O => \N__56084\,
            I => \N__56079\
        );

    \I__12034\ : LocalMux
    port map (
            O => \N__56079\,
            I => \N__56076\
        );

    \I__12033\ : Odrv4
    port map (
            O => \N__56076\,
            I => \c0.n23661\
        );

    \I__12032\ : CascadeMux
    port map (
            O => \N__56073\,
            I => \N__56069\
        );

    \I__12031\ : CascadeMux
    port map (
            O => \N__56072\,
            I => \N__56066\
        );

    \I__12030\ : InMux
    port map (
            O => \N__56069\,
            I => \N__56063\
        );

    \I__12029\ : InMux
    port map (
            O => \N__56066\,
            I => \N__56060\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__56063\,
            I => \N__56057\
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__56060\,
            I => \N__56051\
        );

    \I__12026\ : Span4Mux_h
    port map (
            O => \N__56057\,
            I => \N__56051\
        );

    \I__12025\ : InMux
    port map (
            O => \N__56056\,
            I => \N__56048\
        );

    \I__12024\ : Odrv4
    port map (
            O => \N__56051\,
            I => \c0.data_in_frame_18_5\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__56048\,
            I => \c0.data_in_frame_18_5\
        );

    \I__12022\ : InMux
    port map (
            O => \N__56043\,
            I => \N__56040\
        );

    \I__12021\ : LocalMux
    port map (
            O => \N__56040\,
            I => \N__56035\
        );

    \I__12020\ : InMux
    port map (
            O => \N__56039\,
            I => \N__56030\
        );

    \I__12019\ : InMux
    port map (
            O => \N__56038\,
            I => \N__56030\
        );

    \I__12018\ : Span4Mux_h
    port map (
            O => \N__56035\,
            I => \N__56027\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__56030\,
            I => \c0.data_in_frame_16_3\
        );

    \I__12016\ : Odrv4
    port map (
            O => \N__56027\,
            I => \c0.data_in_frame_16_3\
        );

    \I__12015\ : InMux
    port map (
            O => \N__56022\,
            I => \N__56019\
        );

    \I__12014\ : LocalMux
    port map (
            O => \N__56019\,
            I => \N__56016\
        );

    \I__12013\ : Odrv12
    port map (
            O => \N__56016\,
            I => \c0.n155\
        );

    \I__12012\ : InMux
    port map (
            O => \N__56013\,
            I => \N__56010\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__56010\,
            I => \N__56006\
        );

    \I__12010\ : CascadeMux
    port map (
            O => \N__56009\,
            I => \N__56002\
        );

    \I__12009\ : Span4Mux_v
    port map (
            O => \N__56006\,
            I => \N__55999\
        );

    \I__12008\ : InMux
    port map (
            O => \N__56005\,
            I => \N__55994\
        );

    \I__12007\ : InMux
    port map (
            O => \N__56002\,
            I => \N__55994\
        );

    \I__12006\ : Span4Mux_v
    port map (
            O => \N__55999\,
            I => \N__55991\
        );

    \I__12005\ : LocalMux
    port map (
            O => \N__55994\,
            I => \N__55988\
        );

    \I__12004\ : Odrv4
    port map (
            O => \N__55991\,
            I => \c0.n5_adj_4311\
        );

    \I__12003\ : Odrv4
    port map (
            O => \N__55988\,
            I => \c0.n5_adj_4311\
        );

    \I__12002\ : CascadeMux
    port map (
            O => \N__55983\,
            I => \c0.n5_adj_4311_cascade_\
        );

    \I__12001\ : InMux
    port map (
            O => \N__55980\,
            I => \N__55977\
        );

    \I__12000\ : LocalMux
    port map (
            O => \N__55977\,
            I => \N__55973\
        );

    \I__11999\ : InMux
    port map (
            O => \N__55976\,
            I => \N__55969\
        );

    \I__11998\ : Span4Mux_h
    port map (
            O => \N__55973\,
            I => \N__55966\
        );

    \I__11997\ : InMux
    port map (
            O => \N__55972\,
            I => \N__55962\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__55969\,
            I => \N__55959\
        );

    \I__11995\ : Span4Mux_v
    port map (
            O => \N__55966\,
            I => \N__55956\
        );

    \I__11994\ : InMux
    port map (
            O => \N__55965\,
            I => \N__55953\
        );

    \I__11993\ : LocalMux
    port map (
            O => \N__55962\,
            I => \c0.data_in_frame_10_3\
        );

    \I__11992\ : Odrv4
    port map (
            O => \N__55959\,
            I => \c0.data_in_frame_10_3\
        );

    \I__11991\ : Odrv4
    port map (
            O => \N__55956\,
            I => \c0.data_in_frame_10_3\
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__55953\,
            I => \c0.data_in_frame_10_3\
        );

    \I__11989\ : InMux
    port map (
            O => \N__55944\,
            I => \N__55938\
        );

    \I__11988\ : InMux
    port map (
            O => \N__55943\,
            I => \N__55938\
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__55938\,
            I => \N__55935\
        );

    \I__11986\ : Odrv12
    port map (
            O => \N__55935\,
            I => \c0.n23677\
        );

    \I__11985\ : CascadeMux
    port map (
            O => \N__55932\,
            I => \N__55928\
        );

    \I__11984\ : InMux
    port map (
            O => \N__55931\,
            I => \N__55923\
        );

    \I__11983\ : InMux
    port map (
            O => \N__55928\,
            I => \N__55923\
        );

    \I__11982\ : LocalMux
    port map (
            O => \N__55923\,
            I => \N__55920\
        );

    \I__11981\ : Span4Mux_h
    port map (
            O => \N__55920\,
            I => \N__55916\
        );

    \I__11980\ : InMux
    port map (
            O => \N__55919\,
            I => \N__55913\
        );

    \I__11979\ : Span4Mux_v
    port map (
            O => \N__55916\,
            I => \N__55910\
        );

    \I__11978\ : LocalMux
    port map (
            O => \N__55913\,
            I => data_in_frame_14_4
        );

    \I__11977\ : Odrv4
    port map (
            O => \N__55910\,
            I => data_in_frame_14_4
        );

    \I__11976\ : CascadeMux
    port map (
            O => \N__55905\,
            I => \N__55902\
        );

    \I__11975\ : InMux
    port map (
            O => \N__55902\,
            I => \N__55889\
        );

    \I__11974\ : InMux
    port map (
            O => \N__55901\,
            I => \N__55889\
        );

    \I__11973\ : InMux
    port map (
            O => \N__55900\,
            I => \N__55889\
        );

    \I__11972\ : InMux
    port map (
            O => \N__55899\,
            I => \N__55889\
        );

    \I__11971\ : CascadeMux
    port map (
            O => \N__55898\,
            I => \N__55886\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__55889\,
            I => \N__55883\
        );

    \I__11969\ : InMux
    port map (
            O => \N__55886\,
            I => \N__55879\
        );

    \I__11968\ : Span4Mux_h
    port map (
            O => \N__55883\,
            I => \N__55876\
        );

    \I__11967\ : InMux
    port map (
            O => \N__55882\,
            I => \N__55873\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__55879\,
            I => \c0.data_in_frame_8_2\
        );

    \I__11965\ : Odrv4
    port map (
            O => \N__55876\,
            I => \c0.data_in_frame_8_2\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__55873\,
            I => \c0.data_in_frame_8_2\
        );

    \I__11963\ : CascadeMux
    port map (
            O => \N__55866\,
            I => \c0.n120_cascade_\
        );

    \I__11962\ : InMux
    port map (
            O => \N__55863\,
            I => \N__55860\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__55860\,
            I => \N__55857\
        );

    \I__11960\ : Span4Mux_v
    port map (
            O => \N__55857\,
            I => \N__55854\
        );

    \I__11959\ : Odrv4
    port map (
            O => \N__55854\,
            I => \c0.n142\
        );

    \I__11958\ : CascadeMux
    port map (
            O => \N__55851\,
            I => \c0.n152_cascade_\
        );

    \I__11957\ : InMux
    port map (
            O => \N__55848\,
            I => \N__55845\
        );

    \I__11956\ : LocalMux
    port map (
            O => \N__55845\,
            I => \N__55842\
        );

    \I__11955\ : Odrv4
    port map (
            O => \N__55842\,
            I => \c0.n158\
        );

    \I__11954\ : InMux
    port map (
            O => \N__55839\,
            I => \N__55835\
        );

    \I__11953\ : InMux
    port map (
            O => \N__55838\,
            I => \N__55832\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__55835\,
            I => \N__55827\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__55832\,
            I => \N__55827\
        );

    \I__11950\ : Odrv12
    port map (
            O => \N__55827\,
            I => \c0.n22472\
        );

    \I__11949\ : InMux
    port map (
            O => \N__55824\,
            I => \N__55820\
        );

    \I__11948\ : CascadeMux
    port map (
            O => \N__55823\,
            I => \N__55817\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__55820\,
            I => \N__55814\
        );

    \I__11946\ : InMux
    port map (
            O => \N__55817\,
            I => \N__55811\
        );

    \I__11945\ : Span4Mux_h
    port map (
            O => \N__55814\,
            I => \N__55808\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__55811\,
            I => data_in_frame_14_3
        );

    \I__11943\ : Odrv4
    port map (
            O => \N__55808\,
            I => data_in_frame_14_3
        );

    \I__11942\ : CascadeMux
    port map (
            O => \N__55803\,
            I => \c0.n30_adj_4571_cascade_\
        );

    \I__11941\ : InMux
    port map (
            O => \N__55800\,
            I => \N__55790\
        );

    \I__11940\ : InMux
    port map (
            O => \N__55799\,
            I => \N__55790\
        );

    \I__11939\ : InMux
    port map (
            O => \N__55798\,
            I => \N__55790\
        );

    \I__11938\ : InMux
    port map (
            O => \N__55797\,
            I => \N__55787\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__55790\,
            I => \N__55782\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__55787\,
            I => \N__55782\
        );

    \I__11935\ : Odrv4
    port map (
            O => \N__55782\,
            I => \c0.data_in_frame_4_1\
        );

    \I__11934\ : CascadeMux
    port map (
            O => \N__55779\,
            I => \N__55776\
        );

    \I__11933\ : InMux
    port map (
            O => \N__55776\,
            I => \N__55770\
        );

    \I__11932\ : InMux
    port map (
            O => \N__55775\,
            I => \N__55770\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__55770\,
            I => \c0.data_in_frame_10_4\
        );

    \I__11930\ : InMux
    port map (
            O => \N__55767\,
            I => \N__55761\
        );

    \I__11929\ : InMux
    port map (
            O => \N__55766\,
            I => \N__55761\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__55761\,
            I => \N__55757\
        );

    \I__11927\ : InMux
    port map (
            O => \N__55760\,
            I => \N__55754\
        );

    \I__11926\ : Span4Mux_h
    port map (
            O => \N__55757\,
            I => \N__55751\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__55754\,
            I => \c0.n22455\
        );

    \I__11924\ : Odrv4
    port map (
            O => \N__55751\,
            I => \c0.n22455\
        );

    \I__11923\ : CascadeMux
    port map (
            O => \N__55746\,
            I => \N__55743\
        );

    \I__11922\ : InMux
    port map (
            O => \N__55743\,
            I => \N__55737\
        );

    \I__11921\ : CascadeMux
    port map (
            O => \N__55742\,
            I => \N__55734\
        );

    \I__11920\ : InMux
    port map (
            O => \N__55741\,
            I => \N__55731\
        );

    \I__11919\ : InMux
    port map (
            O => \N__55740\,
            I => \N__55728\
        );

    \I__11918\ : LocalMux
    port map (
            O => \N__55737\,
            I => \N__55724\
        );

    \I__11917\ : InMux
    port map (
            O => \N__55734\,
            I => \N__55721\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__55731\,
            I => \N__55718\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__55728\,
            I => \N__55715\
        );

    \I__11914\ : InMux
    port map (
            O => \N__55727\,
            I => \N__55712\
        );

    \I__11913\ : Span4Mux_h
    port map (
            O => \N__55724\,
            I => \N__55709\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__55721\,
            I => \N__55704\
        );

    \I__11911\ : Span4Mux_v
    port map (
            O => \N__55718\,
            I => \N__55704\
        );

    \I__11910\ : Span4Mux_h
    port map (
            O => \N__55715\,
            I => \N__55701\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__55712\,
            I => \N__55698\
        );

    \I__11908\ : Span4Mux_v
    port map (
            O => \N__55709\,
            I => \N__55695\
        );

    \I__11907\ : Odrv4
    port map (
            O => \N__55704\,
            I => \c0.data_in_frame_12_5\
        );

    \I__11906\ : Odrv4
    port map (
            O => \N__55701\,
            I => \c0.data_in_frame_12_5\
        );

    \I__11905\ : Odrv4
    port map (
            O => \N__55698\,
            I => \c0.data_in_frame_12_5\
        );

    \I__11904\ : Odrv4
    port map (
            O => \N__55695\,
            I => \c0.data_in_frame_12_5\
        );

    \I__11903\ : InMux
    port map (
            O => \N__55686\,
            I => \N__55683\
        );

    \I__11902\ : LocalMux
    port map (
            O => \N__55683\,
            I => \N__55679\
        );

    \I__11901\ : CascadeMux
    port map (
            O => \N__55682\,
            I => \N__55676\
        );

    \I__11900\ : Span4Mux_h
    port map (
            O => \N__55679\,
            I => \N__55673\
        );

    \I__11899\ : InMux
    port map (
            O => \N__55676\,
            I => \N__55670\
        );

    \I__11898\ : Sp12to4
    port map (
            O => \N__55673\,
            I => \N__55665\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__55670\,
            I => \N__55665\
        );

    \I__11896\ : Span12Mux_v
    port map (
            O => \N__55665\,
            I => \N__55661\
        );

    \I__11895\ : InMux
    port map (
            O => \N__55664\,
            I => \N__55658\
        );

    \I__11894\ : Odrv12
    port map (
            O => \N__55661\,
            I => \c0.n42\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__55658\,
            I => \c0.n42\
        );

    \I__11892\ : InMux
    port map (
            O => \N__55653\,
            I => \N__55650\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__55650\,
            I => \N__55647\
        );

    \I__11890\ : Odrv4
    port map (
            O => \N__55647\,
            I => \c0.n58\
        );

    \I__11889\ : InMux
    port map (
            O => \N__55644\,
            I => \N__55641\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__55641\,
            I => \N__55638\
        );

    \I__11887\ : Odrv4
    port map (
            O => \N__55638\,
            I => \c0.n127\
        );

    \I__11886\ : CascadeMux
    port map (
            O => \N__55635\,
            I => \c0.n41_adj_4452_cascade_\
        );

    \I__11885\ : InMux
    port map (
            O => \N__55632\,
            I => \N__55627\
        );

    \I__11884\ : InMux
    port map (
            O => \N__55631\,
            I => \N__55624\
        );

    \I__11883\ : InMux
    port map (
            O => \N__55630\,
            I => \N__55621\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__55627\,
            I => \N__55618\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__55624\,
            I => \N__55615\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__55621\,
            I => \N__55612\
        );

    \I__11879\ : Span4Mux_h
    port map (
            O => \N__55618\,
            I => \N__55604\
        );

    \I__11878\ : Span4Mux_v
    port map (
            O => \N__55615\,
            I => \N__55604\
        );

    \I__11877\ : Span4Mux_v
    port map (
            O => \N__55612\,
            I => \N__55604\
        );

    \I__11876\ : InMux
    port map (
            O => \N__55611\,
            I => \N__55601\
        );

    \I__11875\ : Span4Mux_h
    port map (
            O => \N__55604\,
            I => \N__55598\
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__55601\,
            I => \c0.data_in_frame_11_7\
        );

    \I__11873\ : Odrv4
    port map (
            O => \N__55598\,
            I => \c0.data_in_frame_11_7\
        );

    \I__11872\ : InMux
    port map (
            O => \N__55593\,
            I => \N__55590\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__55590\,
            I => \c0.n39_adj_4453\
        );

    \I__11870\ : InMux
    port map (
            O => \N__55587\,
            I => \N__55584\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__55584\,
            I => \c0.n40_adj_4451\
        );

    \I__11868\ : CascadeMux
    port map (
            O => \N__55581\,
            I => \N__55578\
        );

    \I__11867\ : InMux
    port map (
            O => \N__55578\,
            I => \N__55575\
        );

    \I__11866\ : LocalMux
    port map (
            O => \N__55575\,
            I => \N__55572\
        );

    \I__11865\ : Span4Mux_h
    port map (
            O => \N__55572\,
            I => \N__55569\
        );

    \I__11864\ : Odrv4
    port map (
            O => \N__55569\,
            I => \c0.n14016\
        );

    \I__11863\ : InMux
    port map (
            O => \N__55566\,
            I => \N__55561\
        );

    \I__11862\ : InMux
    port map (
            O => \N__55565\,
            I => \N__55558\
        );

    \I__11861\ : CascadeMux
    port map (
            O => \N__55564\,
            I => \N__55555\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__55561\,
            I => \N__55552\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__55558\,
            I => \N__55549\
        );

    \I__11858\ : InMux
    port map (
            O => \N__55555\,
            I => \N__55546\
        );

    \I__11857\ : Span4Mux_v
    port map (
            O => \N__55552\,
            I => \N__55543\
        );

    \I__11856\ : Span4Mux_v
    port map (
            O => \N__55549\,
            I => \N__55538\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__55546\,
            I => \N__55538\
        );

    \I__11854\ : Odrv4
    port map (
            O => \N__55543\,
            I => \c0.n13223\
        );

    \I__11853\ : Odrv4
    port map (
            O => \N__55538\,
            I => \c0.n13223\
        );

    \I__11852\ : InMux
    port map (
            O => \N__55533\,
            I => \N__55530\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__55530\,
            I => \N__55527\
        );

    \I__11850\ : Odrv4
    port map (
            O => \N__55527\,
            I => \c0.n16_adj_4608\
        );

    \I__11849\ : InMux
    port map (
            O => \N__55524\,
            I => \N__55520\
        );

    \I__11848\ : InMux
    port map (
            O => \N__55523\,
            I => \N__55517\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__55520\,
            I => \N__55514\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__55517\,
            I => \N__55509\
        );

    \I__11845\ : Span4Mux_h
    port map (
            O => \N__55514\,
            I => \N__55505\
        );

    \I__11844\ : InMux
    port map (
            O => \N__55513\,
            I => \N__55500\
        );

    \I__11843\ : InMux
    port map (
            O => \N__55512\,
            I => \N__55500\
        );

    \I__11842\ : Span12Mux_v
    port map (
            O => \N__55509\,
            I => \N__55497\
        );

    \I__11841\ : InMux
    port map (
            O => \N__55508\,
            I => \N__55494\
        );

    \I__11840\ : Sp12to4
    port map (
            O => \N__55505\,
            I => \N__55489\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__55500\,
            I => \N__55489\
        );

    \I__11838\ : Odrv12
    port map (
            O => \N__55497\,
            I => \c0.n21\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__55494\,
            I => \c0.n21\
        );

    \I__11836\ : Odrv12
    port map (
            O => \N__55489\,
            I => \c0.n21\
        );

    \I__11835\ : CascadeMux
    port map (
            O => \N__55482\,
            I => \N__55479\
        );

    \I__11834\ : InMux
    port map (
            O => \N__55479\,
            I => \N__55475\
        );

    \I__11833\ : InMux
    port map (
            O => \N__55478\,
            I => \N__55472\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__55475\,
            I => \N__55469\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__55472\,
            I => \N__55466\
        );

    \I__11830\ : Span4Mux_h
    port map (
            O => \N__55469\,
            I => \N__55463\
        );

    \I__11829\ : Span4Mux_h
    port map (
            O => \N__55466\,
            I => \N__55460\
        );

    \I__11828\ : Odrv4
    port map (
            O => \N__55463\,
            I => \c0.n20\
        );

    \I__11827\ : Odrv4
    port map (
            O => \N__55460\,
            I => \c0.n20\
        );

    \I__11826\ : InMux
    port map (
            O => \N__55455\,
            I => \N__55451\
        );

    \I__11825\ : InMux
    port map (
            O => \N__55454\,
            I => \N__55448\
        );

    \I__11824\ : LocalMux
    port map (
            O => \N__55451\,
            I => \N__55445\
        );

    \I__11823\ : LocalMux
    port map (
            O => \N__55448\,
            I => \N__55442\
        );

    \I__11822\ : Span4Mux_v
    port map (
            O => \N__55445\,
            I => \N__55439\
        );

    \I__11821\ : Odrv12
    port map (
            O => \N__55442\,
            I => \c0.n13_adj_4610\
        );

    \I__11820\ : Odrv4
    port map (
            O => \N__55439\,
            I => \c0.n13_adj_4610\
        );

    \I__11819\ : InMux
    port map (
            O => \N__55434\,
            I => \N__55431\
        );

    \I__11818\ : LocalMux
    port map (
            O => \N__55431\,
            I => \N__55426\
        );

    \I__11817\ : InMux
    port map (
            O => \N__55430\,
            I => \N__55423\
        );

    \I__11816\ : InMux
    port map (
            O => \N__55429\,
            I => \N__55420\
        );

    \I__11815\ : Span4Mux_h
    port map (
            O => \N__55426\,
            I => \N__55415\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__55423\,
            I => \N__55415\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__55420\,
            I => data_in_frame_14_1
        );

    \I__11812\ : Odrv4
    port map (
            O => \N__55415\,
            I => data_in_frame_14_1
        );

    \I__11811\ : InMux
    port map (
            O => \N__55410\,
            I => \N__55407\
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__55407\,
            I => \N__55404\
        );

    \I__11809\ : Odrv4
    port map (
            O => \N__55404\,
            I => \c0.n102\
        );

    \I__11808\ : CascadeMux
    port map (
            O => \N__55401\,
            I => \c0.n147_cascade_\
        );

    \I__11807\ : InMux
    port map (
            O => \N__55398\,
            I => \N__55395\
        );

    \I__11806\ : LocalMux
    port map (
            O => \N__55395\,
            I => \c0.n134\
        );

    \I__11805\ : CascadeMux
    port map (
            O => \N__55392\,
            I => \N__55389\
        );

    \I__11804\ : InMux
    port map (
            O => \N__55389\,
            I => \N__55386\
        );

    \I__11803\ : LocalMux
    port map (
            O => \N__55386\,
            I => \c0.n131\
        );

    \I__11802\ : CascadeMux
    port map (
            O => \N__55383\,
            I => \N__55380\
        );

    \I__11801\ : InMux
    port map (
            O => \N__55380\,
            I => \N__55377\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__55377\,
            I => \N__55374\
        );

    \I__11799\ : Span4Mux_h
    port map (
            O => \N__55374\,
            I => \N__55371\
        );

    \I__11798\ : Odrv4
    port map (
            O => \N__55371\,
            I => \c0.n31_adj_4284\
        );

    \I__11797\ : InMux
    port map (
            O => \N__55368\,
            I => \N__55365\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__55365\,
            I => \c0.n36_adj_4447\
        );

    \I__11795\ : InMux
    port map (
            O => \N__55362\,
            I => \N__55359\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__55359\,
            I => \N__55356\
        );

    \I__11793\ : Span4Mux_v
    port map (
            O => \N__55356\,
            I => \N__55353\
        );

    \I__11792\ : Odrv4
    port map (
            O => \N__55353\,
            I => \c0.n5_adj_4268\
        );

    \I__11791\ : InMux
    port map (
            O => \N__55350\,
            I => \N__55347\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__55347\,
            I => \N__55344\
        );

    \I__11789\ : Span4Mux_h
    port map (
            O => \N__55344\,
            I => \N__55341\
        );

    \I__11788\ : Odrv4
    port map (
            O => \N__55341\,
            I => \c0.n4_adj_4267\
        );

    \I__11787\ : InMux
    port map (
            O => \N__55338\,
            I => \N__55335\
        );

    \I__11786\ : LocalMux
    port map (
            O => \N__55335\,
            I => \c0.n4_adj_4269\
        );

    \I__11785\ : InMux
    port map (
            O => \N__55332\,
            I => \N__55326\
        );

    \I__11784\ : InMux
    port map (
            O => \N__55331\,
            I => \N__55323\
        );

    \I__11783\ : InMux
    port map (
            O => \N__55330\,
            I => \N__55319\
        );

    \I__11782\ : CascadeMux
    port map (
            O => \N__55329\,
            I => \N__55316\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__55326\,
            I => \N__55311\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__55323\,
            I => \N__55311\
        );

    \I__11779\ : InMux
    port map (
            O => \N__55322\,
            I => \N__55308\
        );

    \I__11778\ : LocalMux
    port map (
            O => \N__55319\,
            I => \N__55305\
        );

    \I__11777\ : InMux
    port map (
            O => \N__55316\,
            I => \N__55302\
        );

    \I__11776\ : Span4Mux_v
    port map (
            O => \N__55311\,
            I => \N__55297\
        );

    \I__11775\ : LocalMux
    port map (
            O => \N__55308\,
            I => \N__55297\
        );

    \I__11774\ : Odrv4
    port map (
            O => \N__55305\,
            I => \c0.n22196\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__55302\,
            I => \c0.n22196\
        );

    \I__11772\ : Odrv4
    port map (
            O => \N__55297\,
            I => \c0.n22196\
        );

    \I__11771\ : CascadeMux
    port map (
            O => \N__55290\,
            I => \c0.n4_adj_4269_cascade_\
        );

    \I__11770\ : InMux
    port map (
            O => \N__55287\,
            I => \N__55284\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__55284\,
            I => \c0.n68\
        );

    \I__11768\ : CascadeMux
    port map (
            O => \N__55281\,
            I => \c0.n89_cascade_\
        );

    \I__11767\ : CascadeMux
    port map (
            O => \N__55278\,
            I => \c0.n23_cascade_\
        );

    \I__11766\ : CascadeMux
    port map (
            O => \N__55275\,
            I => \N__55272\
        );

    \I__11765\ : InMux
    port map (
            O => \N__55272\,
            I => \N__55269\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__55269\,
            I => \N__55266\
        );

    \I__11763\ : Span4Mux_v
    port map (
            O => \N__55266\,
            I => \N__55263\
        );

    \I__11762\ : Span4Mux_v
    port map (
            O => \N__55263\,
            I => \N__55260\
        );

    \I__11761\ : Odrv4
    port map (
            O => \N__55260\,
            I => \c0.n26\
        );

    \I__11760\ : CascadeMux
    port map (
            O => \N__55257\,
            I => \c0.n13075_cascade_\
        );

    \I__11759\ : CascadeMux
    port map (
            O => \N__55254\,
            I => \c0.n93_cascade_\
        );

    \I__11758\ : InMux
    port map (
            O => \N__55251\,
            I => \N__55248\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__55248\,
            I => \c0.n12_adj_4299\
        );

    \I__11756\ : CascadeMux
    port map (
            O => \N__55245\,
            I => \c0.n7_adj_4300_cascade_\
        );

    \I__11755\ : InMux
    port map (
            O => \N__55242\,
            I => \N__55238\
        );

    \I__11754\ : CascadeMux
    port map (
            O => \N__55241\,
            I => \N__55235\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__55238\,
            I => \N__55232\
        );

    \I__11752\ : InMux
    port map (
            O => \N__55235\,
            I => \N__55229\
        );

    \I__11751\ : Span4Mux_v
    port map (
            O => \N__55232\,
            I => \N__55226\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__55229\,
            I => \c0.n11_adj_4280\
        );

    \I__11749\ : Odrv4
    port map (
            O => \N__55226\,
            I => \c0.n11_adj_4280\
        );

    \I__11748\ : InMux
    port map (
            O => \N__55221\,
            I => \N__55217\
        );

    \I__11747\ : InMux
    port map (
            O => \N__55220\,
            I => \N__55214\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__55217\,
            I => \N__55211\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__55214\,
            I => \N__55208\
        );

    \I__11744\ : Span4Mux_h
    port map (
            O => \N__55211\,
            I => \N__55203\
        );

    \I__11743\ : Span4Mux_h
    port map (
            O => \N__55208\,
            I => \N__55200\
        );

    \I__11742\ : InMux
    port map (
            O => \N__55207\,
            I => \N__55195\
        );

    \I__11741\ : InMux
    port map (
            O => \N__55206\,
            I => \N__55195\
        );

    \I__11740\ : Odrv4
    port map (
            O => \N__55203\,
            I => \c0.n23251\
        );

    \I__11739\ : Odrv4
    port map (
            O => \N__55200\,
            I => \c0.n23251\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__55195\,
            I => \c0.n23251\
        );

    \I__11737\ : InMux
    port map (
            O => \N__55188\,
            I => \N__55179\
        );

    \I__11736\ : InMux
    port map (
            O => \N__55187\,
            I => \N__55179\
        );

    \I__11735\ : InMux
    port map (
            O => \N__55186\,
            I => \N__55174\
        );

    \I__11734\ : InMux
    port map (
            O => \N__55185\,
            I => \N__55174\
        );

    \I__11733\ : InMux
    port map (
            O => \N__55184\,
            I => \N__55171\
        );

    \I__11732\ : LocalMux
    port map (
            O => \N__55179\,
            I => \N__55168\
        );

    \I__11731\ : LocalMux
    port map (
            O => \N__55174\,
            I => \N__55165\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__55171\,
            I => \N__55162\
        );

    \I__11729\ : Span4Mux_h
    port map (
            O => \N__55168\,
            I => \N__55157\
        );

    \I__11728\ : Span4Mux_v
    port map (
            O => \N__55165\,
            I => \N__55157\
        );

    \I__11727\ : Odrv4
    port map (
            O => \N__55162\,
            I => \c0.n23305\
        );

    \I__11726\ : Odrv4
    port map (
            O => \N__55157\,
            I => \c0.n23305\
        );

    \I__11725\ : CascadeMux
    port map (
            O => \N__55152\,
            I => \c0.n23251_cascade_\
        );

    \I__11724\ : InMux
    port map (
            O => \N__55149\,
            I => \N__55146\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__55146\,
            I => \N__55143\
        );

    \I__11722\ : Span4Mux_v
    port map (
            O => \N__55143\,
            I => \N__55140\
        );

    \I__11721\ : Odrv4
    port map (
            O => \N__55140\,
            I => \c0.n23574\
        );

    \I__11720\ : CascadeMux
    port map (
            O => \N__55137\,
            I => \c0.n7_adj_4282_cascade_\
        );

    \I__11719\ : InMux
    port map (
            O => \N__55134\,
            I => \N__55128\
        );

    \I__11718\ : InMux
    port map (
            O => \N__55133\,
            I => \N__55128\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__55128\,
            I => \c0.n10_adj_4283\
        );

    \I__11716\ : InMux
    port map (
            O => \N__55125\,
            I => \N__55121\
        );

    \I__11715\ : InMux
    port map (
            O => \N__55124\,
            I => \N__55118\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__55121\,
            I => \N__55115\
        );

    \I__11713\ : LocalMux
    port map (
            O => \N__55118\,
            I => \N__55110\
        );

    \I__11712\ : Span4Mux_h
    port map (
            O => \N__55115\,
            I => \N__55107\
        );

    \I__11711\ : InMux
    port map (
            O => \N__55114\,
            I => \N__55104\
        );

    \I__11710\ : CascadeMux
    port map (
            O => \N__55113\,
            I => \N__55101\
        );

    \I__11709\ : Span4Mux_h
    port map (
            O => \N__55110\,
            I => \N__55097\
        );

    \I__11708\ : Span4Mux_v
    port map (
            O => \N__55107\,
            I => \N__55092\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__55104\,
            I => \N__55092\
        );

    \I__11706\ : InMux
    port map (
            O => \N__55101\,
            I => \N__55087\
        );

    \I__11705\ : InMux
    port map (
            O => \N__55100\,
            I => \N__55087\
        );

    \I__11704\ : Odrv4
    port map (
            O => \N__55097\,
            I => \c0.data_in_frame_8_1\
        );

    \I__11703\ : Odrv4
    port map (
            O => \N__55092\,
            I => \c0.data_in_frame_8_1\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__55087\,
            I => \c0.data_in_frame_8_1\
        );

    \I__11701\ : CascadeMux
    port map (
            O => \N__55080\,
            I => \c0.n13_adj_4638_cascade_\
        );

    \I__11700\ : InMux
    port map (
            O => \N__55077\,
            I => \N__55074\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__55074\,
            I => \N__55071\
        );

    \I__11698\ : Span4Mux_h
    port map (
            O => \N__55071\,
            I => \N__55066\
        );

    \I__11697\ : InMux
    port map (
            O => \N__55070\,
            I => \N__55063\
        );

    \I__11696\ : InMux
    port map (
            O => \N__55069\,
            I => \N__55060\
        );

    \I__11695\ : Span4Mux_h
    port map (
            O => \N__55066\,
            I => \N__55057\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__55063\,
            I => \c0.data_in_frame_10_1\
        );

    \I__11693\ : LocalMux
    port map (
            O => \N__55060\,
            I => \c0.data_in_frame_10_1\
        );

    \I__11692\ : Odrv4
    port map (
            O => \N__55057\,
            I => \c0.data_in_frame_10_1\
        );

    \I__11691\ : CascadeMux
    port map (
            O => \N__55050\,
            I => \N__55046\
        );

    \I__11690\ : InMux
    port map (
            O => \N__55049\,
            I => \N__55040\
        );

    \I__11689\ : InMux
    port map (
            O => \N__55046\,
            I => \N__55040\
        );

    \I__11688\ : CascadeMux
    port map (
            O => \N__55045\,
            I => \N__55037\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__55040\,
            I => \N__55034\
        );

    \I__11686\ : InMux
    port map (
            O => \N__55037\,
            I => \N__55031\
        );

    \I__11685\ : Span4Mux_v
    port map (
            O => \N__55034\,
            I => \N__55028\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__55031\,
            I => \c0.data_in_frame_10_2\
        );

    \I__11683\ : Odrv4
    port map (
            O => \N__55028\,
            I => \c0.data_in_frame_10_2\
        );

    \I__11682\ : CascadeMux
    port map (
            O => \N__55023\,
            I => \N__55017\
        );

    \I__11681\ : InMux
    port map (
            O => \N__55022\,
            I => \N__55014\
        );

    \I__11680\ : InMux
    port map (
            O => \N__55021\,
            I => \N__55009\
        );

    \I__11679\ : InMux
    port map (
            O => \N__55020\,
            I => \N__55009\
        );

    \I__11678\ : InMux
    port map (
            O => \N__55017\,
            I => \N__55006\
        );

    \I__11677\ : LocalMux
    port map (
            O => \N__55014\,
            I => \N__55003\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__55009\,
            I => \N__55000\
        );

    \I__11675\ : LocalMux
    port map (
            O => \N__55006\,
            I => \N__54995\
        );

    \I__11674\ : Span4Mux_v
    port map (
            O => \N__55003\,
            I => \N__54995\
        );

    \I__11673\ : Span4Mux_h
    port map (
            O => \N__55000\,
            I => \N__54992\
        );

    \I__11672\ : Odrv4
    port map (
            O => \N__54995\,
            I => \c0.data_in_frame_9_7\
        );

    \I__11671\ : Odrv4
    port map (
            O => \N__54992\,
            I => \c0.data_in_frame_9_7\
        );

    \I__11670\ : CascadeMux
    port map (
            O => \N__54987\,
            I => \c0.n22196_cascade_\
        );

    \I__11669\ : InMux
    port map (
            O => \N__54984\,
            I => \N__54981\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__54981\,
            I => \N__54978\
        );

    \I__11667\ : Span4Mux_h
    port map (
            O => \N__54978\,
            I => \N__54975\
        );

    \I__11666\ : Span4Mux_v
    port map (
            O => \N__54975\,
            I => \N__54972\
        );

    \I__11665\ : Odrv4
    port map (
            O => \N__54972\,
            I => \c0.n12_adj_4258\
        );

    \I__11664\ : InMux
    port map (
            O => \N__54969\,
            I => \N__54963\
        );

    \I__11663\ : InMux
    port map (
            O => \N__54968\,
            I => \N__54963\
        );

    \I__11662\ : LocalMux
    port map (
            O => \N__54963\,
            I => \c0.data_in_frame_3_0\
        );

    \I__11661\ : CascadeMux
    port map (
            O => \N__54960\,
            I => \N__54957\
        );

    \I__11660\ : InMux
    port map (
            O => \N__54957\,
            I => \N__54954\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__54954\,
            I => \c0.n10_adj_4615\
        );

    \I__11658\ : InMux
    port map (
            O => \N__54951\,
            I => \N__54947\
        );

    \I__11657\ : CascadeMux
    port map (
            O => \N__54950\,
            I => \N__54944\
        );

    \I__11656\ : LocalMux
    port map (
            O => \N__54947\,
            I => \N__54940\
        );

    \I__11655\ : InMux
    port map (
            O => \N__54944\,
            I => \N__54937\
        );

    \I__11654\ : InMux
    port map (
            O => \N__54943\,
            I => \N__54933\
        );

    \I__11653\ : Span4Mux_h
    port map (
            O => \N__54940\,
            I => \N__54930\
        );

    \I__11652\ : LocalMux
    port map (
            O => \N__54937\,
            I => \N__54927\
        );

    \I__11651\ : InMux
    port map (
            O => \N__54936\,
            I => \N__54924\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__54933\,
            I => \N__54921\
        );

    \I__11649\ : Span4Mux_v
    port map (
            O => \N__54930\,
            I => \N__54918\
        );

    \I__11648\ : Odrv4
    port map (
            O => \N__54927\,
            I => \c0.data_in_frame_3_1\
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__54924\,
            I => \c0.data_in_frame_3_1\
        );

    \I__11646\ : Odrv12
    port map (
            O => \N__54921\,
            I => \c0.data_in_frame_3_1\
        );

    \I__11645\ : Odrv4
    port map (
            O => \N__54918\,
            I => \c0.data_in_frame_3_1\
        );

    \I__11644\ : InMux
    port map (
            O => \N__54909\,
            I => \N__54906\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__54906\,
            I => \c0.n7_adj_4300\
        );

    \I__11642\ : SRMux
    port map (
            O => \N__54903\,
            I => \N__54900\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__54900\,
            I => \N__54897\
        );

    \I__11640\ : Odrv4
    port map (
            O => \N__54897\,
            I => \c0.n3_adj_4436\
        );

    \I__11639\ : SRMux
    port map (
            O => \N__54894\,
            I => \N__54891\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__54891\,
            I => \N__54888\
        );

    \I__11637\ : Odrv4
    port map (
            O => \N__54888\,
            I => \c0.n3_adj_4376\
        );

    \I__11636\ : InMux
    port map (
            O => \N__54885\,
            I => \N__54872\
        );

    \I__11635\ : InMux
    port map (
            O => \N__54884\,
            I => \N__54872\
        );

    \I__11634\ : InMux
    port map (
            O => \N__54883\,
            I => \N__54872\
        );

    \I__11633\ : InMux
    port map (
            O => \N__54882\,
            I => \N__54863\
        );

    \I__11632\ : InMux
    port map (
            O => \N__54881\,
            I => \N__54863\
        );

    \I__11631\ : InMux
    port map (
            O => \N__54880\,
            I => \N__54863\
        );

    \I__11630\ : InMux
    port map (
            O => \N__54879\,
            I => \N__54863\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__54872\,
            I => \N__54822\
        );

    \I__11628\ : LocalMux
    port map (
            O => \N__54863\,
            I => \N__54822\
        );

    \I__11627\ : InMux
    port map (
            O => \N__54862\,
            I => \N__54815\
        );

    \I__11626\ : InMux
    port map (
            O => \N__54861\,
            I => \N__54815\
        );

    \I__11625\ : InMux
    port map (
            O => \N__54860\,
            I => \N__54815\
        );

    \I__11624\ : InMux
    port map (
            O => \N__54859\,
            I => \N__54806\
        );

    \I__11623\ : InMux
    port map (
            O => \N__54858\,
            I => \N__54806\
        );

    \I__11622\ : InMux
    port map (
            O => \N__54857\,
            I => \N__54806\
        );

    \I__11621\ : InMux
    port map (
            O => \N__54856\,
            I => \N__54806\
        );

    \I__11620\ : InMux
    port map (
            O => \N__54855\,
            I => \N__54799\
        );

    \I__11619\ : InMux
    port map (
            O => \N__54854\,
            I => \N__54799\
        );

    \I__11618\ : InMux
    port map (
            O => \N__54853\,
            I => \N__54799\
        );

    \I__11617\ : InMux
    port map (
            O => \N__54852\,
            I => \N__54790\
        );

    \I__11616\ : InMux
    port map (
            O => \N__54851\,
            I => \N__54790\
        );

    \I__11615\ : InMux
    port map (
            O => \N__54850\,
            I => \N__54790\
        );

    \I__11614\ : InMux
    port map (
            O => \N__54849\,
            I => \N__54790\
        );

    \I__11613\ : InMux
    port map (
            O => \N__54848\,
            I => \N__54783\
        );

    \I__11612\ : InMux
    port map (
            O => \N__54847\,
            I => \N__54783\
        );

    \I__11611\ : InMux
    port map (
            O => \N__54846\,
            I => \N__54783\
        );

    \I__11610\ : InMux
    port map (
            O => \N__54845\,
            I => \N__54774\
        );

    \I__11609\ : InMux
    port map (
            O => \N__54844\,
            I => \N__54774\
        );

    \I__11608\ : InMux
    port map (
            O => \N__54843\,
            I => \N__54774\
        );

    \I__11607\ : InMux
    port map (
            O => \N__54842\,
            I => \N__54774\
        );

    \I__11606\ : InMux
    port map (
            O => \N__54841\,
            I => \N__54767\
        );

    \I__11605\ : InMux
    port map (
            O => \N__54840\,
            I => \N__54767\
        );

    \I__11604\ : InMux
    port map (
            O => \N__54839\,
            I => \N__54767\
        );

    \I__11603\ : InMux
    port map (
            O => \N__54838\,
            I => \N__54758\
        );

    \I__11602\ : InMux
    port map (
            O => \N__54837\,
            I => \N__54758\
        );

    \I__11601\ : InMux
    port map (
            O => \N__54836\,
            I => \N__54758\
        );

    \I__11600\ : InMux
    port map (
            O => \N__54835\,
            I => \N__54758\
        );

    \I__11599\ : CascadeMux
    port map (
            O => \N__54834\,
            I => \N__54755\
        );

    \I__11598\ : CascadeMux
    port map (
            O => \N__54833\,
            I => \N__54751\
        );

    \I__11597\ : CascadeMux
    port map (
            O => \N__54832\,
            I => \N__54747\
        );

    \I__11596\ : CascadeMux
    port map (
            O => \N__54831\,
            I => \N__54743\
        );

    \I__11595\ : CascadeMux
    port map (
            O => \N__54830\,
            I => \N__54733\
        );

    \I__11594\ : CascadeMux
    port map (
            O => \N__54829\,
            I => \N__54729\
        );

    \I__11593\ : CascadeMux
    port map (
            O => \N__54828\,
            I => \N__54725\
        );

    \I__11592\ : CascadeMux
    port map (
            O => \N__54827\,
            I => \N__54721\
        );

    \I__11591\ : Span4Mux_s3_v
    port map (
            O => \N__54822\,
            I => \N__54695\
        );

    \I__11590\ : LocalMux
    port map (
            O => \N__54815\,
            I => \N__54695\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__54806\,
            I => \N__54695\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__54799\,
            I => \N__54695\
        );

    \I__11587\ : LocalMux
    port map (
            O => \N__54790\,
            I => \N__54695\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__54783\,
            I => \N__54695\
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__54774\,
            I => \N__54695\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__54767\,
            I => \N__54695\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__54758\,
            I => \N__54695\
        );

    \I__11582\ : InMux
    port map (
            O => \N__54755\,
            I => \N__54680\
        );

    \I__11581\ : InMux
    port map (
            O => \N__54754\,
            I => \N__54680\
        );

    \I__11580\ : InMux
    port map (
            O => \N__54751\,
            I => \N__54680\
        );

    \I__11579\ : InMux
    port map (
            O => \N__54750\,
            I => \N__54680\
        );

    \I__11578\ : InMux
    port map (
            O => \N__54747\,
            I => \N__54680\
        );

    \I__11577\ : InMux
    port map (
            O => \N__54746\,
            I => \N__54680\
        );

    \I__11576\ : InMux
    port map (
            O => \N__54743\,
            I => \N__54680\
        );

    \I__11575\ : InMux
    port map (
            O => \N__54742\,
            I => \N__54673\
        );

    \I__11574\ : InMux
    port map (
            O => \N__54741\,
            I => \N__54673\
        );

    \I__11573\ : InMux
    port map (
            O => \N__54740\,
            I => \N__54673\
        );

    \I__11572\ : InMux
    port map (
            O => \N__54739\,
            I => \N__54664\
        );

    \I__11571\ : InMux
    port map (
            O => \N__54738\,
            I => \N__54664\
        );

    \I__11570\ : InMux
    port map (
            O => \N__54737\,
            I => \N__54664\
        );

    \I__11569\ : InMux
    port map (
            O => \N__54736\,
            I => \N__54664\
        );

    \I__11568\ : InMux
    port map (
            O => \N__54733\,
            I => \N__54649\
        );

    \I__11567\ : InMux
    port map (
            O => \N__54732\,
            I => \N__54649\
        );

    \I__11566\ : InMux
    port map (
            O => \N__54729\,
            I => \N__54649\
        );

    \I__11565\ : InMux
    port map (
            O => \N__54728\,
            I => \N__54649\
        );

    \I__11564\ : InMux
    port map (
            O => \N__54725\,
            I => \N__54649\
        );

    \I__11563\ : InMux
    port map (
            O => \N__54724\,
            I => \N__54649\
        );

    \I__11562\ : InMux
    port map (
            O => \N__54721\,
            I => \N__54649\
        );

    \I__11561\ : InMux
    port map (
            O => \N__54720\,
            I => \N__54642\
        );

    \I__11560\ : InMux
    port map (
            O => \N__54719\,
            I => \N__54642\
        );

    \I__11559\ : InMux
    port map (
            O => \N__54718\,
            I => \N__54642\
        );

    \I__11558\ : InMux
    port map (
            O => \N__54717\,
            I => \N__54633\
        );

    \I__11557\ : InMux
    port map (
            O => \N__54716\,
            I => \N__54633\
        );

    \I__11556\ : InMux
    port map (
            O => \N__54715\,
            I => \N__54633\
        );

    \I__11555\ : InMux
    port map (
            O => \N__54714\,
            I => \N__54633\
        );

    \I__11554\ : Span4Mux_v
    port map (
            O => \N__54695\,
            I => \N__54615\
        );

    \I__11553\ : LocalMux
    port map (
            O => \N__54680\,
            I => \N__54615\
        );

    \I__11552\ : LocalMux
    port map (
            O => \N__54673\,
            I => \N__54615\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__54664\,
            I => \N__54615\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__54649\,
            I => \N__54615\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__54642\,
            I => \N__54615\
        );

    \I__11548\ : LocalMux
    port map (
            O => \N__54633\,
            I => \N__54615\
        );

    \I__11547\ : CascadeMux
    port map (
            O => \N__54632\,
            I => \N__54590\
        );

    \I__11546\ : CascadeMux
    port map (
            O => \N__54631\,
            I => \N__54586\
        );

    \I__11545\ : CascadeMux
    port map (
            O => \N__54630\,
            I => \N__54582\
        );

    \I__11544\ : Span4Mux_v
    port map (
            O => \N__54615\,
            I => \N__54566\
        );

    \I__11543\ : InMux
    port map (
            O => \N__54614\,
            I => \N__54559\
        );

    \I__11542\ : InMux
    port map (
            O => \N__54613\,
            I => \N__54559\
        );

    \I__11541\ : InMux
    port map (
            O => \N__54612\,
            I => \N__54559\
        );

    \I__11540\ : InMux
    port map (
            O => \N__54611\,
            I => \N__54550\
        );

    \I__11539\ : InMux
    port map (
            O => \N__54610\,
            I => \N__54550\
        );

    \I__11538\ : InMux
    port map (
            O => \N__54609\,
            I => \N__54550\
        );

    \I__11537\ : InMux
    port map (
            O => \N__54608\,
            I => \N__54550\
        );

    \I__11536\ : InMux
    port map (
            O => \N__54607\,
            I => \N__54543\
        );

    \I__11535\ : InMux
    port map (
            O => \N__54606\,
            I => \N__54543\
        );

    \I__11534\ : InMux
    port map (
            O => \N__54605\,
            I => \N__54543\
        );

    \I__11533\ : InMux
    port map (
            O => \N__54604\,
            I => \N__54534\
        );

    \I__11532\ : InMux
    port map (
            O => \N__54603\,
            I => \N__54534\
        );

    \I__11531\ : InMux
    port map (
            O => \N__54602\,
            I => \N__54534\
        );

    \I__11530\ : InMux
    port map (
            O => \N__54601\,
            I => \N__54534\
        );

    \I__11529\ : InMux
    port map (
            O => \N__54600\,
            I => \N__54527\
        );

    \I__11528\ : InMux
    port map (
            O => \N__54599\,
            I => \N__54527\
        );

    \I__11527\ : InMux
    port map (
            O => \N__54598\,
            I => \N__54527\
        );

    \I__11526\ : InMux
    port map (
            O => \N__54597\,
            I => \N__54518\
        );

    \I__11525\ : InMux
    port map (
            O => \N__54596\,
            I => \N__54518\
        );

    \I__11524\ : InMux
    port map (
            O => \N__54595\,
            I => \N__54518\
        );

    \I__11523\ : InMux
    port map (
            O => \N__54594\,
            I => \N__54518\
        );

    \I__11522\ : InMux
    port map (
            O => \N__54593\,
            I => \N__54475\
        );

    \I__11521\ : InMux
    port map (
            O => \N__54590\,
            I => \N__54475\
        );

    \I__11520\ : InMux
    port map (
            O => \N__54589\,
            I => \N__54475\
        );

    \I__11519\ : InMux
    port map (
            O => \N__54586\,
            I => \N__54475\
        );

    \I__11518\ : InMux
    port map (
            O => \N__54585\,
            I => \N__54475\
        );

    \I__11517\ : InMux
    port map (
            O => \N__54582\,
            I => \N__54475\
        );

    \I__11516\ : InMux
    port map (
            O => \N__54581\,
            I => \N__54475\
        );

    \I__11515\ : CascadeMux
    port map (
            O => \N__54580\,
            I => \N__54471\
        );

    \I__11514\ : CascadeMux
    port map (
            O => \N__54579\,
            I => \N__54467\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__54578\,
            I => \N__54463\
        );

    \I__11512\ : CascadeMux
    port map (
            O => \N__54577\,
            I => \N__54458\
        );

    \I__11511\ : CascadeMux
    port map (
            O => \N__54576\,
            I => \N__54454\
        );

    \I__11510\ : CascadeMux
    port map (
            O => \N__54575\,
            I => \N__54450\
        );

    \I__11509\ : CascadeMux
    port map (
            O => \N__54574\,
            I => \N__54445\
        );

    \I__11508\ : CascadeMux
    port map (
            O => \N__54573\,
            I => \N__54441\
        );

    \I__11507\ : CascadeMux
    port map (
            O => \N__54572\,
            I => \N__54437\
        );

    \I__11506\ : CascadeMux
    port map (
            O => \N__54571\,
            I => \N__54432\
        );

    \I__11505\ : CascadeMux
    port map (
            O => \N__54570\,
            I => \N__54428\
        );

    \I__11504\ : CascadeMux
    port map (
            O => \N__54569\,
            I => \N__54424\
        );

    \I__11503\ : Span4Mux_h
    port map (
            O => \N__54566\,
            I => \N__54402\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__54559\,
            I => \N__54402\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__54550\,
            I => \N__54402\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__54543\,
            I => \N__54402\
        );

    \I__11499\ : LocalMux
    port map (
            O => \N__54534\,
            I => \N__54402\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__54527\,
            I => \N__54402\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__54518\,
            I => \N__54402\
        );

    \I__11496\ : InMux
    port map (
            O => \N__54517\,
            I => \N__54395\
        );

    \I__11495\ : InMux
    port map (
            O => \N__54516\,
            I => \N__54395\
        );

    \I__11494\ : InMux
    port map (
            O => \N__54515\,
            I => \N__54395\
        );

    \I__11493\ : InMux
    port map (
            O => \N__54514\,
            I => \N__54386\
        );

    \I__11492\ : InMux
    port map (
            O => \N__54513\,
            I => \N__54386\
        );

    \I__11491\ : InMux
    port map (
            O => \N__54512\,
            I => \N__54386\
        );

    \I__11490\ : InMux
    port map (
            O => \N__54511\,
            I => \N__54386\
        );

    \I__11489\ : InMux
    port map (
            O => \N__54510\,
            I => \N__54379\
        );

    \I__11488\ : InMux
    port map (
            O => \N__54509\,
            I => \N__54379\
        );

    \I__11487\ : InMux
    port map (
            O => \N__54508\,
            I => \N__54379\
        );

    \I__11486\ : InMux
    port map (
            O => \N__54507\,
            I => \N__54370\
        );

    \I__11485\ : InMux
    port map (
            O => \N__54506\,
            I => \N__54370\
        );

    \I__11484\ : InMux
    port map (
            O => \N__54505\,
            I => \N__54370\
        );

    \I__11483\ : InMux
    port map (
            O => \N__54504\,
            I => \N__54370\
        );

    \I__11482\ : InMux
    port map (
            O => \N__54503\,
            I => \N__54363\
        );

    \I__11481\ : InMux
    port map (
            O => \N__54502\,
            I => \N__54363\
        );

    \I__11480\ : InMux
    port map (
            O => \N__54501\,
            I => \N__54363\
        );

    \I__11479\ : InMux
    port map (
            O => \N__54500\,
            I => \N__54354\
        );

    \I__11478\ : InMux
    port map (
            O => \N__54499\,
            I => \N__54354\
        );

    \I__11477\ : InMux
    port map (
            O => \N__54498\,
            I => \N__54354\
        );

    \I__11476\ : InMux
    port map (
            O => \N__54497\,
            I => \N__54354\
        );

    \I__11475\ : InMux
    port map (
            O => \N__54496\,
            I => \N__54347\
        );

    \I__11474\ : InMux
    port map (
            O => \N__54495\,
            I => \N__54347\
        );

    \I__11473\ : InMux
    port map (
            O => \N__54494\,
            I => \N__54347\
        );

    \I__11472\ : InMux
    port map (
            O => \N__54493\,
            I => \N__54338\
        );

    \I__11471\ : InMux
    port map (
            O => \N__54492\,
            I => \N__54338\
        );

    \I__11470\ : InMux
    port map (
            O => \N__54491\,
            I => \N__54338\
        );

    \I__11469\ : InMux
    port map (
            O => \N__54490\,
            I => \N__54338\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__54475\,
            I => \N__54304\
        );

    \I__11467\ : InMux
    port map (
            O => \N__54474\,
            I => \N__54289\
        );

    \I__11466\ : InMux
    port map (
            O => \N__54471\,
            I => \N__54289\
        );

    \I__11465\ : InMux
    port map (
            O => \N__54470\,
            I => \N__54289\
        );

    \I__11464\ : InMux
    port map (
            O => \N__54467\,
            I => \N__54289\
        );

    \I__11463\ : InMux
    port map (
            O => \N__54466\,
            I => \N__54289\
        );

    \I__11462\ : InMux
    port map (
            O => \N__54463\,
            I => \N__54289\
        );

    \I__11461\ : InMux
    port map (
            O => \N__54462\,
            I => \N__54289\
        );

    \I__11460\ : InMux
    port map (
            O => \N__54461\,
            I => \N__54274\
        );

    \I__11459\ : InMux
    port map (
            O => \N__54458\,
            I => \N__54274\
        );

    \I__11458\ : InMux
    port map (
            O => \N__54457\,
            I => \N__54274\
        );

    \I__11457\ : InMux
    port map (
            O => \N__54454\,
            I => \N__54274\
        );

    \I__11456\ : InMux
    port map (
            O => \N__54453\,
            I => \N__54274\
        );

    \I__11455\ : InMux
    port map (
            O => \N__54450\,
            I => \N__54274\
        );

    \I__11454\ : InMux
    port map (
            O => \N__54449\,
            I => \N__54274\
        );

    \I__11453\ : InMux
    port map (
            O => \N__54448\,
            I => \N__54259\
        );

    \I__11452\ : InMux
    port map (
            O => \N__54445\,
            I => \N__54259\
        );

    \I__11451\ : InMux
    port map (
            O => \N__54444\,
            I => \N__54259\
        );

    \I__11450\ : InMux
    port map (
            O => \N__54441\,
            I => \N__54259\
        );

    \I__11449\ : InMux
    port map (
            O => \N__54440\,
            I => \N__54259\
        );

    \I__11448\ : InMux
    port map (
            O => \N__54437\,
            I => \N__54259\
        );

    \I__11447\ : InMux
    port map (
            O => \N__54436\,
            I => \N__54259\
        );

    \I__11446\ : InMux
    port map (
            O => \N__54435\,
            I => \N__54244\
        );

    \I__11445\ : InMux
    port map (
            O => \N__54432\,
            I => \N__54244\
        );

    \I__11444\ : InMux
    port map (
            O => \N__54431\,
            I => \N__54244\
        );

    \I__11443\ : InMux
    port map (
            O => \N__54428\,
            I => \N__54244\
        );

    \I__11442\ : InMux
    port map (
            O => \N__54427\,
            I => \N__54244\
        );

    \I__11441\ : InMux
    port map (
            O => \N__54424\,
            I => \N__54244\
        );

    \I__11440\ : InMux
    port map (
            O => \N__54423\,
            I => \N__54244\
        );

    \I__11439\ : CascadeMux
    port map (
            O => \N__54422\,
            I => \N__54240\
        );

    \I__11438\ : CascadeMux
    port map (
            O => \N__54421\,
            I => \N__54236\
        );

    \I__11437\ : CascadeMux
    port map (
            O => \N__54420\,
            I => \N__54232\
        );

    \I__11436\ : CascadeMux
    port map (
            O => \N__54419\,
            I => \N__54227\
        );

    \I__11435\ : CascadeMux
    port map (
            O => \N__54418\,
            I => \N__54223\
        );

    \I__11434\ : CascadeMux
    port map (
            O => \N__54417\,
            I => \N__54219\
        );

    \I__11433\ : Span4Mux_v
    port map (
            O => \N__54402\,
            I => \N__54199\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__54395\,
            I => \N__54199\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__54386\,
            I => \N__54199\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__54379\,
            I => \N__54199\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__54370\,
            I => \N__54199\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__54363\,
            I => \N__54199\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__54354\,
            I => \N__54199\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__54347\,
            I => \N__54199\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__54338\,
            I => \N__54199\
        );

    \I__11424\ : InMux
    port map (
            O => \N__54337\,
            I => \N__54192\
        );

    \I__11423\ : InMux
    port map (
            O => \N__54336\,
            I => \N__54192\
        );

    \I__11422\ : InMux
    port map (
            O => \N__54335\,
            I => \N__54192\
        );

    \I__11421\ : InMux
    port map (
            O => \N__54334\,
            I => \N__54183\
        );

    \I__11420\ : InMux
    port map (
            O => \N__54333\,
            I => \N__54183\
        );

    \I__11419\ : InMux
    port map (
            O => \N__54332\,
            I => \N__54183\
        );

    \I__11418\ : InMux
    port map (
            O => \N__54331\,
            I => \N__54183\
        );

    \I__11417\ : InMux
    port map (
            O => \N__54330\,
            I => \N__54176\
        );

    \I__11416\ : InMux
    port map (
            O => \N__54329\,
            I => \N__54176\
        );

    \I__11415\ : InMux
    port map (
            O => \N__54328\,
            I => \N__54176\
        );

    \I__11414\ : InMux
    port map (
            O => \N__54327\,
            I => \N__54167\
        );

    \I__11413\ : InMux
    port map (
            O => \N__54326\,
            I => \N__54167\
        );

    \I__11412\ : InMux
    port map (
            O => \N__54325\,
            I => \N__54167\
        );

    \I__11411\ : InMux
    port map (
            O => \N__54324\,
            I => \N__54167\
        );

    \I__11410\ : InMux
    port map (
            O => \N__54323\,
            I => \N__54160\
        );

    \I__11409\ : InMux
    port map (
            O => \N__54322\,
            I => \N__54160\
        );

    \I__11408\ : InMux
    port map (
            O => \N__54321\,
            I => \N__54160\
        );

    \I__11407\ : InMux
    port map (
            O => \N__54320\,
            I => \N__54151\
        );

    \I__11406\ : InMux
    port map (
            O => \N__54319\,
            I => \N__54151\
        );

    \I__11405\ : InMux
    port map (
            O => \N__54318\,
            I => \N__54151\
        );

    \I__11404\ : InMux
    port map (
            O => \N__54317\,
            I => \N__54151\
        );

    \I__11403\ : CascadeMux
    port map (
            O => \N__54316\,
            I => \N__54147\
        );

    \I__11402\ : CascadeMux
    port map (
            O => \N__54315\,
            I => \N__54143\
        );

    \I__11401\ : CascadeMux
    port map (
            O => \N__54314\,
            I => \N__54139\
        );

    \I__11400\ : InMux
    port map (
            O => \N__54313\,
            I => \N__54124\
        );

    \I__11399\ : InMux
    port map (
            O => \N__54312\,
            I => \N__54124\
        );

    \I__11398\ : InMux
    port map (
            O => \N__54311\,
            I => \N__54124\
        );

    \I__11397\ : InMux
    port map (
            O => \N__54310\,
            I => \N__54115\
        );

    \I__11396\ : InMux
    port map (
            O => \N__54309\,
            I => \N__54115\
        );

    \I__11395\ : InMux
    port map (
            O => \N__54308\,
            I => \N__54115\
        );

    \I__11394\ : InMux
    port map (
            O => \N__54307\,
            I => \N__54115\
        );

    \I__11393\ : Span4Mux_s0_v
    port map (
            O => \N__54304\,
            I => \N__54106\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__54289\,
            I => \N__54106\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__54274\,
            I => \N__54106\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__54259\,
            I => \N__54106\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__54244\,
            I => \N__54103\
        );

    \I__11388\ : InMux
    port map (
            O => \N__54243\,
            I => \N__54088\
        );

    \I__11387\ : InMux
    port map (
            O => \N__54240\,
            I => \N__54088\
        );

    \I__11386\ : InMux
    port map (
            O => \N__54239\,
            I => \N__54088\
        );

    \I__11385\ : InMux
    port map (
            O => \N__54236\,
            I => \N__54088\
        );

    \I__11384\ : InMux
    port map (
            O => \N__54235\,
            I => \N__54088\
        );

    \I__11383\ : InMux
    port map (
            O => \N__54232\,
            I => \N__54088\
        );

    \I__11382\ : InMux
    port map (
            O => \N__54231\,
            I => \N__54088\
        );

    \I__11381\ : InMux
    port map (
            O => \N__54230\,
            I => \N__54073\
        );

    \I__11380\ : InMux
    port map (
            O => \N__54227\,
            I => \N__54073\
        );

    \I__11379\ : InMux
    port map (
            O => \N__54226\,
            I => \N__54073\
        );

    \I__11378\ : InMux
    port map (
            O => \N__54223\,
            I => \N__54073\
        );

    \I__11377\ : InMux
    port map (
            O => \N__54222\,
            I => \N__54073\
        );

    \I__11376\ : InMux
    port map (
            O => \N__54219\,
            I => \N__54073\
        );

    \I__11375\ : InMux
    port map (
            O => \N__54218\,
            I => \N__54073\
        );

    \I__11374\ : Span4Mux_v
    port map (
            O => \N__54199\,
            I => \N__54058\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__54192\,
            I => \N__54058\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__54183\,
            I => \N__54058\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__54176\,
            I => \N__54058\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__54167\,
            I => \N__54058\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__54160\,
            I => \N__54058\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__54151\,
            I => \N__54058\
        );

    \I__11367\ : InMux
    port map (
            O => \N__54150\,
            I => \N__54043\
        );

    \I__11366\ : InMux
    port map (
            O => \N__54147\,
            I => \N__54043\
        );

    \I__11365\ : InMux
    port map (
            O => \N__54146\,
            I => \N__54043\
        );

    \I__11364\ : InMux
    port map (
            O => \N__54143\,
            I => \N__54043\
        );

    \I__11363\ : InMux
    port map (
            O => \N__54142\,
            I => \N__54043\
        );

    \I__11362\ : InMux
    port map (
            O => \N__54139\,
            I => \N__54043\
        );

    \I__11361\ : InMux
    port map (
            O => \N__54138\,
            I => \N__54043\
        );

    \I__11360\ : InMux
    port map (
            O => \N__54137\,
            I => \N__54036\
        );

    \I__11359\ : InMux
    port map (
            O => \N__54136\,
            I => \N__54036\
        );

    \I__11358\ : InMux
    port map (
            O => \N__54135\,
            I => \N__54036\
        );

    \I__11357\ : InMux
    port map (
            O => \N__54134\,
            I => \N__54027\
        );

    \I__11356\ : InMux
    port map (
            O => \N__54133\,
            I => \N__54027\
        );

    \I__11355\ : InMux
    port map (
            O => \N__54132\,
            I => \N__54027\
        );

    \I__11354\ : InMux
    port map (
            O => \N__54131\,
            I => \N__54027\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__54124\,
            I => \N__54015\
        );

    \I__11352\ : LocalMux
    port map (
            O => \N__54115\,
            I => \N__54015\
        );

    \I__11351\ : Span4Mux_v
    port map (
            O => \N__54106\,
            I => \N__54002\
        );

    \I__11350\ : Span4Mux_h
    port map (
            O => \N__54103\,
            I => \N__54002\
        );

    \I__11349\ : LocalMux
    port map (
            O => \N__54088\,
            I => \N__54002\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__54073\,
            I => \N__54002\
        );

    \I__11347\ : Span4Mux_v
    port map (
            O => \N__54058\,
            I => \N__54002\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__54043\,
            I => \N__54002\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__54036\,
            I => \N__53990\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__54027\,
            I => \N__53990\
        );

    \I__11343\ : InMux
    port map (
            O => \N__54026\,
            I => \N__53983\
        );

    \I__11342\ : InMux
    port map (
            O => \N__54025\,
            I => \N__53983\
        );

    \I__11341\ : InMux
    port map (
            O => \N__54024\,
            I => \N__53983\
        );

    \I__11340\ : InMux
    port map (
            O => \N__54023\,
            I => \N__53974\
        );

    \I__11339\ : InMux
    port map (
            O => \N__54022\,
            I => \N__53974\
        );

    \I__11338\ : InMux
    port map (
            O => \N__54021\,
            I => \N__53974\
        );

    \I__11337\ : InMux
    port map (
            O => \N__54020\,
            I => \N__53974\
        );

    \I__11336\ : Span4Mux_h
    port map (
            O => \N__54015\,
            I => \N__53971\
        );

    \I__11335\ : Span4Mux_v
    port map (
            O => \N__54002\,
            I => \N__53968\
        );

    \I__11334\ : InMux
    port map (
            O => \N__54001\,
            I => \N__53961\
        );

    \I__11333\ : InMux
    port map (
            O => \N__54000\,
            I => \N__53961\
        );

    \I__11332\ : InMux
    port map (
            O => \N__53999\,
            I => \N__53961\
        );

    \I__11331\ : InMux
    port map (
            O => \N__53998\,
            I => \N__53952\
        );

    \I__11330\ : InMux
    port map (
            O => \N__53997\,
            I => \N__53952\
        );

    \I__11329\ : InMux
    port map (
            O => \N__53996\,
            I => \N__53952\
        );

    \I__11328\ : InMux
    port map (
            O => \N__53995\,
            I => \N__53952\
        );

    \I__11327\ : Span12Mux_h
    port map (
            O => \N__53990\,
            I => \N__53949\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__53983\,
            I => \N__53944\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__53974\,
            I => \N__53944\
        );

    \I__11324\ : Sp12to4
    port map (
            O => \N__53971\,
            I => \N__53941\
        );

    \I__11323\ : Sp12to4
    port map (
            O => \N__53968\,
            I => \N__53934\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__53961\,
            I => \N__53934\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__53952\,
            I => \N__53934\
        );

    \I__11320\ : Span12Mux_v
    port map (
            O => \N__53949\,
            I => \N__53929\
        );

    \I__11319\ : Span12Mux_h
    port map (
            O => \N__53944\,
            I => \N__53929\
        );

    \I__11318\ : Span12Mux_s8_v
    port map (
            O => \N__53941\,
            I => \N__53924\
        );

    \I__11317\ : Span12Mux_h
    port map (
            O => \N__53934\,
            I => \N__53924\
        );

    \I__11316\ : Odrv12
    port map (
            O => \N__53929\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11315\ : Odrv12
    port map (
            O => \N__53924\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11314\ : InMux
    port map (
            O => \N__53919\,
            I => \bfn_19_32_0_\
        );

    \I__11313\ : CascadeMux
    port map (
            O => \N__53916\,
            I => \N__53912\
        );

    \I__11312\ : InMux
    port map (
            O => \N__53915\,
            I => \N__53905\
        );

    \I__11311\ : InMux
    port map (
            O => \N__53912\,
            I => \N__53902\
        );

    \I__11310\ : InMux
    port map (
            O => \N__53911\,
            I => \N__53895\
        );

    \I__11309\ : InMux
    port map (
            O => \N__53910\,
            I => \N__53895\
        );

    \I__11308\ : InMux
    port map (
            O => \N__53909\,
            I => \N__53895\
        );

    \I__11307\ : InMux
    port map (
            O => \N__53908\,
            I => \N__53891\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__53905\,
            I => \N__53888\
        );

    \I__11305\ : LocalMux
    port map (
            O => \N__53902\,
            I => \N__53885\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__53895\,
            I => \N__53882\
        );

    \I__11303\ : InMux
    port map (
            O => \N__53894\,
            I => \N__53878\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__53891\,
            I => \N__53874\
        );

    \I__11301\ : Span4Mux_v
    port map (
            O => \N__53888\,
            I => \N__53871\
        );

    \I__11300\ : Span4Mux_h
    port map (
            O => \N__53885\,
            I => \N__53866\
        );

    \I__11299\ : Span4Mux_v
    port map (
            O => \N__53882\,
            I => \N__53866\
        );

    \I__11298\ : InMux
    port map (
            O => \N__53881\,
            I => \N__53863\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__53878\,
            I => \N__53860\
        );

    \I__11296\ : InMux
    port map (
            O => \N__53877\,
            I => \N__53857\
        );

    \I__11295\ : Span4Mux_v
    port map (
            O => \N__53874\,
            I => \N__53854\
        );

    \I__11294\ : Span4Mux_v
    port map (
            O => \N__53871\,
            I => \N__53851\
        );

    \I__11293\ : Span4Mux_v
    port map (
            O => \N__53866\,
            I => \N__53848\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__53863\,
            I => \N__53843\
        );

    \I__11291\ : Span12Mux_v
    port map (
            O => \N__53860\,
            I => \N__53843\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__53857\,
            I => \N__53838\
        );

    \I__11289\ : Span4Mux_v
    port map (
            O => \N__53854\,
            I => \N__53838\
        );

    \I__11288\ : Span4Mux_h
    port map (
            O => \N__53851\,
            I => \N__53835\
        );

    \I__11287\ : Span4Mux_h
    port map (
            O => \N__53848\,
            I => \N__53832\
        );

    \I__11286\ : Odrv12
    port map (
            O => \N__53843\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__11285\ : Odrv4
    port map (
            O => \N__53838\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__11284\ : Odrv4
    port map (
            O => \N__53835\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__11283\ : Odrv4
    port map (
            O => \N__53832\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__11282\ : SRMux
    port map (
            O => \N__53823\,
            I => \N__53820\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__53820\,
            I => \N__53817\
        );

    \I__11280\ : Odrv12
    port map (
            O => \N__53817\,
            I => \c0.n3_adj_4373\
        );

    \I__11279\ : InMux
    port map (
            O => \N__53814\,
            I => \N__53811\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__53811\,
            I => \N__53808\
        );

    \I__11277\ : Span4Mux_h
    port map (
            O => \N__53808\,
            I => \N__53804\
        );

    \I__11276\ : InMux
    port map (
            O => \N__53807\,
            I => \N__53799\
        );

    \I__11275\ : Span4Mux_v
    port map (
            O => \N__53804\,
            I => \N__53796\
        );

    \I__11274\ : InMux
    port map (
            O => \N__53803\,
            I => \N__53793\
        );

    \I__11273\ : InMux
    port map (
            O => \N__53802\,
            I => \N__53790\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__53799\,
            I => \N__53787\
        );

    \I__11271\ : Span4Mux_v
    port map (
            O => \N__53796\,
            I => \N__53782\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__53793\,
            I => \N__53782\
        );

    \I__11269\ : LocalMux
    port map (
            O => \N__53790\,
            I => \N__53779\
        );

    \I__11268\ : Span4Mux_h
    port map (
            O => \N__53787\,
            I => \N__53776\
        );

    \I__11267\ : Odrv4
    port map (
            O => \N__53782\,
            I => \c0.n17856\
        );

    \I__11266\ : Odrv4
    port map (
            O => \N__53779\,
            I => \c0.n17856\
        );

    \I__11265\ : Odrv4
    port map (
            O => \N__53776\,
            I => \c0.n17856\
        );

    \I__11264\ : InMux
    port map (
            O => \N__53769\,
            I => \N__53761\
        );

    \I__11263\ : InMux
    port map (
            O => \N__53768\,
            I => \N__53756\
        );

    \I__11262\ : InMux
    port map (
            O => \N__53767\,
            I => \N__53753\
        );

    \I__11261\ : InMux
    port map (
            O => \N__53766\,
            I => \N__53750\
        );

    \I__11260\ : InMux
    port map (
            O => \N__53765\,
            I => \N__53737\
        );

    \I__11259\ : InMux
    port map (
            O => \N__53764\,
            I => \N__53734\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__53761\,
            I => \N__53731\
        );

    \I__11257\ : InMux
    port map (
            O => \N__53760\,
            I => \N__53728\
        );

    \I__11256\ : InMux
    port map (
            O => \N__53759\,
            I => \N__53725\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__53756\,
            I => \N__53717\
        );

    \I__11254\ : LocalMux
    port map (
            O => \N__53753\,
            I => \N__53717\
        );

    \I__11253\ : LocalMux
    port map (
            O => \N__53750\,
            I => \N__53717\
        );

    \I__11252\ : InMux
    port map (
            O => \N__53749\,
            I => \N__53714\
        );

    \I__11251\ : InMux
    port map (
            O => \N__53748\,
            I => \N__53709\
        );

    \I__11250\ : InMux
    port map (
            O => \N__53747\,
            I => \N__53706\
        );

    \I__11249\ : InMux
    port map (
            O => \N__53746\,
            I => \N__53703\
        );

    \I__11248\ : InMux
    port map (
            O => \N__53745\,
            I => \N__53700\
        );

    \I__11247\ : InMux
    port map (
            O => \N__53744\,
            I => \N__53689\
        );

    \I__11246\ : InMux
    port map (
            O => \N__53743\,
            I => \N__53686\
        );

    \I__11245\ : InMux
    port map (
            O => \N__53742\,
            I => \N__53683\
        );

    \I__11244\ : InMux
    port map (
            O => \N__53741\,
            I => \N__53680\
        );

    \I__11243\ : InMux
    port map (
            O => \N__53740\,
            I => \N__53677\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__53737\,
            I => \N__53666\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__53734\,
            I => \N__53666\
        );

    \I__11240\ : Sp12to4
    port map (
            O => \N__53731\,
            I => \N__53666\
        );

    \I__11239\ : LocalMux
    port map (
            O => \N__53728\,
            I => \N__53666\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__53725\,
            I => \N__53666\
        );

    \I__11237\ : InMux
    port map (
            O => \N__53724\,
            I => \N__53662\
        );

    \I__11236\ : Span4Mux_v
    port map (
            O => \N__53717\,
            I => \N__53657\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__53714\,
            I => \N__53657\
        );

    \I__11234\ : InMux
    port map (
            O => \N__53713\,
            I => \N__53654\
        );

    \I__11233\ : InMux
    port map (
            O => \N__53712\,
            I => \N__53651\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__53709\,
            I => \N__53642\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__53706\,
            I => \N__53642\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__53703\,
            I => \N__53642\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__53700\,
            I => \N__53642\
        );

    \I__11228\ : InMux
    port map (
            O => \N__53699\,
            I => \N__53637\
        );

    \I__11227\ : InMux
    port map (
            O => \N__53698\,
            I => \N__53634\
        );

    \I__11226\ : InMux
    port map (
            O => \N__53697\,
            I => \N__53631\
        );

    \I__11225\ : InMux
    port map (
            O => \N__53696\,
            I => \N__53628\
        );

    \I__11224\ : InMux
    port map (
            O => \N__53695\,
            I => \N__53625\
        );

    \I__11223\ : InMux
    port map (
            O => \N__53694\,
            I => \N__53622\
        );

    \I__11222\ : InMux
    port map (
            O => \N__53693\,
            I => \N__53619\
        );

    \I__11221\ : InMux
    port map (
            O => \N__53692\,
            I => \N__53616\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__53689\,
            I => \N__53603\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__53686\,
            I => \N__53603\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__53683\,
            I => \N__53603\
        );

    \I__11217\ : LocalMux
    port map (
            O => \N__53680\,
            I => \N__53603\
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__53677\,
            I => \N__53603\
        );

    \I__11215\ : Span12Mux_s8_v
    port map (
            O => \N__53666\,
            I => \N__53603\
        );

    \I__11214\ : InMux
    port map (
            O => \N__53665\,
            I => \N__53600\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__53662\,
            I => \N__53589\
        );

    \I__11212\ : Sp12to4
    port map (
            O => \N__53657\,
            I => \N__53589\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__53654\,
            I => \N__53589\
        );

    \I__11210\ : LocalMux
    port map (
            O => \N__53651\,
            I => \N__53589\
        );

    \I__11209\ : Span12Mux_v
    port map (
            O => \N__53642\,
            I => \N__53589\
        );

    \I__11208\ : InMux
    port map (
            O => \N__53641\,
            I => \N__53586\
        );

    \I__11207\ : InMux
    port map (
            O => \N__53640\,
            I => \N__53583\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__53637\,
            I => \N__53580\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__53634\,
            I => \N__53563\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__53631\,
            I => \N__53563\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__53628\,
            I => \N__53563\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__53625\,
            I => \N__53563\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__53622\,
            I => \N__53563\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__53619\,
            I => \N__53563\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__53616\,
            I => \N__53563\
        );

    \I__11198\ : Span12Mux_v
    port map (
            O => \N__53603\,
            I => \N__53563\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__53600\,
            I => \N__53558\
        );

    \I__11196\ : Span12Mux_v
    port map (
            O => \N__53589\,
            I => \N__53558\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__53586\,
            I => \c0.n1306\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__53583\,
            I => \c0.n1306\
        );

    \I__11193\ : Odrv4
    port map (
            O => \N__53580\,
            I => \c0.n1306\
        );

    \I__11192\ : Odrv12
    port map (
            O => \N__53563\,
            I => \c0.n1306\
        );

    \I__11191\ : Odrv12
    port map (
            O => \N__53558\,
            I => \c0.n1306\
        );

    \I__11190\ : InMux
    port map (
            O => \N__53547\,
            I => \N__53544\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__53544\,
            I => \N__53539\
        );

    \I__11188\ : InMux
    port map (
            O => \N__53543\,
            I => \N__53536\
        );

    \I__11187\ : InMux
    port map (
            O => \N__53542\,
            I => \N__53533\
        );

    \I__11186\ : Span4Mux_h
    port map (
            O => \N__53539\,
            I => \N__53530\
        );

    \I__11185\ : LocalMux
    port map (
            O => \N__53536\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__53533\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__11183\ : Odrv4
    port map (
            O => \N__53530\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__11182\ : InMux
    port map (
            O => \N__53523\,
            I => \bfn_19_30_0_\
        );

    \I__11181\ : SRMux
    port map (
            O => \N__53520\,
            I => \N__53517\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__53517\,
            I => \c0.n3_adj_4378\
        );

    \I__11179\ : InMux
    port map (
            O => \N__53514\,
            I => \N__53511\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__53511\,
            I => \N__53506\
        );

    \I__11177\ : InMux
    port map (
            O => \N__53510\,
            I => \N__53503\
        );

    \I__11176\ : InMux
    port map (
            O => \N__53509\,
            I => \N__53500\
        );

    \I__11175\ : Span4Mux_v
    port map (
            O => \N__53506\,
            I => \N__53497\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__53503\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__53500\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__11172\ : Odrv4
    port map (
            O => \N__53497\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__11171\ : InMux
    port map (
            O => \N__53490\,
            I => \bfn_19_31_0_\
        );

    \I__11170\ : CascadeMux
    port map (
            O => \N__53487\,
            I => \N__53484\
        );

    \I__11169\ : InMux
    port map (
            O => \N__53484\,
            I => \N__53481\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__53481\,
            I => \N__53476\
        );

    \I__11167\ : InMux
    port map (
            O => \N__53480\,
            I => \N__53473\
        );

    \I__11166\ : InMux
    port map (
            O => \N__53479\,
            I => \N__53470\
        );

    \I__11165\ : Span4Mux_h
    port map (
            O => \N__53476\,
            I => \N__53467\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__53473\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__53470\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__11162\ : Odrv4
    port map (
            O => \N__53467\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__11161\ : InMux
    port map (
            O => \N__53460\,
            I => \bfn_19_29_0_\
        );

    \I__11160\ : SRMux
    port map (
            O => \N__53457\,
            I => \N__53454\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__53454\,
            I => \N__53451\
        );

    \I__11158\ : Odrv12
    port map (
            O => \N__53451\,
            I => \c0.n3_adj_4380\
        );

    \I__11157\ : InMux
    port map (
            O => \N__53448\,
            I => \N__53445\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__53445\,
            I => \N__53442\
        );

    \I__11155\ : Span4Mux_v
    port map (
            O => \N__53442\,
            I => \N__53437\
        );

    \I__11154\ : InMux
    port map (
            O => \N__53441\,
            I => \N__53434\
        );

    \I__11153\ : InMux
    port map (
            O => \N__53440\,
            I => \N__53431\
        );

    \I__11152\ : Span4Mux_h
    port map (
            O => \N__53437\,
            I => \N__53428\
        );

    \I__11151\ : LocalMux
    port map (
            O => \N__53434\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__53431\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__11149\ : Odrv4
    port map (
            O => \N__53428\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__11148\ : InMux
    port map (
            O => \N__53421\,
            I => \bfn_19_28_0_\
        );

    \I__11147\ : SRMux
    port map (
            O => \N__53418\,
            I => \N__53415\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__53415\,
            I => \N__53412\
        );

    \I__11145\ : Odrv4
    port map (
            O => \N__53412\,
            I => \c0.n3_adj_4382\
        );

    \I__11144\ : InMux
    port map (
            O => \N__53409\,
            I => \N__53405\
        );

    \I__11143\ : InMux
    port map (
            O => \N__53408\,
            I => \N__53401\
        );

    \I__11142\ : LocalMux
    port map (
            O => \N__53405\,
            I => \N__53398\
        );

    \I__11141\ : InMux
    port map (
            O => \N__53404\,
            I => \N__53395\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__53401\,
            I => \N__53390\
        );

    \I__11139\ : Span4Mux_v
    port map (
            O => \N__53398\,
            I => \N__53390\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__53395\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__11137\ : Odrv4
    port map (
            O => \N__53390\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__11136\ : InMux
    port map (
            O => \N__53385\,
            I => \bfn_19_27_0_\
        );

    \I__11135\ : SRMux
    port map (
            O => \N__53382\,
            I => \N__53379\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__53379\,
            I => \c0.n3_adj_4384\
        );

    \I__11133\ : InMux
    port map (
            O => \N__53376\,
            I => \N__53371\
        );

    \I__11132\ : InMux
    port map (
            O => \N__53375\,
            I => \N__53368\
        );

    \I__11131\ : InMux
    port map (
            O => \N__53374\,
            I => \N__53365\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__53371\,
            I => \N__53362\
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__53368\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__53365\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__11127\ : Odrv4
    port map (
            O => \N__53362\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__11126\ : InMux
    port map (
            O => \N__53355\,
            I => \bfn_19_26_0_\
        );

    \I__11125\ : SRMux
    port map (
            O => \N__53352\,
            I => \N__53349\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__53349\,
            I => \c0.n3_adj_4386\
        );

    \I__11123\ : InMux
    port map (
            O => \N__53346\,
            I => \N__53343\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__53343\,
            I => \N__53338\
        );

    \I__11121\ : InMux
    port map (
            O => \N__53342\,
            I => \N__53335\
        );

    \I__11120\ : InMux
    port map (
            O => \N__53341\,
            I => \N__53332\
        );

    \I__11119\ : Odrv4
    port map (
            O => \N__53338\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__11118\ : LocalMux
    port map (
            O => \N__53335\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__53332\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__11116\ : InMux
    port map (
            O => \N__53325\,
            I => \bfn_19_25_0_\
        );

    \I__11115\ : SRMux
    port map (
            O => \N__53322\,
            I => \N__53319\
        );

    \I__11114\ : LocalMux
    port map (
            O => \N__53319\,
            I => \N__53316\
        );

    \I__11113\ : Odrv12
    port map (
            O => \N__53316\,
            I => \c0.n3_adj_4388\
        );

    \I__11112\ : CascadeMux
    port map (
            O => \N__53313\,
            I => \N__53310\
        );

    \I__11111\ : InMux
    port map (
            O => \N__53310\,
            I => \N__53306\
        );

    \I__11110\ : InMux
    port map (
            O => \N__53309\,
            I => \N__53303\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__53306\,
            I => \N__53299\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__53303\,
            I => \N__53296\
        );

    \I__11107\ : InMux
    port map (
            O => \N__53302\,
            I => \N__53293\
        );

    \I__11106\ : Span4Mux_h
    port map (
            O => \N__53299\,
            I => \N__53290\
        );

    \I__11105\ : Odrv4
    port map (
            O => \N__53296\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__53293\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__11103\ : Odrv4
    port map (
            O => \N__53290\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__11102\ : InMux
    port map (
            O => \N__53283\,
            I => \bfn_19_24_0_\
        );

    \I__11101\ : SRMux
    port map (
            O => \N__53280\,
            I => \N__53277\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__53277\,
            I => \N__53274\
        );

    \I__11099\ : Odrv12
    port map (
            O => \N__53274\,
            I => \c0.n3_adj_4390\
        );

    \I__11098\ : InMux
    port map (
            O => \N__53271\,
            I => \N__53267\
        );

    \I__11097\ : InMux
    port map (
            O => \N__53270\,
            I => \N__53264\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__53267\,
            I => \N__53258\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__53264\,
            I => \N__53258\
        );

    \I__11094\ : InMux
    port map (
            O => \N__53263\,
            I => \N__53255\
        );

    \I__11093\ : Span4Mux_v
    port map (
            O => \N__53258\,
            I => \N__53252\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__53255\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__11091\ : Odrv4
    port map (
            O => \N__53252\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__11090\ : InMux
    port map (
            O => \N__53247\,
            I => \bfn_19_23_0_\
        );

    \I__11089\ : SRMux
    port map (
            O => \N__53244\,
            I => \N__53241\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__53241\,
            I => \N__53238\
        );

    \I__11087\ : Span4Mux_h
    port map (
            O => \N__53238\,
            I => \N__53235\
        );

    \I__11086\ : Odrv4
    port map (
            O => \N__53235\,
            I => \c0.n3_adj_4392\
        );

    \I__11085\ : SRMux
    port map (
            O => \N__53232\,
            I => \N__53229\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__53229\,
            I => \N__53226\
        );

    \I__11083\ : Span4Mux_v
    port map (
            O => \N__53226\,
            I => \N__53223\
        );

    \I__11082\ : Odrv4
    port map (
            O => \N__53223\,
            I => \c0.n3_adj_4396\
        );

    \I__11081\ : InMux
    port map (
            O => \N__53220\,
            I => \N__53216\
        );

    \I__11080\ : InMux
    port map (
            O => \N__53219\,
            I => \N__53213\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__53216\,
            I => \N__53207\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__53213\,
            I => \N__53207\
        );

    \I__11077\ : InMux
    port map (
            O => \N__53212\,
            I => \N__53204\
        );

    \I__11076\ : Span4Mux_v
    port map (
            O => \N__53207\,
            I => \N__53201\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__53204\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__11074\ : Odrv4
    port map (
            O => \N__53201\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__11073\ : InMux
    port map (
            O => \N__53196\,
            I => \bfn_19_22_0_\
        );

    \I__11072\ : SRMux
    port map (
            O => \N__53193\,
            I => \N__53190\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__53190\,
            I => \N__53187\
        );

    \I__11070\ : Span4Mux_h
    port map (
            O => \N__53187\,
            I => \N__53184\
        );

    \I__11069\ : Odrv4
    port map (
            O => \N__53184\,
            I => \c0.n3_adj_4394\
        );

    \I__11068\ : CascadeMux
    port map (
            O => \N__53181\,
            I => \N__53177\
        );

    \I__11067\ : InMux
    port map (
            O => \N__53180\,
            I => \N__53174\
        );

    \I__11066\ : InMux
    port map (
            O => \N__53177\,
            I => \N__53171\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__53174\,
            I => \N__53165\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__53171\,
            I => \N__53165\
        );

    \I__11063\ : InMux
    port map (
            O => \N__53170\,
            I => \N__53162\
        );

    \I__11062\ : Span4Mux_v
    port map (
            O => \N__53165\,
            I => \N__53159\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__53162\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__11060\ : Odrv4
    port map (
            O => \N__53159\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__11059\ : InMux
    port map (
            O => \N__53154\,
            I => \bfn_19_20_0_\
        );

    \I__11058\ : SRMux
    port map (
            O => \N__53151\,
            I => \N__53148\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__53148\,
            I => \N__53145\
        );

    \I__11056\ : Span4Mux_v
    port map (
            O => \N__53145\,
            I => \N__53142\
        );

    \I__11055\ : Span4Mux_h
    port map (
            O => \N__53142\,
            I => \N__53139\
        );

    \I__11054\ : Odrv4
    port map (
            O => \N__53139\,
            I => \c0.n3_adj_4398\
        );

    \I__11053\ : InMux
    port map (
            O => \N__53136\,
            I => \N__53133\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__53133\,
            I => \N__53129\
        );

    \I__11051\ : InMux
    port map (
            O => \N__53132\,
            I => \N__53126\
        );

    \I__11050\ : Span4Mux_v
    port map (
            O => \N__53129\,
            I => \N__53120\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__53126\,
            I => \N__53120\
        );

    \I__11048\ : InMux
    port map (
            O => \N__53125\,
            I => \N__53117\
        );

    \I__11047\ : Sp12to4
    port map (
            O => \N__53120\,
            I => \N__53114\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__53117\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__11045\ : Odrv12
    port map (
            O => \N__53114\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__11044\ : InMux
    port map (
            O => \N__53109\,
            I => \bfn_19_21_0_\
        );

    \I__11043\ : InMux
    port map (
            O => \N__53106\,
            I => \bfn_19_19_0_\
        );

    \I__11042\ : CascadeMux
    port map (
            O => \N__53103\,
            I => \N__53100\
        );

    \I__11041\ : InMux
    port map (
            O => \N__53100\,
            I => \N__53096\
        );

    \I__11040\ : InMux
    port map (
            O => \N__53099\,
            I => \N__53093\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__53096\,
            I => \N__53090\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__53093\,
            I => \N__53084\
        );

    \I__11037\ : Span4Mux_v
    port map (
            O => \N__53090\,
            I => \N__53084\
        );

    \I__11036\ : InMux
    port map (
            O => \N__53089\,
            I => \N__53081\
        );

    \I__11035\ : Span4Mux_v
    port map (
            O => \N__53084\,
            I => \N__53078\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__53081\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__11033\ : Odrv4
    port map (
            O => \N__53078\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__11032\ : InMux
    port map (
            O => \N__53073\,
            I => \bfn_19_18_0_\
        );

    \I__11031\ : SRMux
    port map (
            O => \N__53070\,
            I => \N__53067\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__53067\,
            I => \N__53064\
        );

    \I__11029\ : Span4Mux_v
    port map (
            O => \N__53064\,
            I => \N__53061\
        );

    \I__11028\ : Odrv4
    port map (
            O => \N__53061\,
            I => \c0.n3_adj_4402\
        );

    \I__11027\ : CascadeMux
    port map (
            O => \N__53058\,
            I => \N__53055\
        );

    \I__11026\ : InMux
    port map (
            O => \N__53055\,
            I => \N__53051\
        );

    \I__11025\ : InMux
    port map (
            O => \N__53054\,
            I => \N__53048\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__53051\,
            I => \N__53045\
        );

    \I__11023\ : LocalMux
    port map (
            O => \N__53048\,
            I => \N__53042\
        );

    \I__11022\ : Span4Mux_h
    port map (
            O => \N__53045\,
            I => \N__53039\
        );

    \I__11021\ : Span4Mux_h
    port map (
            O => \N__53042\,
            I => \N__53033\
        );

    \I__11020\ : Span4Mux_v
    port map (
            O => \N__53039\,
            I => \N__53033\
        );

    \I__11019\ : InMux
    port map (
            O => \N__53038\,
            I => \N__53030\
        );

    \I__11018\ : Span4Mux_v
    port map (
            O => \N__53033\,
            I => \N__53027\
        );

    \I__11017\ : LocalMux
    port map (
            O => \N__53030\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__11016\ : Odrv4
    port map (
            O => \N__53027\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__11015\ : InMux
    port map (
            O => \N__53022\,
            I => \bfn_19_17_0_\
        );

    \I__11014\ : SRMux
    port map (
            O => \N__53019\,
            I => \N__53016\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__53016\,
            I => \N__53013\
        );

    \I__11012\ : Span4Mux_h
    port map (
            O => \N__53013\,
            I => \N__53010\
        );

    \I__11011\ : Odrv4
    port map (
            O => \N__53010\,
            I => \c0.n3_adj_4404\
        );

    \I__11010\ : InMux
    port map (
            O => \N__53007\,
            I => \N__53003\
        );

    \I__11009\ : InMux
    port map (
            O => \N__53006\,
            I => \N__53000\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__53003\,
            I => \N__52997\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__53000\,
            I => \N__52993\
        );

    \I__11006\ : Span4Mux_v
    port map (
            O => \N__52997\,
            I => \N__52990\
        );

    \I__11005\ : InMux
    port map (
            O => \N__52996\,
            I => \N__52987\
        );

    \I__11004\ : Span12Mux_h
    port map (
            O => \N__52993\,
            I => \N__52982\
        );

    \I__11003\ : Sp12to4
    port map (
            O => \N__52990\,
            I => \N__52982\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__52987\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__11001\ : Odrv12
    port map (
            O => \N__52982\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__11000\ : InMux
    port map (
            O => \N__52977\,
            I => \bfn_19_16_0_\
        );

    \I__10999\ : SRMux
    port map (
            O => \N__52974\,
            I => \N__52971\
        );

    \I__10998\ : LocalMux
    port map (
            O => \N__52971\,
            I => \N__52968\
        );

    \I__10997\ : Span4Mux_h
    port map (
            O => \N__52968\,
            I => \N__52965\
        );

    \I__10996\ : Span4Mux_v
    port map (
            O => \N__52965\,
            I => \N__52962\
        );

    \I__10995\ : Odrv4
    port map (
            O => \N__52962\,
            I => \c0.n3_adj_4406\
        );

    \I__10994\ : CascadeMux
    port map (
            O => \N__52959\,
            I => \N__52956\
        );

    \I__10993\ : InMux
    port map (
            O => \N__52956\,
            I => \N__52952\
        );

    \I__10992\ : InMux
    port map (
            O => \N__52955\,
            I => \N__52949\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__52952\,
            I => \N__52946\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__52949\,
            I => \N__52943\
        );

    \I__10989\ : Sp12to4
    port map (
            O => \N__52946\,
            I => \N__52939\
        );

    \I__10988\ : Span4Mux_v
    port map (
            O => \N__52943\,
            I => \N__52936\
        );

    \I__10987\ : InMux
    port map (
            O => \N__52942\,
            I => \N__52933\
        );

    \I__10986\ : Span12Mux_s9_v
    port map (
            O => \N__52939\,
            I => \N__52930\
        );

    \I__10985\ : Odrv4
    port map (
            O => \N__52936\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__52933\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__10983\ : Odrv12
    port map (
            O => \N__52930\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__10982\ : InMux
    port map (
            O => \N__52923\,
            I => \bfn_19_15_0_\
        );

    \I__10981\ : SRMux
    port map (
            O => \N__52920\,
            I => \N__52917\
        );

    \I__10980\ : LocalMux
    port map (
            O => \N__52917\,
            I => \N__52914\
        );

    \I__10979\ : Span4Mux_v
    port map (
            O => \N__52914\,
            I => \N__52911\
        );

    \I__10978\ : Odrv4
    port map (
            O => \N__52911\,
            I => \c0.n3_adj_4408\
        );

    \I__10977\ : InMux
    port map (
            O => \N__52908\,
            I => \bfn_19_14_0_\
        );

    \I__10976\ : InMux
    port map (
            O => \N__52905\,
            I => \N__52901\
        );

    \I__10975\ : InMux
    port map (
            O => \N__52904\,
            I => \N__52898\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__52901\,
            I => \N__52895\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__52898\,
            I => \N__52892\
        );

    \I__10972\ : Sp12to4
    port map (
            O => \N__52895\,
            I => \N__52886\
        );

    \I__10971\ : Sp12to4
    port map (
            O => \N__52892\,
            I => \N__52886\
        );

    \I__10970\ : InMux
    port map (
            O => \N__52891\,
            I => \N__52883\
        );

    \I__10969\ : Span12Mux_s11_v
    port map (
            O => \N__52886\,
            I => \N__52880\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__52883\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__10967\ : Odrv12
    port map (
            O => \N__52880\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__10966\ : InMux
    port map (
            O => \N__52875\,
            I => \bfn_19_13_0_\
        );

    \I__10965\ : SRMux
    port map (
            O => \N__52872\,
            I => \N__52869\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__52869\,
            I => \N__52866\
        );

    \I__10963\ : Span4Mux_v
    port map (
            O => \N__52866\,
            I => \N__52863\
        );

    \I__10962\ : Span4Mux_v
    port map (
            O => \N__52863\,
            I => \N__52860\
        );

    \I__10961\ : Span4Mux_v
    port map (
            O => \N__52860\,
            I => \N__52857\
        );

    \I__10960\ : Odrv4
    port map (
            O => \N__52857\,
            I => \c0.n3_adj_4412\
        );

    \I__10959\ : SRMux
    port map (
            O => \N__52854\,
            I => \N__52851\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__52851\,
            I => \N__52848\
        );

    \I__10957\ : Span4Mux_v
    port map (
            O => \N__52848\,
            I => \N__52845\
        );

    \I__10956\ : Span4Mux_v
    port map (
            O => \N__52845\,
            I => \N__52842\
        );

    \I__10955\ : Span4Mux_v
    port map (
            O => \N__52842\,
            I => \N__52839\
        );

    \I__10954\ : Odrv4
    port map (
            O => \N__52839\,
            I => \c0.n3_adj_4416\
        );

    \I__10953\ : InMux
    port map (
            O => \N__52836\,
            I => \N__52832\
        );

    \I__10952\ : InMux
    port map (
            O => \N__52835\,
            I => \N__52829\
        );

    \I__10951\ : LocalMux
    port map (
            O => \N__52832\,
            I => \N__52826\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__52829\,
            I => \N__52823\
        );

    \I__10949\ : Span4Mux_h
    port map (
            O => \N__52826\,
            I => \N__52820\
        );

    \I__10948\ : Span4Mux_h
    port map (
            O => \N__52823\,
            I => \N__52817\
        );

    \I__10947\ : Sp12to4
    port map (
            O => \N__52820\,
            I => \N__52811\
        );

    \I__10946\ : Sp12to4
    port map (
            O => \N__52817\,
            I => \N__52811\
        );

    \I__10945\ : InMux
    port map (
            O => \N__52816\,
            I => \N__52808\
        );

    \I__10944\ : Span12Mux_v
    port map (
            O => \N__52811\,
            I => \N__52805\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__52808\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__10942\ : Odrv12
    port map (
            O => \N__52805\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__10941\ : InMux
    port map (
            O => \N__52800\,
            I => \bfn_19_12_0_\
        );

    \I__10940\ : SRMux
    port map (
            O => \N__52797\,
            I => \N__52794\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__52794\,
            I => \N__52791\
        );

    \I__10938\ : Span4Mux_h
    port map (
            O => \N__52791\,
            I => \N__52788\
        );

    \I__10937\ : Span4Mux_v
    port map (
            O => \N__52788\,
            I => \N__52785\
        );

    \I__10936\ : Span4Mux_v
    port map (
            O => \N__52785\,
            I => \N__52782\
        );

    \I__10935\ : Span4Mux_h
    port map (
            O => \N__52782\,
            I => \N__52779\
        );

    \I__10934\ : Odrv4
    port map (
            O => \N__52779\,
            I => \c0.n3_adj_4414\
        );

    \I__10933\ : InMux
    port map (
            O => \N__52776\,
            I => \N__52773\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__52773\,
            I => \N__52770\
        );

    \I__10931\ : Span4Mux_h
    port map (
            O => \N__52770\,
            I => \N__52766\
        );

    \I__10930\ : InMux
    port map (
            O => \N__52769\,
            I => \N__52763\
        );

    \I__10929\ : Span4Mux_v
    port map (
            O => \N__52766\,
            I => \N__52760\
        );

    \I__10928\ : LocalMux
    port map (
            O => \N__52763\,
            I => \N__52757\
        );

    \I__10927\ : Sp12to4
    port map (
            O => \N__52760\,
            I => \N__52751\
        );

    \I__10926\ : Span12Mux_h
    port map (
            O => \N__52757\,
            I => \N__52751\
        );

    \I__10925\ : InMux
    port map (
            O => \N__52756\,
            I => \N__52748\
        );

    \I__10924\ : Span12Mux_v
    port map (
            O => \N__52751\,
            I => \N__52745\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__52748\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__10922\ : Odrv12
    port map (
            O => \N__52745\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__10921\ : InMux
    port map (
            O => \N__52740\,
            I => \bfn_19_10_0_\
        );

    \I__10920\ : SRMux
    port map (
            O => \N__52737\,
            I => \N__52734\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__52734\,
            I => \N__52731\
        );

    \I__10918\ : Span4Mux_v
    port map (
            O => \N__52731\,
            I => \N__52728\
        );

    \I__10917\ : Span4Mux_v
    port map (
            O => \N__52728\,
            I => \N__52725\
        );

    \I__10916\ : Odrv4
    port map (
            O => \N__52725\,
            I => \c0.n3_adj_4418\
        );

    \I__10915\ : InMux
    port map (
            O => \N__52722\,
            I => \N__52716\
        );

    \I__10914\ : InMux
    port map (
            O => \N__52721\,
            I => \N__52716\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__52716\,
            I => \N__52713\
        );

    \I__10912\ : Sp12to4
    port map (
            O => \N__52713\,
            I => \N__52709\
        );

    \I__10911\ : InMux
    port map (
            O => \N__52712\,
            I => \N__52706\
        );

    \I__10910\ : Span12Mux_v
    port map (
            O => \N__52709\,
            I => \N__52703\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__52706\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__10908\ : Odrv12
    port map (
            O => \N__52703\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__10907\ : InMux
    port map (
            O => \N__52698\,
            I => \bfn_19_11_0_\
        );

    \I__10906\ : InMux
    port map (
            O => \N__52695\,
            I => \N__52691\
        );

    \I__10905\ : InMux
    port map (
            O => \N__52694\,
            I => \N__52688\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__52691\,
            I => \N__52685\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__52688\,
            I => \N__52682\
        );

    \I__10902\ : Span4Mux_v
    port map (
            O => \N__52685\,
            I => \N__52679\
        );

    \I__10901\ : Span4Mux_v
    port map (
            O => \N__52682\,
            I => \N__52676\
        );

    \I__10900\ : Span4Mux_h
    port map (
            O => \N__52679\,
            I => \N__52673\
        );

    \I__10899\ : Span4Mux_v
    port map (
            O => \N__52676\,
            I => \N__52670\
        );

    \I__10898\ : Span4Mux_v
    port map (
            O => \N__52673\,
            I => \N__52666\
        );

    \I__10897\ : Sp12to4
    port map (
            O => \N__52670\,
            I => \N__52663\
        );

    \I__10896\ : InMux
    port map (
            O => \N__52669\,
            I => \N__52660\
        );

    \I__10895\ : Odrv4
    port map (
            O => \N__52666\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__10894\ : Odrv12
    port map (
            O => \N__52663\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__52660\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__10892\ : InMux
    port map (
            O => \N__52653\,
            I => \bfn_19_9_0_\
        );

    \I__10891\ : SRMux
    port map (
            O => \N__52650\,
            I => \N__52647\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__52647\,
            I => \N__52644\
        );

    \I__10889\ : Span4Mux_h
    port map (
            O => \N__52644\,
            I => \N__52641\
        );

    \I__10888\ : Span4Mux_h
    port map (
            O => \N__52641\,
            I => \N__52638\
        );

    \I__10887\ : Span4Mux_v
    port map (
            O => \N__52638\,
            I => \N__52635\
        );

    \I__10886\ : Odrv4
    port map (
            O => \N__52635\,
            I => \c0.n3_adj_4420\
        );

    \I__10885\ : InMux
    port map (
            O => \N__52632\,
            I => \N__52629\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__52629\,
            I => \N__52625\
        );

    \I__10883\ : InMux
    port map (
            O => \N__52628\,
            I => \N__52622\
        );

    \I__10882\ : Span4Mux_h
    port map (
            O => \N__52625\,
            I => \N__52619\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__52622\,
            I => \N__52616\
        );

    \I__10880\ : Sp12to4
    port map (
            O => \N__52619\,
            I => \N__52610\
        );

    \I__10879\ : Sp12to4
    port map (
            O => \N__52616\,
            I => \N__52610\
        );

    \I__10878\ : InMux
    port map (
            O => \N__52615\,
            I => \N__52607\
        );

    \I__10877\ : Span12Mux_v
    port map (
            O => \N__52610\,
            I => \N__52604\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__52607\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__10875\ : Odrv12
    port map (
            O => \N__52604\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__10874\ : InMux
    port map (
            O => \N__52599\,
            I => \bfn_19_8_0_\
        );

    \I__10873\ : SRMux
    port map (
            O => \N__52596\,
            I => \N__52593\
        );

    \I__10872\ : LocalMux
    port map (
            O => \N__52593\,
            I => \N__52590\
        );

    \I__10871\ : Span4Mux_v
    port map (
            O => \N__52590\,
            I => \N__52587\
        );

    \I__10870\ : Span4Mux_v
    port map (
            O => \N__52587\,
            I => \N__52584\
        );

    \I__10869\ : Span4Mux_v
    port map (
            O => \N__52584\,
            I => \N__52581\
        );

    \I__10868\ : Span4Mux_h
    port map (
            O => \N__52581\,
            I => \N__52578\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__52578\,
            I => \c0.n3_adj_4422\
        );

    \I__10866\ : InMux
    port map (
            O => \N__52575\,
            I => \N__52572\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__52572\,
            I => \N__52569\
        );

    \I__10864\ : Span4Mux_v
    port map (
            O => \N__52569\,
            I => \N__52565\
        );

    \I__10863\ : InMux
    port map (
            O => \N__52568\,
            I => \N__52562\
        );

    \I__10862\ : Span4Mux_v
    port map (
            O => \N__52565\,
            I => \N__52556\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__52562\,
            I => \N__52556\
        );

    \I__10860\ : InMux
    port map (
            O => \N__52561\,
            I => \N__52553\
        );

    \I__10859\ : Span4Mux_v
    port map (
            O => \N__52556\,
            I => \N__52549\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__52553\,
            I => \N__52546\
        );

    \I__10857\ : InMux
    port map (
            O => \N__52552\,
            I => \N__52543\
        );

    \I__10856\ : Span4Mux_v
    port map (
            O => \N__52549\,
            I => \N__52540\
        );

    \I__10855\ : Span4Mux_h
    port map (
            O => \N__52546\,
            I => \N__52537\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__52543\,
            I => \N__52534\
        );

    \I__10853\ : Span4Mux_v
    port map (
            O => \N__52540\,
            I => \N__52531\
        );

    \I__10852\ : Sp12to4
    port map (
            O => \N__52537\,
            I => \N__52526\
        );

    \I__10851\ : Sp12to4
    port map (
            O => \N__52534\,
            I => \N__52526\
        );

    \I__10850\ : Span4Mux_h
    port map (
            O => \N__52531\,
            I => \N__52522\
        );

    \I__10849\ : Span12Mux_v
    port map (
            O => \N__52526\,
            I => \N__52519\
        );

    \I__10848\ : InMux
    port map (
            O => \N__52525\,
            I => \N__52516\
        );

    \I__10847\ : Odrv4
    port map (
            O => \N__52522\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__10846\ : Odrv12
    port map (
            O => \N__52519\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__52516\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__10844\ : InMux
    port map (
            O => \N__52509\,
            I => \bfn_19_7_0_\
        );

    \I__10843\ : SRMux
    port map (
            O => \N__52506\,
            I => \N__52503\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__52503\,
            I => \N__52500\
        );

    \I__10841\ : Span4Mux_v
    port map (
            O => \N__52500\,
            I => \N__52497\
        );

    \I__10840\ : Span4Mux_v
    port map (
            O => \N__52497\,
            I => \N__52494\
        );

    \I__10839\ : Sp12to4
    port map (
            O => \N__52494\,
            I => \N__52491\
        );

    \I__10838\ : Span12Mux_h
    port map (
            O => \N__52491\,
            I => \N__52488\
        );

    \I__10837\ : Odrv12
    port map (
            O => \N__52488\,
            I => \c0.n3_adj_4424\
        );

    \I__10836\ : InMux
    port map (
            O => \N__52485\,
            I => \N__52482\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__52482\,
            I => \N__52477\
        );

    \I__10834\ : InMux
    port map (
            O => \N__52481\,
            I => \N__52474\
        );

    \I__10833\ : InMux
    port map (
            O => \N__52480\,
            I => \N__52471\
        );

    \I__10832\ : Span4Mux_v
    port map (
            O => \N__52477\,
            I => \N__52468\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__52474\,
            I => \N__52465\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__52471\,
            I => \N__52462\
        );

    \I__10829\ : Sp12to4
    port map (
            O => \N__52468\,
            I => \N__52459\
        );

    \I__10828\ : Span4Mux_h
    port map (
            O => \N__52465\,
            I => \N__52456\
        );

    \I__10827\ : Span12Mux_h
    port map (
            O => \N__52462\,
            I => \N__52451\
        );

    \I__10826\ : Span12Mux_h
    port map (
            O => \N__52459\,
            I => \N__52446\
        );

    \I__10825\ : Sp12to4
    port map (
            O => \N__52456\,
            I => \N__52446\
        );

    \I__10824\ : InMux
    port map (
            O => \N__52455\,
            I => \N__52443\
        );

    \I__10823\ : InMux
    port map (
            O => \N__52454\,
            I => \N__52440\
        );

    \I__10822\ : Span12Mux_v
    port map (
            O => \N__52451\,
            I => \N__52437\
        );

    \I__10821\ : Span12Mux_v
    port map (
            O => \N__52446\,
            I => \N__52434\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__52443\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__52440\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__10818\ : Odrv12
    port map (
            O => \N__52437\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__10817\ : Odrv12
    port map (
            O => \N__52434\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__10816\ : InMux
    port map (
            O => \N__52425\,
            I => \bfn_19_6_0_\
        );

    \I__10815\ : SRMux
    port map (
            O => \N__52422\,
            I => \N__52419\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__52419\,
            I => \N__52416\
        );

    \I__10813\ : Span4Mux_v
    port map (
            O => \N__52416\,
            I => \N__52413\
        );

    \I__10812\ : Odrv4
    port map (
            O => \N__52413\,
            I => \c0.n3_adj_4426\
        );

    \I__10811\ : InMux
    port map (
            O => \N__52410\,
            I => \N__52404\
        );

    \I__10810\ : InMux
    port map (
            O => \N__52409\,
            I => \N__52401\
        );

    \I__10809\ : InMux
    port map (
            O => \N__52408\,
            I => \N__52398\
        );

    \I__10808\ : InMux
    port map (
            O => \N__52407\,
            I => \N__52395\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__52404\,
            I => \N__52392\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__52401\,
            I => \N__52389\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__52398\,
            I => \N__52384\
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__52395\,
            I => \N__52384\
        );

    \I__10803\ : Span4Mux_h
    port map (
            O => \N__52392\,
            I => \N__52381\
        );

    \I__10802\ : Span4Mux_h
    port map (
            O => \N__52389\,
            I => \N__52378\
        );

    \I__10801\ : Span4Mux_h
    port map (
            O => \N__52384\,
            I => \N__52375\
        );

    \I__10800\ : Span4Mux_v
    port map (
            O => \N__52381\,
            I => \N__52371\
        );

    \I__10799\ : Sp12to4
    port map (
            O => \N__52378\,
            I => \N__52366\
        );

    \I__10798\ : Sp12to4
    port map (
            O => \N__52375\,
            I => \N__52366\
        );

    \I__10797\ : InMux
    port map (
            O => \N__52374\,
            I => \N__52363\
        );

    \I__10796\ : Span4Mux_v
    port map (
            O => \N__52371\,
            I => \N__52359\
        );

    \I__10795\ : Span12Mux_s7_v
    port map (
            O => \N__52366\,
            I => \N__52356\
        );

    \I__10794\ : LocalMux
    port map (
            O => \N__52363\,
            I => \N__52353\
        );

    \I__10793\ : InMux
    port map (
            O => \N__52362\,
            I => \N__52350\
        );

    \I__10792\ : Span4Mux_v
    port map (
            O => \N__52359\,
            I => \N__52347\
        );

    \I__10791\ : Span12Mux_v
    port map (
            O => \N__52356\,
            I => \N__52344\
        );

    \I__10790\ : Odrv4
    port map (
            O => \N__52353\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__52350\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__10788\ : Odrv4
    port map (
            O => \N__52347\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__10787\ : Odrv12
    port map (
            O => \N__52344\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__10786\ : InMux
    port map (
            O => \N__52335\,
            I => \bfn_19_5_0_\
        );

    \I__10785\ : SRMux
    port map (
            O => \N__52332\,
            I => \N__52329\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__52329\,
            I => \N__52326\
        );

    \I__10783\ : Span4Mux_h
    port map (
            O => \N__52326\,
            I => \N__52323\
        );

    \I__10782\ : Odrv4
    port map (
            O => \N__52323\,
            I => \c0.n3_adj_4428\
        );

    \I__10781\ : InMux
    port map (
            O => \N__52320\,
            I => \bfn_19_4_0_\
        );

    \I__10780\ : SRMux
    port map (
            O => \N__52317\,
            I => \N__52314\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__52314\,
            I => \N__52311\
        );

    \I__10778\ : Span4Mux_h
    port map (
            O => \N__52311\,
            I => \N__52308\
        );

    \I__10777\ : Span4Mux_v
    port map (
            O => \N__52308\,
            I => \N__52305\
        );

    \I__10776\ : Odrv4
    port map (
            O => \N__52305\,
            I => \c0.n3_adj_4434\
        );

    \I__10775\ : InMux
    port map (
            O => \N__52302\,
            I => \bfn_19_3_0_\
        );

    \I__10774\ : SRMux
    port map (
            O => \N__52299\,
            I => \N__52296\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__52296\,
            I => \N__52293\
        );

    \I__10772\ : Span4Mux_v
    port map (
            O => \N__52293\,
            I => \N__52290\
        );

    \I__10771\ : Span4Mux_v
    port map (
            O => \N__52290\,
            I => \N__52287\
        );

    \I__10770\ : Odrv4
    port map (
            O => \N__52287\,
            I => \c0.n3_adj_4432\
        );

    \I__10769\ : CascadeMux
    port map (
            O => \N__52284\,
            I => \N__52281\
        );

    \I__10768\ : InMux
    port map (
            O => \N__52281\,
            I => \N__52278\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__52278\,
            I => \c0.n161\
        );

    \I__10766\ : InMux
    port map (
            O => \N__52275\,
            I => \bfn_19_2_0_\
        );

    \I__10765\ : InMux
    port map (
            O => \N__52272\,
            I => \N__52269\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__52269\,
            I => \c0.n41_adj_4292\
        );

    \I__10763\ : CascadeMux
    port map (
            O => \N__52266\,
            I => \c0.n42_adj_4272_cascade_\
        );

    \I__10762\ : InMux
    port map (
            O => \N__52263\,
            I => \N__52260\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__52260\,
            I => \c0.n44_adj_4270\
        );

    \I__10760\ : InMux
    port map (
            O => \N__52257\,
            I => \N__52254\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__52254\,
            I => \c0.n50_adj_4296\
        );

    \I__10758\ : InMux
    port map (
            O => \N__52251\,
            I => \N__52248\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__52248\,
            I => \c0.n43_adj_4275\
        );

    \I__10756\ : CascadeMux
    port map (
            O => \N__52245\,
            I => \N__52242\
        );

    \I__10755\ : InMux
    port map (
            O => \N__52242\,
            I => \N__52238\
        );

    \I__10754\ : CascadeMux
    port map (
            O => \N__52241\,
            I => \N__52235\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__52238\,
            I => \N__52232\
        );

    \I__10752\ : InMux
    port map (
            O => \N__52235\,
            I => \N__52229\
        );

    \I__10751\ : Span4Mux_v
    port map (
            O => \N__52232\,
            I => \N__52226\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__52229\,
            I => \N__52223\
        );

    \I__10749\ : Sp12to4
    port map (
            O => \N__52226\,
            I => \N__52220\
        );

    \I__10748\ : Odrv4
    port map (
            O => \N__52223\,
            I => \c0.data_in_frame_28_7\
        );

    \I__10747\ : Odrv12
    port map (
            O => \N__52220\,
            I => \c0.data_in_frame_28_7\
        );

    \I__10746\ : CascadeMux
    port map (
            O => \N__52215\,
            I => \N__52212\
        );

    \I__10745\ : InMux
    port map (
            O => \N__52212\,
            I => \N__52209\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__52209\,
            I => \c0.n45_adj_4298\
        );

    \I__10743\ : InMux
    port map (
            O => \N__52206\,
            I => \N__52201\
        );

    \I__10742\ : InMux
    port map (
            O => \N__52205\,
            I => \N__52198\
        );

    \I__10741\ : CascadeMux
    port map (
            O => \N__52204\,
            I => \N__52195\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__52201\,
            I => \N__52192\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__52198\,
            I => \N__52188\
        );

    \I__10738\ : InMux
    port map (
            O => \N__52195\,
            I => \N__52185\
        );

    \I__10737\ : Span4Mux_h
    port map (
            O => \N__52192\,
            I => \N__52182\
        );

    \I__10736\ : InMux
    port map (
            O => \N__52191\,
            I => \N__52179\
        );

    \I__10735\ : Span4Mux_v
    port map (
            O => \N__52188\,
            I => \N__52176\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__52185\,
            I => \c0.data_in_frame_25_3\
        );

    \I__10733\ : Odrv4
    port map (
            O => \N__52182\,
            I => \c0.data_in_frame_25_3\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__52179\,
            I => \c0.data_in_frame_25_3\
        );

    \I__10731\ : Odrv4
    port map (
            O => \N__52176\,
            I => \c0.data_in_frame_25_3\
        );

    \I__10730\ : InMux
    port map (
            O => \N__52167\,
            I => \N__52162\
        );

    \I__10729\ : InMux
    port map (
            O => \N__52166\,
            I => \N__52159\
        );

    \I__10728\ : CascadeMux
    port map (
            O => \N__52165\,
            I => \N__52156\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__52162\,
            I => \N__52150\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__52159\,
            I => \N__52150\
        );

    \I__10725\ : InMux
    port map (
            O => \N__52156\,
            I => \N__52145\
        );

    \I__10724\ : InMux
    port map (
            O => \N__52155\,
            I => \N__52145\
        );

    \I__10723\ : Odrv12
    port map (
            O => \N__52150\,
            I => \c0.data_in_frame_25_2\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__52145\,
            I => \c0.data_in_frame_25_2\
        );

    \I__10721\ : InMux
    port map (
            O => \N__52140\,
            I => \N__52137\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__52137\,
            I => \c0.n40_adj_4294\
        );

    \I__10719\ : InMux
    port map (
            O => \N__52134\,
            I => \N__52129\
        );

    \I__10718\ : InMux
    port map (
            O => \N__52133\,
            I => \N__52124\
        );

    \I__10717\ : InMux
    port map (
            O => \N__52132\,
            I => \N__52124\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__52129\,
            I => \N__52121\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__52124\,
            I => \N__52118\
        );

    \I__10714\ : Odrv4
    port map (
            O => \N__52121\,
            I => \c0.n5_adj_4349\
        );

    \I__10713\ : Odrv4
    port map (
            O => \N__52118\,
            I => \c0.n5_adj_4349\
        );

    \I__10712\ : CascadeMux
    port map (
            O => \N__52113\,
            I => \c0.n10_adj_4371_cascade_\
        );

    \I__10711\ : InMux
    port map (
            O => \N__52110\,
            I => \N__52107\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__52107\,
            I => \c0.n12_adj_4372\
        );

    \I__10709\ : CascadeMux
    port map (
            O => \N__52104\,
            I => \c0.n12_adj_4671_cascade_\
        );

    \I__10708\ : CascadeMux
    port map (
            O => \N__52101\,
            I => \N__52098\
        );

    \I__10707\ : InMux
    port map (
            O => \N__52098\,
            I => \N__52094\
        );

    \I__10706\ : CascadeMux
    port map (
            O => \N__52097\,
            I => \N__52091\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__52094\,
            I => \N__52087\
        );

    \I__10704\ : InMux
    port map (
            O => \N__52091\,
            I => \N__52084\
        );

    \I__10703\ : InMux
    port map (
            O => \N__52090\,
            I => \N__52081\
        );

    \I__10702\ : Span4Mux_v
    port map (
            O => \N__52087\,
            I => \N__52078\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__52084\,
            I => \N__52075\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__52081\,
            I => \N__52072\
        );

    \I__10699\ : Sp12to4
    port map (
            O => \N__52078\,
            I => \N__52068\
        );

    \I__10698\ : Span4Mux_h
    port map (
            O => \N__52075\,
            I => \N__52065\
        );

    \I__10697\ : Span4Mux_h
    port map (
            O => \N__52072\,
            I => \N__52062\
        );

    \I__10696\ : CascadeMux
    port map (
            O => \N__52071\,
            I => \N__52059\
        );

    \I__10695\ : Span12Mux_h
    port map (
            O => \N__52068\,
            I => \N__52056\
        );

    \I__10694\ : Sp12to4
    port map (
            O => \N__52065\,
            I => \N__52051\
        );

    \I__10693\ : Sp12to4
    port map (
            O => \N__52062\,
            I => \N__52051\
        );

    \I__10692\ : InMux
    port map (
            O => \N__52059\,
            I => \N__52048\
        );

    \I__10691\ : Span12Mux_v
    port map (
            O => \N__52056\,
            I => \N__52045\
        );

    \I__10690\ : Span12Mux_v
    port map (
            O => \N__52051\,
            I => \N__52042\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__52048\,
            I => \c0.data_in_frame_24_7\
        );

    \I__10688\ : Odrv12
    port map (
            O => \N__52045\,
            I => \c0.data_in_frame_24_7\
        );

    \I__10687\ : Odrv12
    port map (
            O => \N__52042\,
            I => \c0.data_in_frame_24_7\
        );

    \I__10686\ : InMux
    port map (
            O => \N__52035\,
            I => \N__52032\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__52032\,
            I => \c0.n25467\
        );

    \I__10684\ : InMux
    port map (
            O => \N__52029\,
            I => \N__52025\
        );

    \I__10683\ : InMux
    port map (
            O => \N__52028\,
            I => \N__52022\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__52025\,
            I => \c0.n24098\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__52022\,
            I => \c0.n24098\
        );

    \I__10680\ : CascadeMux
    port map (
            O => \N__52017\,
            I => \N__52014\
        );

    \I__10679\ : InMux
    port map (
            O => \N__52014\,
            I => \N__52010\
        );

    \I__10678\ : InMux
    port map (
            O => \N__52013\,
            I => \N__52007\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__52010\,
            I => \N__52004\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__52007\,
            I => \c0.data_in_frame_29_4\
        );

    \I__10675\ : Odrv12
    port map (
            O => \N__52004\,
            I => \c0.data_in_frame_29_4\
        );

    \I__10674\ : InMux
    port map (
            O => \N__51999\,
            I => \N__51995\
        );

    \I__10673\ : InMux
    port map (
            O => \N__51998\,
            I => \N__51992\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__51995\,
            I => \N__51987\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__51992\,
            I => \N__51987\
        );

    \I__10670\ : Odrv4
    port map (
            O => \N__51987\,
            I => \c0.n23533\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__51984\,
            I => \N__51981\
        );

    \I__10668\ : InMux
    port map (
            O => \N__51981\,
            I => \N__51978\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__51978\,
            I => \N__51975\
        );

    \I__10666\ : Span4Mux_v
    port map (
            O => \N__51975\,
            I => \N__51972\
        );

    \I__10665\ : Odrv4
    port map (
            O => \N__51972\,
            I => \c0.n5_adj_4370\
        );

    \I__10664\ : InMux
    port map (
            O => \N__51969\,
            I => \N__51966\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__51966\,
            I => \N__51963\
        );

    \I__10662\ : Odrv4
    port map (
            O => \N__51963\,
            I => \c0.n10_adj_4371\
        );

    \I__10661\ : CascadeMux
    port map (
            O => \N__51960\,
            I => \c0.n10_adj_4439_cascade_\
        );

    \I__10660\ : InMux
    port map (
            O => \N__51957\,
            I => \N__51954\
        );

    \I__10659\ : LocalMux
    port map (
            O => \N__51954\,
            I => \c0.n20_adj_4441\
        );

    \I__10658\ : CascadeMux
    port map (
            O => \N__51951\,
            I => \c0.n13_adj_4442_cascade_\
        );

    \I__10657\ : CascadeMux
    port map (
            O => \N__51948\,
            I => \c0.n24528_cascade_\
        );

    \I__10656\ : InMux
    port map (
            O => \N__51945\,
            I => \N__51940\
        );

    \I__10655\ : InMux
    port map (
            O => \N__51944\,
            I => \N__51937\
        );

    \I__10654\ : InMux
    port map (
            O => \N__51943\,
            I => \N__51934\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__51940\,
            I => \N__51931\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__51937\,
            I => \c0.n23718\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__51934\,
            I => \c0.n23718\
        );

    \I__10650\ : Odrv4
    port map (
            O => \N__51931\,
            I => \c0.n23718\
        );

    \I__10649\ : InMux
    port map (
            O => \N__51924\,
            I => \N__51921\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__51921\,
            I => \N__51918\
        );

    \I__10647\ : Odrv4
    port map (
            O => \N__51918\,
            I => \c0.n12_adj_4506\
        );

    \I__10646\ : InMux
    port map (
            O => \N__51915\,
            I => \N__51912\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__51912\,
            I => \c0.n20_adj_4512\
        );

    \I__10644\ : InMux
    port map (
            O => \N__51909\,
            I => \N__51906\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__51906\,
            I => \c0.n24_adj_4509\
        );

    \I__10642\ : InMux
    port map (
            O => \N__51903\,
            I => \N__51900\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__51900\,
            I => \c0.n22_adj_4507\
        );

    \I__10640\ : InMux
    port map (
            O => \N__51897\,
            I => \N__51894\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__51894\,
            I => \c0.n23627\
        );

    \I__10638\ : CascadeMux
    port map (
            O => \N__51891\,
            I => \c0.n23627_cascade_\
        );

    \I__10637\ : InMux
    port map (
            O => \N__51888\,
            I => \N__51882\
        );

    \I__10636\ : InMux
    port map (
            O => \N__51887\,
            I => \N__51882\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__51882\,
            I => \N__51878\
        );

    \I__10634\ : InMux
    port map (
            O => \N__51881\,
            I => \N__51875\
        );

    \I__10633\ : Odrv4
    port map (
            O => \N__51878\,
            I => \c0.n24528\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__51875\,
            I => \c0.n24528\
        );

    \I__10631\ : InMux
    port map (
            O => \N__51870\,
            I => \N__51867\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__51867\,
            I => \c0.n10_adj_4575\
        );

    \I__10629\ : InMux
    port map (
            O => \N__51864\,
            I => \N__51861\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__51861\,
            I => \c0.n23_adj_4598\
        );

    \I__10627\ : CascadeMux
    port map (
            O => \N__51858\,
            I => \N__51855\
        );

    \I__10626\ : InMux
    port map (
            O => \N__51855\,
            I => \N__51852\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__51852\,
            I => \N__51849\
        );

    \I__10624\ : Span4Mux_v
    port map (
            O => \N__51849\,
            I => \N__51846\
        );

    \I__10623\ : Odrv4
    port map (
            O => \N__51846\,
            I => \c0.n4_adj_4352\
        );

    \I__10622\ : InMux
    port map (
            O => \N__51843\,
            I => \N__51840\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__51840\,
            I => \c0.n23_adj_4353\
        );

    \I__10620\ : CascadeMux
    port map (
            O => \N__51837\,
            I => \c0.n23_adj_4353_cascade_\
        );

    \I__10619\ : InMux
    port map (
            O => \N__51834\,
            I => \N__51828\
        );

    \I__10618\ : InMux
    port map (
            O => \N__51833\,
            I => \N__51828\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__51828\,
            I => \c0.n15_adj_4344\
        );

    \I__10616\ : InMux
    port map (
            O => \N__51825\,
            I => \N__51822\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__51822\,
            I => \c0.n21428\
        );

    \I__10614\ : CascadeMux
    port map (
            O => \N__51819\,
            I => \c0.n11_adj_4438_cascade_\
        );

    \I__10613\ : InMux
    port map (
            O => \N__51816\,
            I => \N__51813\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__51813\,
            I => \c0.n16_adj_4437\
        );

    \I__10611\ : InMux
    port map (
            O => \N__51810\,
            I => \N__51804\
        );

    \I__10610\ : InMux
    port map (
            O => \N__51809\,
            I => \N__51804\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__51804\,
            I => \c0.n22420\
        );

    \I__10608\ : CascadeMux
    port map (
            O => \N__51801\,
            I => \N__51797\
        );

    \I__10607\ : CascadeMux
    port map (
            O => \N__51800\,
            I => \N__51794\
        );

    \I__10606\ : InMux
    port map (
            O => \N__51797\,
            I => \N__51791\
        );

    \I__10605\ : InMux
    port map (
            O => \N__51794\,
            I => \N__51788\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__51791\,
            I => \N__51785\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__51788\,
            I => \c0.data_in_frame_28_0\
        );

    \I__10602\ : Odrv4
    port map (
            O => \N__51785\,
            I => \c0.data_in_frame_28_0\
        );

    \I__10601\ : InMux
    port map (
            O => \N__51780\,
            I => \N__51774\
        );

    \I__10600\ : InMux
    port map (
            O => \N__51779\,
            I => \N__51770\
        );

    \I__10599\ : InMux
    port map (
            O => \N__51778\,
            I => \N__51767\
        );

    \I__10598\ : InMux
    port map (
            O => \N__51777\,
            I => \N__51764\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__51774\,
            I => \N__51761\
        );

    \I__10596\ : InMux
    port map (
            O => \N__51773\,
            I => \N__51758\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__51770\,
            I => \N__51751\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__51767\,
            I => \N__51751\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__51764\,
            I => \N__51751\
        );

    \I__10592\ : Span4Mux_v
    port map (
            O => \N__51761\,
            I => \N__51748\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__51758\,
            I => \c0.n21491\
        );

    \I__10590\ : Odrv12
    port map (
            O => \N__51751\,
            I => \c0.n21491\
        );

    \I__10589\ : Odrv4
    port map (
            O => \N__51748\,
            I => \c0.n21491\
        );

    \I__10588\ : CascadeMux
    port map (
            O => \N__51741\,
            I => \c0.n23187_cascade_\
        );

    \I__10587\ : CascadeMux
    port map (
            O => \N__51738\,
            I => \c0.n10_adj_4591_cascade_\
        );

    \I__10586\ : InMux
    port map (
            O => \N__51735\,
            I => \N__51732\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__51732\,
            I => \c0.n10_adj_4591\
        );

    \I__10584\ : InMux
    port map (
            O => \N__51729\,
            I => \N__51724\
        );

    \I__10583\ : InMux
    port map (
            O => \N__51728\,
            I => \N__51719\
        );

    \I__10582\ : InMux
    port map (
            O => \N__51727\,
            I => \N__51719\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__51724\,
            I => data_in_frame_21_2
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__51719\,
            I => data_in_frame_21_2
        );

    \I__10579\ : CascadeMux
    port map (
            O => \N__51714\,
            I => \c0.n12_adj_4606_cascade_\
        );

    \I__10578\ : CascadeMux
    port map (
            O => \N__51711\,
            I => \c0.n21325_cascade_\
        );

    \I__10577\ : InMux
    port map (
            O => \N__51708\,
            I => \N__51705\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__51705\,
            I => \N__51702\
        );

    \I__10575\ : Span4Mux_h
    port map (
            O => \N__51702\,
            I => \N__51699\
        );

    \I__10574\ : Span4Mux_v
    port map (
            O => \N__51699\,
            I => \N__51696\
        );

    \I__10573\ : Odrv4
    port map (
            O => \N__51696\,
            I => \c0.n24384\
        );

    \I__10572\ : CascadeMux
    port map (
            O => \N__51693\,
            I => \c0.n4_adj_4464_cascade_\
        );

    \I__10571\ : CascadeMux
    port map (
            O => \N__51690\,
            I => \c0.n21428_cascade_\
        );

    \I__10570\ : InMux
    port map (
            O => \N__51687\,
            I => \N__51684\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__51684\,
            I => \c0.n24_adj_4593\
        );

    \I__10568\ : InMux
    port map (
            O => \N__51681\,
            I => \N__51678\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__51678\,
            I => \c0.n154\
        );

    \I__10566\ : CascadeMux
    port map (
            O => \N__51675\,
            I => \N__51672\
        );

    \I__10565\ : InMux
    port map (
            O => \N__51672\,
            I => \N__51668\
        );

    \I__10564\ : InMux
    port map (
            O => \N__51671\,
            I => \N__51665\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__51668\,
            I => \N__51662\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__51665\,
            I => \c0.n15_adj_4301\
        );

    \I__10561\ : Odrv4
    port map (
            O => \N__51662\,
            I => \c0.n15_adj_4301\
        );

    \I__10560\ : InMux
    port map (
            O => \N__51657\,
            I => \N__51654\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__51654\,
            I => \c0.n21_adj_4605\
        );

    \I__10558\ : CascadeMux
    port map (
            O => \N__51651\,
            I => \N__51648\
        );

    \I__10557\ : InMux
    port map (
            O => \N__51648\,
            I => \N__51645\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__51645\,
            I => \c0.n19_adj_4604\
        );

    \I__10555\ : InMux
    port map (
            O => \N__51642\,
            I => \N__51639\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__51639\,
            I => \N__51636\
        );

    \I__10553\ : Odrv12
    port map (
            O => \N__51636\,
            I => \c0.n16_adj_4256\
        );

    \I__10552\ : InMux
    port map (
            O => \N__51633\,
            I => \N__51630\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__51630\,
            I => \c0.n22\
        );

    \I__10550\ : InMux
    port map (
            O => \N__51627\,
            I => \N__51623\
        );

    \I__10549\ : InMux
    port map (
            O => \N__51626\,
            I => \N__51620\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__51623\,
            I => \N__51617\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__51620\,
            I => \N__51614\
        );

    \I__10546\ : Span4Mux_v
    port map (
            O => \N__51617\,
            I => \N__51610\
        );

    \I__10545\ : Sp12to4
    port map (
            O => \N__51614\,
            I => \N__51607\
        );

    \I__10544\ : InMux
    port map (
            O => \N__51613\,
            I => \N__51604\
        );

    \I__10543\ : Odrv4
    port map (
            O => \N__51610\,
            I => \c0.n13280\
        );

    \I__10542\ : Odrv12
    port map (
            O => \N__51607\,
            I => \c0.n13280\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__51604\,
            I => \c0.n13280\
        );

    \I__10540\ : CascadeMux
    port map (
            O => \N__51597\,
            I => \c0.n13_cascade_\
        );

    \I__10539\ : InMux
    port map (
            O => \N__51594\,
            I => \N__51591\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__51591\,
            I => \N__51588\
        );

    \I__10537\ : Odrv12
    port map (
            O => \N__51588\,
            I => \c0.n20_adj_4222\
        );

    \I__10536\ : InMux
    port map (
            O => \N__51585\,
            I => \N__51582\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__51582\,
            I => \N__51578\
        );

    \I__10534\ : InMux
    port map (
            O => \N__51581\,
            I => \N__51575\
        );

    \I__10533\ : Span4Mux_v
    port map (
            O => \N__51578\,
            I => \N__51568\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__51575\,
            I => \N__51568\
        );

    \I__10531\ : InMux
    port map (
            O => \N__51574\,
            I => \N__51565\
        );

    \I__10530\ : InMux
    port map (
            O => \N__51573\,
            I => \N__51559\
        );

    \I__10529\ : Span4Mux_v
    port map (
            O => \N__51568\,
            I => \N__51556\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__51565\,
            I => \N__51553\
        );

    \I__10527\ : InMux
    port map (
            O => \N__51564\,
            I => \N__51550\
        );

    \I__10526\ : InMux
    port map (
            O => \N__51563\,
            I => \N__51547\
        );

    \I__10525\ : InMux
    port map (
            O => \N__51562\,
            I => \N__51544\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__51559\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10523\ : Odrv4
    port map (
            O => \N__51556\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10522\ : Odrv12
    port map (
            O => \N__51553\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__51550\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__51547\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__51544\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10518\ : CascadeMux
    port map (
            O => \N__51531\,
            I => \c0.n22_adj_4223_cascade_\
        );

    \I__10517\ : CascadeMux
    port map (
            O => \N__51528\,
            I => \c0.n21_adj_4225_cascade_\
        );

    \I__10516\ : CascadeMux
    port map (
            O => \N__51525\,
            I => \c0.n10_adj_4277_cascade_\
        );

    \I__10515\ : CascadeMux
    port map (
            O => \N__51522\,
            I => \N__51518\
        );

    \I__10514\ : InMux
    port map (
            O => \N__51521\,
            I => \N__51510\
        );

    \I__10513\ : InMux
    port map (
            O => \N__51518\,
            I => \N__51510\
        );

    \I__10512\ : InMux
    port map (
            O => \N__51517\,
            I => \N__51510\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__51510\,
            I => \c0.n23116\
        );

    \I__10510\ : InMux
    port map (
            O => \N__51507\,
            I => \N__51504\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__51504\,
            I => \N__51501\
        );

    \I__10508\ : Span4Mux_h
    port map (
            O => \N__51501\,
            I => \N__51498\
        );

    \I__10507\ : Span4Mux_v
    port map (
            O => \N__51498\,
            I => \N__51495\
        );

    \I__10506\ : Odrv4
    port map (
            O => \N__51495\,
            I => \c0.n128\
        );

    \I__10505\ : CascadeMux
    port map (
            O => \N__51492\,
            I => \c0.n129_cascade_\
        );

    \I__10504\ : InMux
    port map (
            O => \N__51489\,
            I => \N__51486\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__51486\,
            I => \c0.n11_adj_4614\
        );

    \I__10502\ : CascadeMux
    port map (
            O => \N__51483\,
            I => \c0.n16_adj_4613_cascade_\
        );

    \I__10501\ : InMux
    port map (
            O => \N__51480\,
            I => \N__51477\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__51477\,
            I => \N__51474\
        );

    \I__10499\ : Span4Mux_v
    port map (
            O => \N__51474\,
            I => \N__51471\
        );

    \I__10498\ : Span4Mux_v
    port map (
            O => \N__51471\,
            I => \N__51468\
        );

    \I__10497\ : Span4Mux_h
    port map (
            O => \N__51468\,
            I => \N__51461\
        );

    \I__10496\ : InMux
    port map (
            O => \N__51467\,
            I => \N__51455\
        );

    \I__10495\ : InMux
    port map (
            O => \N__51466\,
            I => \N__51455\
        );

    \I__10494\ : CascadeMux
    port map (
            O => \N__51465\,
            I => \N__51452\
        );

    \I__10493\ : CascadeMux
    port map (
            O => \N__51464\,
            I => \N__51449\
        );

    \I__10492\ : Span4Mux_v
    port map (
            O => \N__51461\,
            I => \N__51443\
        );

    \I__10491\ : InMux
    port map (
            O => \N__51460\,
            I => \N__51440\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__51455\,
            I => \N__51436\
        );

    \I__10489\ : InMux
    port map (
            O => \N__51452\,
            I => \N__51433\
        );

    \I__10488\ : InMux
    port map (
            O => \N__51449\,
            I => \N__51428\
        );

    \I__10487\ : InMux
    port map (
            O => \N__51448\,
            I => \N__51428\
        );

    \I__10486\ : CascadeMux
    port map (
            O => \N__51447\,
            I => \N__51425\
        );

    \I__10485\ : CascadeMux
    port map (
            O => \N__51446\,
            I => \N__51421\
        );

    \I__10484\ : Span4Mux_h
    port map (
            O => \N__51443\,
            I => \N__51415\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__51440\,
            I => \N__51412\
        );

    \I__10482\ : InMux
    port map (
            O => \N__51439\,
            I => \N__51409\
        );

    \I__10481\ : Span4Mux_v
    port map (
            O => \N__51436\,
            I => \N__51402\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__51433\,
            I => \N__51402\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__51428\,
            I => \N__51402\
        );

    \I__10478\ : InMux
    port map (
            O => \N__51425\,
            I => \N__51397\
        );

    \I__10477\ : InMux
    port map (
            O => \N__51424\,
            I => \N__51397\
        );

    \I__10476\ : InMux
    port map (
            O => \N__51421\,
            I => \N__51390\
        );

    \I__10475\ : InMux
    port map (
            O => \N__51420\,
            I => \N__51390\
        );

    \I__10474\ : InMux
    port map (
            O => \N__51419\,
            I => \N__51390\
        );

    \I__10473\ : InMux
    port map (
            O => \N__51418\,
            I => \N__51387\
        );

    \I__10472\ : Odrv4
    port map (
            O => \N__51415\,
            I => data_in_frame_1_3
        );

    \I__10471\ : Odrv4
    port map (
            O => \N__51412\,
            I => data_in_frame_1_3
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__51409\,
            I => data_in_frame_1_3
        );

    \I__10469\ : Odrv4
    port map (
            O => \N__51402\,
            I => data_in_frame_1_3
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__51397\,
            I => data_in_frame_1_3
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__51390\,
            I => data_in_frame_1_3
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__51387\,
            I => data_in_frame_1_3
        );

    \I__10465\ : InMux
    port map (
            O => \N__51372\,
            I => \N__51369\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__51369\,
            I => \N__51366\
        );

    \I__10463\ : Odrv12
    port map (
            O => \N__51366\,
            I => \c0.n126\
        );

    \I__10462\ : InMux
    port map (
            O => \N__51363\,
            I => \N__51360\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__51360\,
            I => \c0.n123\
        );

    \I__10460\ : CascadeMux
    port map (
            O => \N__51357\,
            I => \c0.n144_cascade_\
        );

    \I__10459\ : InMux
    port map (
            O => \N__51354\,
            I => \N__51351\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__51351\,
            I => \N__51348\
        );

    \I__10457\ : Odrv4
    port map (
            O => \N__51348\,
            I => \c0.n7_adj_4221\
        );

    \I__10456\ : InMux
    port map (
            O => \N__51345\,
            I => \N__51342\
        );

    \I__10455\ : LocalMux
    port map (
            O => \N__51342\,
            I => \c0.n16_adj_4641\
        );

    \I__10454\ : CascadeMux
    port map (
            O => \N__51339\,
            I => \c0.n23116_cascade_\
        );

    \I__10453\ : InMux
    port map (
            O => \N__51336\,
            I => \N__51332\
        );

    \I__10452\ : InMux
    port map (
            O => \N__51335\,
            I => \N__51329\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__51332\,
            I => \N__51323\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__51329\,
            I => \N__51323\
        );

    \I__10449\ : InMux
    port map (
            O => \N__51328\,
            I => \N__51320\
        );

    \I__10448\ : Span4Mux_v
    port map (
            O => \N__51323\,
            I => \N__51317\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__51320\,
            I => \c0.n7_adj_4337\
        );

    \I__10446\ : Odrv4
    port map (
            O => \N__51317\,
            I => \c0.n7_adj_4337\
        );

    \I__10445\ : CascadeMux
    port map (
            O => \N__51312\,
            I => \c0.n38_adj_4573_cascade_\
        );

    \I__10444\ : InMux
    port map (
            O => \N__51309\,
            I => \N__51306\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__51306\,
            I => \N__51303\
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__51303\,
            I => \c0.n44_adj_4744\
        );

    \I__10441\ : CascadeMux
    port map (
            O => \N__51300\,
            I => \c0.n43_adj_4574_cascade_\
        );

    \I__10440\ : InMux
    port map (
            O => \N__51297\,
            I => \N__51294\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__51294\,
            I => \c0.n41_adj_4745\
        );

    \I__10438\ : InMux
    port map (
            O => \N__51291\,
            I => \N__51288\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__51288\,
            I => \N__51285\
        );

    \I__10436\ : Odrv4
    port map (
            O => \N__51285\,
            I => \c0.n24048\
        );

    \I__10435\ : CascadeMux
    port map (
            O => \N__51282\,
            I => \c0.n24048_cascade_\
        );

    \I__10434\ : InMux
    port map (
            O => \N__51279\,
            I => \N__51276\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__51276\,
            I => \N__51272\
        );

    \I__10432\ : InMux
    port map (
            O => \N__51275\,
            I => \N__51269\
        );

    \I__10431\ : Odrv4
    port map (
            O => \N__51272\,
            I => \c0.n109\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__51269\,
            I => \c0.n109\
        );

    \I__10429\ : CascadeMux
    port map (
            O => \N__51264\,
            I => \N__51261\
        );

    \I__10428\ : InMux
    port map (
            O => \N__51261\,
            I => \N__51258\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__51258\,
            I => \N__51255\
        );

    \I__10426\ : Odrv4
    port map (
            O => \N__51255\,
            I => \c0.n23_adj_4590\
        );

    \I__10425\ : InMux
    port map (
            O => \N__51252\,
            I => \N__51249\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__51249\,
            I => \N__51246\
        );

    \I__10423\ : Span4Mux_h
    port map (
            O => \N__51246\,
            I => \N__51243\
        );

    \I__10422\ : Odrv4
    port map (
            O => \N__51243\,
            I => \c0.n29_adj_4734\
        );

    \I__10421\ : CascadeMux
    port map (
            O => \N__51240\,
            I => \c0.n20_adj_4290_cascade_\
        );

    \I__10420\ : InMux
    port map (
            O => \N__51237\,
            I => \N__51234\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__51234\,
            I => \N__51229\
        );

    \I__10418\ : InMux
    port map (
            O => \N__51233\,
            I => \N__51224\
        );

    \I__10417\ : InMux
    port map (
            O => \N__51232\,
            I => \N__51224\
        );

    \I__10416\ : Span4Mux_v
    port map (
            O => \N__51229\,
            I => \N__51220\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__51224\,
            I => \N__51213\
        );

    \I__10414\ : InMux
    port map (
            O => \N__51223\,
            I => \N__51208\
        );

    \I__10413\ : Sp12to4
    port map (
            O => \N__51220\,
            I => \N__51203\
        );

    \I__10412\ : InMux
    port map (
            O => \N__51219\,
            I => \N__51200\
        );

    \I__10411\ : InMux
    port map (
            O => \N__51218\,
            I => \N__51197\
        );

    \I__10410\ : InMux
    port map (
            O => \N__51217\,
            I => \N__51192\
        );

    \I__10409\ : InMux
    port map (
            O => \N__51216\,
            I => \N__51192\
        );

    \I__10408\ : Span4Mux_v
    port map (
            O => \N__51213\,
            I => \N__51189\
        );

    \I__10407\ : InMux
    port map (
            O => \N__51212\,
            I => \N__51184\
        );

    \I__10406\ : InMux
    port map (
            O => \N__51211\,
            I => \N__51184\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__51208\,
            I => \N__51181\
        );

    \I__10404\ : InMux
    port map (
            O => \N__51207\,
            I => \N__51176\
        );

    \I__10403\ : InMux
    port map (
            O => \N__51206\,
            I => \N__51176\
        );

    \I__10402\ : Odrv12
    port map (
            O => \N__51203\,
            I => data_in_frame_1_1
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__51200\,
            I => data_in_frame_1_1
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__51197\,
            I => data_in_frame_1_1
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__51192\,
            I => data_in_frame_1_1
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__51189\,
            I => data_in_frame_1_1
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__51184\,
            I => data_in_frame_1_1
        );

    \I__10396\ : Odrv4
    port map (
            O => \N__51181\,
            I => data_in_frame_1_1
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__51176\,
            I => data_in_frame_1_1
        );

    \I__10394\ : InMux
    port map (
            O => \N__51159\,
            I => \N__51156\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__51156\,
            I => \N__51153\
        );

    \I__10392\ : Odrv12
    port map (
            O => \N__51153\,
            I => \c0.n51\
        );

    \I__10391\ : InMux
    port map (
            O => \N__51150\,
            I => \N__51144\
        );

    \I__10390\ : InMux
    port map (
            O => \N__51149\,
            I => \N__51144\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__51144\,
            I => \c0.n29\
        );

    \I__10388\ : CascadeMux
    port map (
            O => \N__51141\,
            I => \c0.n51_cascade_\
        );

    \I__10387\ : InMux
    port map (
            O => \N__51138\,
            I => \N__51131\
        );

    \I__10386\ : InMux
    port map (
            O => \N__51137\,
            I => \N__51131\
        );

    \I__10385\ : InMux
    port map (
            O => \N__51136\,
            I => \N__51128\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__51131\,
            I => \N__51125\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__51128\,
            I => \c0.n22_adj_4647\
        );

    \I__10382\ : Odrv4
    port map (
            O => \N__51125\,
            I => \c0.n22_adj_4647\
        );

    \I__10381\ : CascadeMux
    port map (
            O => \N__51120\,
            I => \c0.n102_cascade_\
        );

    \I__10380\ : InMux
    port map (
            O => \N__51117\,
            I => \N__51114\
        );

    \I__10379\ : LocalMux
    port map (
            O => \N__51114\,
            I => \c0.n32\
        );

    \I__10378\ : CascadeMux
    port map (
            O => \N__51111\,
            I => \c0.n16_adj_4256_cascade_\
        );

    \I__10377\ : CascadeMux
    port map (
            O => \N__51108\,
            I => \N__51105\
        );

    \I__10376\ : InMux
    port map (
            O => \N__51105\,
            I => \N__51102\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__51102\,
            I => \c0.n9_adj_4279\
        );

    \I__10374\ : CascadeMux
    port map (
            O => \N__51099\,
            I => \N__51096\
        );

    \I__10373\ : InMux
    port map (
            O => \N__51096\,
            I => \N__51093\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__51093\,
            I => \N__51089\
        );

    \I__10371\ : InMux
    port map (
            O => \N__51092\,
            I => \N__51086\
        );

    \I__10370\ : Span4Mux_h
    port map (
            O => \N__51089\,
            I => \N__51082\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__51086\,
            I => \N__51079\
        );

    \I__10368\ : InMux
    port map (
            O => \N__51085\,
            I => \N__51076\
        );

    \I__10367\ : Odrv4
    port map (
            O => \N__51082\,
            I => \c0.n13141\
        );

    \I__10366\ : Odrv12
    port map (
            O => \N__51079\,
            I => \c0.n13141\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__51076\,
            I => \c0.n13141\
        );

    \I__10364\ : CascadeMux
    port map (
            O => \N__51069\,
            I => \c0.n9_adj_4279_cascade_\
        );

    \I__10363\ : CascadeMux
    port map (
            O => \N__51066\,
            I => \c0.n23574_cascade_\
        );

    \I__10362\ : InMux
    port map (
            O => \N__51063\,
            I => \N__51060\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__51060\,
            I => \c0.n11_adj_4257\
        );

    \I__10360\ : CascadeMux
    port map (
            O => \N__51057\,
            I => \c0.n38_adj_4285_cascade_\
        );

    \I__10359\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51051\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__51051\,
            I => \c0.n26_adj_4289\
        );

    \I__10357\ : CascadeMux
    port map (
            O => \N__51048\,
            I => \c0.n26_adj_4289_cascade_\
        );

    \I__10356\ : InMux
    port map (
            O => \N__51045\,
            I => \N__51041\
        );

    \I__10355\ : InMux
    port map (
            O => \N__51044\,
            I => \N__51038\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__51041\,
            I => \N__51035\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__51038\,
            I => \c0.data_out_frame_0__7__N_2626\
        );

    \I__10352\ : Odrv4
    port map (
            O => \N__51035\,
            I => \c0.data_out_frame_0__7__N_2626\
        );

    \I__10351\ : InMux
    port map (
            O => \N__51030\,
            I => \N__51024\
        );

    \I__10350\ : InMux
    port map (
            O => \N__51029\,
            I => \N__51024\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__51024\,
            I => \c0.n20_adj_4290\
        );

    \I__10348\ : InMux
    port map (
            O => \N__51021\,
            I => \N__51018\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__51018\,
            I => \c0.n12_adj_4657\
        );

    \I__10346\ : CascadeMux
    port map (
            O => \N__51015\,
            I => \N__51012\
        );

    \I__10345\ : InMux
    port map (
            O => \N__51012\,
            I => \N__51009\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__51009\,
            I => \N__51006\
        );

    \I__10343\ : Span4Mux_h
    port map (
            O => \N__51006\,
            I => \N__51003\
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__51003\,
            I => \c0.n23_adj_4648\
        );

    \I__10341\ : InMux
    port map (
            O => \N__51000\,
            I => \N__50997\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__50997\,
            I => \c0.n39_adj_4737\
        );

    \I__10339\ : InMux
    port map (
            O => \N__50994\,
            I => \N__50991\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__50991\,
            I => \c0.n38_adj_4736\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__50988\,
            I => \N__50985\
        );

    \I__10336\ : InMux
    port map (
            O => \N__50985\,
            I => \N__50979\
        );

    \I__10335\ : InMux
    port map (
            O => \N__50984\,
            I => \N__50979\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__50979\,
            I => \c0.n23562\
        );

    \I__10333\ : CascadeMux
    port map (
            O => \N__50976\,
            I => \c0.n23562_cascade_\
        );

    \I__10332\ : InMux
    port map (
            O => \N__50973\,
            I => \N__50966\
        );

    \I__10331\ : InMux
    port map (
            O => \N__50972\,
            I => \N__50961\
        );

    \I__10330\ : InMux
    port map (
            O => \N__50971\,
            I => \N__50961\
        );

    \I__10329\ : InMux
    port map (
            O => \N__50970\,
            I => \N__50956\
        );

    \I__10328\ : InMux
    port map (
            O => \N__50969\,
            I => \N__50956\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__50966\,
            I => data_in_frame_5_5
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__50961\,
            I => data_in_frame_5_5
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__50956\,
            I => data_in_frame_5_5
        );

    \I__10324\ : CascadeMux
    port map (
            O => \N__50949\,
            I => \N__50946\
        );

    \I__10323\ : InMux
    port map (
            O => \N__50946\,
            I => \N__50937\
        );

    \I__10322\ : InMux
    port map (
            O => \N__50945\,
            I => \N__50932\
        );

    \I__10321\ : InMux
    port map (
            O => \N__50944\,
            I => \N__50932\
        );

    \I__10320\ : InMux
    port map (
            O => \N__50943\,
            I => \N__50927\
        );

    \I__10319\ : InMux
    port map (
            O => \N__50942\,
            I => \N__50927\
        );

    \I__10318\ : InMux
    port map (
            O => \N__50941\,
            I => \N__50922\
        );

    \I__10317\ : InMux
    port map (
            O => \N__50940\,
            I => \N__50922\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__50937\,
            I => \c0.data_in_frame_3_4\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__50932\,
            I => \c0.data_in_frame_3_4\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__50927\,
            I => \c0.data_in_frame_3_4\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__50922\,
            I => \c0.data_in_frame_3_4\
        );

    \I__10312\ : CascadeMux
    port map (
            O => \N__50913\,
            I => \N__50905\
        );

    \I__10311\ : CascadeMux
    port map (
            O => \N__50912\,
            I => \N__50901\
        );

    \I__10310\ : CascadeMux
    port map (
            O => \N__50911\,
            I => \N__50898\
        );

    \I__10309\ : CascadeMux
    port map (
            O => \N__50910\,
            I => \N__50895\
        );

    \I__10308\ : InMux
    port map (
            O => \N__50909\,
            I => \N__50892\
        );

    \I__10307\ : CascadeMux
    port map (
            O => \N__50908\,
            I => \N__50889\
        );

    \I__10306\ : InMux
    port map (
            O => \N__50905\,
            I => \N__50886\
        );

    \I__10305\ : CascadeMux
    port map (
            O => \N__50904\,
            I => \N__50883\
        );

    \I__10304\ : InMux
    port map (
            O => \N__50901\,
            I => \N__50880\
        );

    \I__10303\ : InMux
    port map (
            O => \N__50898\,
            I => \N__50877\
        );

    \I__10302\ : InMux
    port map (
            O => \N__50895\,
            I => \N__50874\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__50892\,
            I => \N__50871\
        );

    \I__10300\ : InMux
    port map (
            O => \N__50889\,
            I => \N__50868\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__50886\,
            I => \N__50861\
        );

    \I__10298\ : InMux
    port map (
            O => \N__50883\,
            I => \N__50858\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__50880\,
            I => \N__50851\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__50877\,
            I => \N__50851\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__50874\,
            I => \N__50851\
        );

    \I__10294\ : Span4Mux_s3_v
    port map (
            O => \N__50871\,
            I => \N__50848\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__50868\,
            I => \N__50845\
        );

    \I__10292\ : InMux
    port map (
            O => \N__50867\,
            I => \N__50842\
        );

    \I__10291\ : InMux
    port map (
            O => \N__50866\,
            I => \N__50837\
        );

    \I__10290\ : InMux
    port map (
            O => \N__50865\,
            I => \N__50837\
        );

    \I__10289\ : CascadeMux
    port map (
            O => \N__50864\,
            I => \N__50834\
        );

    \I__10288\ : Span4Mux_v
    port map (
            O => \N__50861\,
            I => \N__50829\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__50858\,
            I => \N__50829\
        );

    \I__10286\ : Span4Mux_h
    port map (
            O => \N__50851\,
            I => \N__50826\
        );

    \I__10285\ : Span4Mux_h
    port map (
            O => \N__50848\,
            I => \N__50822\
        );

    \I__10284\ : Span4Mux_v
    port map (
            O => \N__50845\,
            I => \N__50817\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__50842\,
            I => \N__50817\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__50837\,
            I => \N__50814\
        );

    \I__10281\ : InMux
    port map (
            O => \N__50834\,
            I => \N__50811\
        );

    \I__10280\ : Span4Mux_v
    port map (
            O => \N__50829\,
            I => \N__50808\
        );

    \I__10279\ : Span4Mux_h
    port map (
            O => \N__50826\,
            I => \N__50805\
        );

    \I__10278\ : InMux
    port map (
            O => \N__50825\,
            I => \N__50802\
        );

    \I__10277\ : Sp12to4
    port map (
            O => \N__50822\,
            I => \N__50799\
        );

    \I__10276\ : Span4Mux_h
    port map (
            O => \N__50817\,
            I => \N__50796\
        );

    \I__10275\ : Span4Mux_v
    port map (
            O => \N__50814\,
            I => \N__50793\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__50811\,
            I => \N__50790\
        );

    \I__10273\ : Span4Mux_h
    port map (
            O => \N__50808\,
            I => \N__50787\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__50805\,
            I => \N__50782\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__50802\,
            I => \N__50782\
        );

    \I__10270\ : Span12Mux_h
    port map (
            O => \N__50799\,
            I => \N__50779\
        );

    \I__10269\ : Span4Mux_h
    port map (
            O => \N__50796\,
            I => \N__50776\
        );

    \I__10268\ : Span4Mux_h
    port map (
            O => \N__50793\,
            I => \N__50773\
        );

    \I__10267\ : Sp12to4
    port map (
            O => \N__50790\,
            I => \N__50770\
        );

    \I__10266\ : Span4Mux_h
    port map (
            O => \N__50787\,
            I => \N__50767\
        );

    \I__10265\ : Sp12to4
    port map (
            O => \N__50782\,
            I => \N__50760\
        );

    \I__10264\ : Span12Mux_v
    port map (
            O => \N__50779\,
            I => \N__50760\
        );

    \I__10263\ : Sp12to4
    port map (
            O => \N__50776\,
            I => \N__50760\
        );

    \I__10262\ : Span4Mux_h
    port map (
            O => \N__50773\,
            I => \N__50757\
        );

    \I__10261\ : Span12Mux_h
    port map (
            O => \N__50770\,
            I => \N__50754\
        );

    \I__10260\ : Span4Mux_h
    port map (
            O => \N__50767\,
            I => \N__50751\
        );

    \I__10259\ : Span12Mux_v
    port map (
            O => \N__50760\,
            I => \N__50748\
        );

    \I__10258\ : Span4Mux_v
    port map (
            O => \N__50757\,
            I => \N__50745\
        );

    \I__10257\ : Odrv12
    port map (
            O => \N__50754\,
            I => \r_Rx_Data\
        );

    \I__10256\ : Odrv4
    port map (
            O => \N__50751\,
            I => \r_Rx_Data\
        );

    \I__10255\ : Odrv12
    port map (
            O => \N__50748\,
            I => \r_Rx_Data\
        );

    \I__10254\ : Odrv4
    port map (
            O => \N__50745\,
            I => \r_Rx_Data\
        );

    \I__10253\ : CascadeMux
    port map (
            O => \N__50736\,
            I => \n4_cascade_\
        );

    \I__10252\ : InMux
    port map (
            O => \N__50733\,
            I => \N__50730\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__50730\,
            I => \N__50727\
        );

    \I__10250\ : Span4Mux_s2_v
    port map (
            O => \N__50727\,
            I => \N__50723\
        );

    \I__10249\ : InMux
    port map (
            O => \N__50726\,
            I => \N__50720\
        );

    \I__10248\ : Sp12to4
    port map (
            O => \N__50723\,
            I => \N__50715\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__50720\,
            I => \N__50712\
        );

    \I__10246\ : InMux
    port map (
            O => \N__50719\,
            I => \N__50709\
        );

    \I__10245\ : InMux
    port map (
            O => \N__50718\,
            I => \N__50706\
        );

    \I__10244\ : Span12Mux_h
    port map (
            O => \N__50715\,
            I => \N__50703\
        );

    \I__10243\ : Span4Mux_h
    port map (
            O => \N__50712\,
            I => \N__50698\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__50709\,
            I => \N__50698\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__50706\,
            I => \N__50695\
        );

    \I__10240\ : Span12Mux_v
    port map (
            O => \N__50703\,
            I => \N__50692\
        );

    \I__10239\ : Span4Mux_v
    port map (
            O => \N__50698\,
            I => \N__50689\
        );

    \I__10238\ : Span4Mux_v
    port map (
            O => \N__50695\,
            I => \N__50686\
        );

    \I__10237\ : Odrv12
    port map (
            O => \N__50692\,
            I => n12904
        );

    \I__10236\ : Odrv4
    port map (
            O => \N__50689\,
            I => n12904
        );

    \I__10235\ : Odrv4
    port map (
            O => \N__50686\,
            I => n12904
        );

    \I__10234\ : InMux
    port map (
            O => \N__50679\,
            I => \N__50676\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__50676\,
            I => \N__50673\
        );

    \I__10232\ : Span12Mux_s4_v
    port map (
            O => \N__50673\,
            I => \N__50670\
        );

    \I__10231\ : Span12Mux_v
    port map (
            O => \N__50670\,
            I => \N__50667\
        );

    \I__10230\ : Odrv12
    port map (
            O => \N__50667\,
            I => \c0.rx.n14277\
        );

    \I__10229\ : InMux
    port map (
            O => \N__50664\,
            I => \N__50661\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__50661\,
            I => \N__50658\
        );

    \I__10227\ : Sp12to4
    port map (
            O => \N__50658\,
            I => \N__50655\
        );

    \I__10226\ : Span12Mux_s3_v
    port map (
            O => \N__50655\,
            I => \N__50652\
        );

    \I__10225\ : Span12Mux_v
    port map (
            O => \N__50652\,
            I => \N__50647\
        );

    \I__10224\ : InMux
    port map (
            O => \N__50651\,
            I => \N__50644\
        );

    \I__10223\ : InMux
    port map (
            O => \N__50650\,
            I => \N__50641\
        );

    \I__10222\ : Odrv12
    port map (
            O => \N__50647\,
            I => \c0.n12514\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__50644\,
            I => \c0.n12514\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__50641\,
            I => \c0.n12514\
        );

    \I__10219\ : InMux
    port map (
            O => \N__50634\,
            I => \N__50631\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__50631\,
            I => \N__50628\
        );

    \I__10217\ : Span4Mux_h
    port map (
            O => \N__50628\,
            I => \N__50625\
        );

    \I__10216\ : Span4Mux_v
    port map (
            O => \N__50625\,
            I => \N__50622\
        );

    \I__10215\ : Span4Mux_v
    port map (
            O => \N__50622\,
            I => \N__50617\
        );

    \I__10214\ : InMux
    port map (
            O => \N__50621\,
            I => \N__50614\
        );

    \I__10213\ : InMux
    port map (
            O => \N__50620\,
            I => \N__50611\
        );

    \I__10212\ : Span4Mux_v
    port map (
            O => \N__50617\,
            I => \N__50606\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__50614\,
            I => \N__50606\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__50611\,
            I => \N__50601\
        );

    \I__10209\ : Span4Mux_h
    port map (
            O => \N__50606\,
            I => \N__50601\
        );

    \I__10208\ : Odrv4
    port map (
            O => \N__50601\,
            I => \c0.n20641\
        );

    \I__10207\ : CascadeMux
    port map (
            O => \N__50598\,
            I => \N__50595\
        );

    \I__10206\ : InMux
    port map (
            O => \N__50595\,
            I => \N__50592\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__50592\,
            I => \N__50589\
        );

    \I__10204\ : Span4Mux_s3_v
    port map (
            O => \N__50589\,
            I => \N__50585\
        );

    \I__10203\ : InMux
    port map (
            O => \N__50588\,
            I => \N__50581\
        );

    \I__10202\ : Span4Mux_h
    port map (
            O => \N__50585\,
            I => \N__50578\
        );

    \I__10201\ : InMux
    port map (
            O => \N__50584\,
            I => \N__50575\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__50581\,
            I => \N__50571\
        );

    \I__10199\ : Span4Mux_h
    port map (
            O => \N__50578\,
            I => \N__50568\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__50575\,
            I => \N__50565\
        );

    \I__10197\ : InMux
    port map (
            O => \N__50574\,
            I => \N__50562\
        );

    \I__10196\ : Span4Mux_h
    port map (
            O => \N__50571\,
            I => \N__50559\
        );

    \I__10195\ : Sp12to4
    port map (
            O => \N__50568\,
            I => \N__50556\
        );

    \I__10194\ : Span4Mux_h
    port map (
            O => \N__50565\,
            I => \N__50553\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__50562\,
            I => \N__50550\
        );

    \I__10192\ : Odrv4
    port map (
            O => \N__50559\,
            I => \c0.n21391\
        );

    \I__10191\ : Odrv12
    port map (
            O => \N__50556\,
            I => \c0.n21391\
        );

    \I__10190\ : Odrv4
    port map (
            O => \N__50553\,
            I => \c0.n21391\
        );

    \I__10189\ : Odrv4
    port map (
            O => \N__50550\,
            I => \c0.n21391\
        );

    \I__10188\ : InMux
    port map (
            O => \N__50541\,
            I => \N__50538\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__50538\,
            I => \N__50535\
        );

    \I__10186\ : Span4Mux_h
    port map (
            O => \N__50535\,
            I => \N__50532\
        );

    \I__10185\ : Sp12to4
    port map (
            O => \N__50532\,
            I => \N__50529\
        );

    \I__10184\ : Span12Mux_v
    port map (
            O => \N__50529\,
            I => \N__50523\
        );

    \I__10183\ : InMux
    port map (
            O => \N__50528\,
            I => \N__50520\
        );

    \I__10182\ : InMux
    port map (
            O => \N__50527\,
            I => \N__50517\
        );

    \I__10181\ : InMux
    port map (
            O => \N__50526\,
            I => \N__50514\
        );

    \I__10180\ : Odrv12
    port map (
            O => \N__50523\,
            I => \c0.n21360\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__50520\,
            I => \c0.n21360\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__50517\,
            I => \c0.n21360\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__50514\,
            I => \c0.n21360\
        );

    \I__10176\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50502\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__50502\,
            I => \N__50499\
        );

    \I__10174\ : Span4Mux_h
    port map (
            O => \N__50499\,
            I => \N__50496\
        );

    \I__10173\ : Span4Mux_h
    port map (
            O => \N__50496\,
            I => \N__50493\
        );

    \I__10172\ : Sp12to4
    port map (
            O => \N__50493\,
            I => \N__50490\
        );

    \I__10171\ : Span12Mux_v
    port map (
            O => \N__50490\,
            I => \N__50487\
        );

    \I__10170\ : Odrv12
    port map (
            O => \N__50487\,
            I => \c0.n21_adj_4719\
        );

    \I__10169\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50477\
        );

    \I__10168\ : InMux
    port map (
            O => \N__50483\,
            I => \N__50474\
        );

    \I__10167\ : InMux
    port map (
            O => \N__50482\,
            I => \N__50467\
        );

    \I__10166\ : InMux
    port map (
            O => \N__50481\,
            I => \N__50467\
        );

    \I__10165\ : InMux
    port map (
            O => \N__50480\,
            I => \N__50455\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__50477\,
            I => \N__50448\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__50474\,
            I => \N__50448\
        );

    \I__10162\ : InMux
    port map (
            O => \N__50473\,
            I => \N__50445\
        );

    \I__10161\ : InMux
    port map (
            O => \N__50472\,
            I => \N__50442\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__50467\,
            I => \N__50439\
        );

    \I__10159\ : InMux
    port map (
            O => \N__50466\,
            I => \N__50433\
        );

    \I__10158\ : CascadeMux
    port map (
            O => \N__50465\,
            I => \N__50430\
        );

    \I__10157\ : InMux
    port map (
            O => \N__50464\,
            I => \N__50420\
        );

    \I__10156\ : InMux
    port map (
            O => \N__50463\,
            I => \N__50417\
        );

    \I__10155\ : InMux
    port map (
            O => \N__50462\,
            I => \N__50410\
        );

    \I__10154\ : InMux
    port map (
            O => \N__50461\,
            I => \N__50410\
        );

    \I__10153\ : InMux
    port map (
            O => \N__50460\,
            I => \N__50410\
        );

    \I__10152\ : InMux
    port map (
            O => \N__50459\,
            I => \N__50405\
        );

    \I__10151\ : InMux
    port map (
            O => \N__50458\,
            I => \N__50405\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__50455\,
            I => \N__50398\
        );

    \I__10149\ : InMux
    port map (
            O => \N__50454\,
            I => \N__50395\
        );

    \I__10148\ : InMux
    port map (
            O => \N__50453\,
            I => \N__50392\
        );

    \I__10147\ : Span4Mux_h
    port map (
            O => \N__50448\,
            I => \N__50386\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__50445\,
            I => \N__50386\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__50442\,
            I => \N__50381\
        );

    \I__10144\ : Span4Mux_v
    port map (
            O => \N__50439\,
            I => \N__50381\
        );

    \I__10143\ : InMux
    port map (
            O => \N__50438\,
            I => \N__50378\
        );

    \I__10142\ : InMux
    port map (
            O => \N__50437\,
            I => \N__50375\
        );

    \I__10141\ : InMux
    port map (
            O => \N__50436\,
            I => \N__50372\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__50433\,
            I => \N__50369\
        );

    \I__10139\ : InMux
    port map (
            O => \N__50430\,
            I => \N__50362\
        );

    \I__10138\ : InMux
    port map (
            O => \N__50429\,
            I => \N__50362\
        );

    \I__10137\ : InMux
    port map (
            O => \N__50428\,
            I => \N__50362\
        );

    \I__10136\ : InMux
    port map (
            O => \N__50427\,
            I => \N__50359\
        );

    \I__10135\ : InMux
    port map (
            O => \N__50426\,
            I => \N__50356\
        );

    \I__10134\ : InMux
    port map (
            O => \N__50425\,
            I => \N__50353\
        );

    \I__10133\ : InMux
    port map (
            O => \N__50424\,
            I => \N__50348\
        );

    \I__10132\ : InMux
    port map (
            O => \N__50423\,
            I => \N__50348\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__50420\,
            I => \N__50339\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__50417\,
            I => \N__50339\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__50410\,
            I => \N__50339\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__50405\,
            I => \N__50339\
        );

    \I__10127\ : InMux
    port map (
            O => \N__50404\,
            I => \N__50334\
        );

    \I__10126\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50334\
        );

    \I__10125\ : InMux
    port map (
            O => \N__50402\,
            I => \N__50329\
        );

    \I__10124\ : InMux
    port map (
            O => \N__50401\,
            I => \N__50329\
        );

    \I__10123\ : Span4Mux_v
    port map (
            O => \N__50398\,
            I => \N__50326\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__50395\,
            I => \N__50323\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__50392\,
            I => \N__50320\
        );

    \I__10120\ : InMux
    port map (
            O => \N__50391\,
            I => \N__50317\
        );

    \I__10119\ : Span4Mux_v
    port map (
            O => \N__50386\,
            I => \N__50314\
        );

    \I__10118\ : Span4Mux_v
    port map (
            O => \N__50381\,
            I => \N__50311\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__50378\,
            I => \N__50306\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__50375\,
            I => \N__50306\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__50372\,
            I => \N__50301\
        );

    \I__10114\ : Span4Mux_v
    port map (
            O => \N__50369\,
            I => \N__50301\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__50362\,
            I => \N__50286\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__50359\,
            I => \N__50286\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__50356\,
            I => \N__50286\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__50353\,
            I => \N__50286\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__50348\,
            I => \N__50286\
        );

    \I__10108\ : Span4Mux_v
    port map (
            O => \N__50339\,
            I => \N__50286\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__50334\,
            I => \N__50286\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__50329\,
            I => \N__50283\
        );

    \I__10105\ : Span4Mux_h
    port map (
            O => \N__50326\,
            I => \N__50278\
        );

    \I__10104\ : Span4Mux_v
    port map (
            O => \N__50323\,
            I => \N__50278\
        );

    \I__10103\ : Span4Mux_v
    port map (
            O => \N__50320\,
            I => \N__50273\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__50317\,
            I => \N__50273\
        );

    \I__10101\ : Span4Mux_v
    port map (
            O => \N__50314\,
            I => \N__50268\
        );

    \I__10100\ : Span4Mux_v
    port map (
            O => \N__50311\,
            I => \N__50268\
        );

    \I__10099\ : Span4Mux_v
    port map (
            O => \N__50306\,
            I => \N__50261\
        );

    \I__10098\ : Span4Mux_v
    port map (
            O => \N__50301\,
            I => \N__50261\
        );

    \I__10097\ : Span4Mux_v
    port map (
            O => \N__50286\,
            I => \N__50261\
        );

    \I__10096\ : Span4Mux_h
    port map (
            O => \N__50283\,
            I => \N__50256\
        );

    \I__10095\ : Span4Mux_v
    port map (
            O => \N__50278\,
            I => \N__50256\
        );

    \I__10094\ : Sp12to4
    port map (
            O => \N__50273\,
            I => \N__50253\
        );

    \I__10093\ : Span4Mux_h
    port map (
            O => \N__50268\,
            I => \N__50250\
        );

    \I__10092\ : Sp12to4
    port map (
            O => \N__50261\,
            I => \N__50247\
        );

    \I__10091\ : Span4Mux_v
    port map (
            O => \N__50256\,
            I => \N__50244\
        );

    \I__10090\ : Span12Mux_v
    port map (
            O => \N__50253\,
            I => \N__50241\
        );

    \I__10089\ : Sp12to4
    port map (
            O => \N__50250\,
            I => \N__50236\
        );

    \I__10088\ : Span12Mux_h
    port map (
            O => \N__50247\,
            I => \N__50236\
        );

    \I__10087\ : Span4Mux_v
    port map (
            O => \N__50244\,
            I => \N__50230\
        );

    \I__10086\ : Span12Mux_v
    port map (
            O => \N__50241\,
            I => \N__50227\
        );

    \I__10085\ : Span12Mux_v
    port map (
            O => \N__50236\,
            I => \N__50224\
        );

    \I__10084\ : InMux
    port map (
            O => \N__50235\,
            I => \N__50217\
        );

    \I__10083\ : InMux
    port map (
            O => \N__50234\,
            I => \N__50217\
        );

    \I__10082\ : InMux
    port map (
            O => \N__50233\,
            I => \N__50217\
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__50230\,
            I => rx_data_ready
        );

    \I__10080\ : Odrv12
    port map (
            O => \N__50227\,
            I => rx_data_ready
        );

    \I__10079\ : Odrv12
    port map (
            O => \N__50224\,
            I => rx_data_ready
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__50217\,
            I => rx_data_ready
        );

    \I__10077\ : InMux
    port map (
            O => \N__50208\,
            I => \N__50205\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__50205\,
            I => \N__50202\
        );

    \I__10075\ : Sp12to4
    port map (
            O => \N__50202\,
            I => \N__50199\
        );

    \I__10074\ : Span12Mux_h
    port map (
            O => \N__50199\,
            I => \N__50195\
        );

    \I__10073\ : InMux
    port map (
            O => \N__50198\,
            I => \N__50192\
        );

    \I__10072\ : Span12Mux_v
    port map (
            O => \N__50195\,
            I => \N__50189\
        );

    \I__10071\ : LocalMux
    port map (
            O => \N__50192\,
            I => \c0.FRAME_MATCHER_rx_data_ready_prev\
        );

    \I__10070\ : Odrv12
    port map (
            O => \N__50189\,
            I => \c0.FRAME_MATCHER_rx_data_ready_prev\
        );

    \I__10069\ : CascadeMux
    port map (
            O => \N__50184\,
            I => \N__50180\
        );

    \I__10068\ : CascadeMux
    port map (
            O => \N__50183\,
            I => \N__50174\
        );

    \I__10067\ : InMux
    port map (
            O => \N__50180\,
            I => \N__50169\
        );

    \I__10066\ : InMux
    port map (
            O => \N__50179\,
            I => \N__50169\
        );

    \I__10065\ : CascadeMux
    port map (
            O => \N__50178\,
            I => \N__50166\
        );

    \I__10064\ : CascadeMux
    port map (
            O => \N__50177\,
            I => \N__50163\
        );

    \I__10063\ : InMux
    port map (
            O => \N__50174\,
            I => \N__50158\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__50169\,
            I => \N__50154\
        );

    \I__10061\ : InMux
    port map (
            O => \N__50166\,
            I => \N__50150\
        );

    \I__10060\ : InMux
    port map (
            O => \N__50163\,
            I => \N__50147\
        );

    \I__10059\ : CascadeMux
    port map (
            O => \N__50162\,
            I => \N__50144\
        );

    \I__10058\ : InMux
    port map (
            O => \N__50161\,
            I => \N__50141\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__50158\,
            I => \N__50138\
        );

    \I__10056\ : CascadeMux
    port map (
            O => \N__50157\,
            I => \N__50135\
        );

    \I__10055\ : Span12Mux_h
    port map (
            O => \N__50154\,
            I => \N__50132\
        );

    \I__10054\ : InMux
    port map (
            O => \N__50153\,
            I => \N__50129\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__50150\,
            I => \N__50126\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__50147\,
            I => \N__50123\
        );

    \I__10051\ : InMux
    port map (
            O => \N__50144\,
            I => \N__50120\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__50141\,
            I => \N__50117\
        );

    \I__10049\ : Span4Mux_v
    port map (
            O => \N__50138\,
            I => \N__50114\
        );

    \I__10048\ : InMux
    port map (
            O => \N__50135\,
            I => \N__50111\
        );

    \I__10047\ : Span12Mux_v
    port map (
            O => \N__50132\,
            I => \N__50108\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__50129\,
            I => \N__50103\
        );

    \I__10045\ : Span4Mux_h
    port map (
            O => \N__50126\,
            I => \N__50100\
        );

    \I__10044\ : Span4Mux_h
    port map (
            O => \N__50123\,
            I => \N__50095\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__50120\,
            I => \N__50095\
        );

    \I__10042\ : Span4Mux_v
    port map (
            O => \N__50117\,
            I => \N__50090\
        );

    \I__10041\ : Span4Mux_v
    port map (
            O => \N__50114\,
            I => \N__50090\
        );

    \I__10040\ : LocalMux
    port map (
            O => \N__50111\,
            I => \N__50087\
        );

    \I__10039\ : Span12Mux_v
    port map (
            O => \N__50108\,
            I => \N__50084\
        );

    \I__10038\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50079\
        );

    \I__10037\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50079\
        );

    \I__10036\ : Span12Mux_h
    port map (
            O => \N__50103\,
            I => \N__50076\
        );

    \I__10035\ : Span4Mux_v
    port map (
            O => \N__50100\,
            I => \N__50071\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__50095\,
            I => \N__50071\
        );

    \I__10033\ : Span4Mux_h
    port map (
            O => \N__50090\,
            I => \N__50066\
        );

    \I__10032\ : Span4Mux_v
    port map (
            O => \N__50087\,
            I => \N__50066\
        );

    \I__10031\ : Odrv12
    port map (
            O => \N__50084\,
            I => \r_SM_Main_1\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__50079\,
            I => \r_SM_Main_1\
        );

    \I__10029\ : Odrv12
    port map (
            O => \N__50076\,
            I => \r_SM_Main_1\
        );

    \I__10028\ : Odrv4
    port map (
            O => \N__50071\,
            I => \r_SM_Main_1\
        );

    \I__10027\ : Odrv4
    port map (
            O => \N__50066\,
            I => \r_SM_Main_1\
        );

    \I__10026\ : InMux
    port map (
            O => \N__50055\,
            I => \N__50052\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__50052\,
            I => \N__50049\
        );

    \I__10024\ : Span4Mux_s0_v
    port map (
            O => \N__50049\,
            I => \N__50045\
        );

    \I__10023\ : InMux
    port map (
            O => \N__50048\,
            I => \N__50039\
        );

    \I__10022\ : Sp12to4
    port map (
            O => \N__50045\,
            I => \N__50036\
        );

    \I__10021\ : InMux
    port map (
            O => \N__50044\,
            I => \N__50031\
        );

    \I__10020\ : InMux
    port map (
            O => \N__50043\,
            I => \N__50026\
        );

    \I__10019\ : InMux
    port map (
            O => \N__50042\,
            I => \N__50026\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__50039\,
            I => \N__50022\
        );

    \I__10017\ : Span12Mux_s4_v
    port map (
            O => \N__50036\,
            I => \N__50019\
        );

    \I__10016\ : InMux
    port map (
            O => \N__50035\,
            I => \N__50016\
        );

    \I__10015\ : InMux
    port map (
            O => \N__50034\,
            I => \N__50013\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__50031\,
            I => \N__50010\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__50026\,
            I => \N__50007\
        );

    \I__10012\ : InMux
    port map (
            O => \N__50025\,
            I => \N__50004\
        );

    \I__10011\ : Span4Mux_v
    port map (
            O => \N__50022\,
            I => \N__50001\
        );

    \I__10010\ : Span12Mux_h
    port map (
            O => \N__50019\,
            I => \N__49997\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__50016\,
            I => \N__49992\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__50013\,
            I => \N__49992\
        );

    \I__10007\ : Span4Mux_h
    port map (
            O => \N__50010\,
            I => \N__49985\
        );

    \I__10006\ : Span4Mux_v
    port map (
            O => \N__50007\,
            I => \N__49985\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__50004\,
            I => \N__49985\
        );

    \I__10004\ : Span4Mux_h
    port map (
            O => \N__50001\,
            I => \N__49982\
        );

    \I__10003\ : InMux
    port map (
            O => \N__50000\,
            I => \N__49979\
        );

    \I__10002\ : Span12Mux_v
    port map (
            O => \N__49997\,
            I => \N__49974\
        );

    \I__10001\ : Span12Mux_h
    port map (
            O => \N__49992\,
            I => \N__49974\
        );

    \I__10000\ : Span4Mux_h
    port map (
            O => \N__49985\,
            I => \N__49971\
        );

    \I__9999\ : Odrv4
    port map (
            O => \N__49982\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__49979\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__9997\ : Odrv12
    port map (
            O => \N__49974\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__9996\ : Odrv4
    port map (
            O => \N__49971\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__9995\ : InMux
    port map (
            O => \N__49962\,
            I => \N__49959\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__49959\,
            I => \N__49953\
        );

    \I__9993\ : InMux
    port map (
            O => \N__49958\,
            I => \N__49948\
        );

    \I__9992\ : InMux
    port map (
            O => \N__49957\,
            I => \N__49948\
        );

    \I__9991\ : InMux
    port map (
            O => \N__49956\,
            I => \N__49945\
        );

    \I__9990\ : Span4Mux_h
    port map (
            O => \N__49953\,
            I => \N__49935\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__49948\,
            I => \N__49935\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__49945\,
            I => \N__49932\
        );

    \I__9987\ : InMux
    port map (
            O => \N__49944\,
            I => \N__49929\
        );

    \I__9986\ : InMux
    port map (
            O => \N__49943\,
            I => \N__49924\
        );

    \I__9985\ : InMux
    port map (
            O => \N__49942\,
            I => \N__49924\
        );

    \I__9984\ : InMux
    port map (
            O => \N__49941\,
            I => \N__49921\
        );

    \I__9983\ : InMux
    port map (
            O => \N__49940\,
            I => \N__49918\
        );

    \I__9982\ : Span4Mux_h
    port map (
            O => \N__49935\,
            I => \N__49915\
        );

    \I__9981\ : Span4Mux_h
    port map (
            O => \N__49932\,
            I => \N__49910\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__49929\,
            I => \N__49910\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__49924\,
            I => \N__49907\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__49921\,
            I => \N__49904\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__49918\,
            I => \N__49901\
        );

    \I__9976\ : Sp12to4
    port map (
            O => \N__49915\,
            I => \N__49896\
        );

    \I__9975\ : Sp12to4
    port map (
            O => \N__49910\,
            I => \N__49896\
        );

    \I__9974\ : Span12Mux_s8_v
    port map (
            O => \N__49907\,
            I => \N__49893\
        );

    \I__9973\ : Span12Mux_s9_h
    port map (
            O => \N__49904\,
            I => \N__49886\
        );

    \I__9972\ : Span12Mux_h
    port map (
            O => \N__49901\,
            I => \N__49886\
        );

    \I__9971\ : Span12Mux_v
    port map (
            O => \N__49896\,
            I => \N__49886\
        );

    \I__9970\ : Odrv12
    port map (
            O => \N__49893\,
            I => \r_SM_Main_2\
        );

    \I__9969\ : Odrv12
    port map (
            O => \N__49886\,
            I => \r_SM_Main_2\
        );

    \I__9968\ : SRMux
    port map (
            O => \N__49881\,
            I => \N__49878\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__49878\,
            I => \N__49875\
        );

    \I__9966\ : Span4Mux_h
    port map (
            O => \N__49875\,
            I => \N__49872\
        );

    \I__9965\ : Sp12to4
    port map (
            O => \N__49872\,
            I => \N__49869\
        );

    \I__9964\ : Span12Mux_v
    port map (
            O => \N__49869\,
            I => \N__49866\
        );

    \I__9963\ : Odrv12
    port map (
            O => \N__49866\,
            I => \c0.rx.n22094\
        );

    \I__9962\ : InMux
    port map (
            O => \N__49863\,
            I => \N__49860\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__49860\,
            I => \c0.n46_adj_4739\
        );

    \I__9960\ : InMux
    port map (
            O => \N__49857\,
            I => \N__49854\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__49854\,
            I => \N__49851\
        );

    \I__9958\ : Span4Mux_v
    port map (
            O => \N__49851\,
            I => \N__49848\
        );

    \I__9957\ : Odrv4
    port map (
            O => \N__49848\,
            I => \c0.n39_adj_4295\
        );

    \I__9956\ : InMux
    port map (
            O => \N__49845\,
            I => \N__49841\
        );

    \I__9955\ : InMux
    port map (
            O => \N__49844\,
            I => \N__49838\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__49841\,
            I => \N__49833\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__49838\,
            I => \N__49833\
        );

    \I__9952\ : Odrv4
    port map (
            O => \N__49833\,
            I => \c0.n13043\
        );

    \I__9951\ : InMux
    port map (
            O => \N__49830\,
            I => \N__49824\
        );

    \I__9950\ : InMux
    port map (
            O => \N__49829\,
            I => \N__49821\
        );

    \I__9949\ : InMux
    port map (
            O => \N__49828\,
            I => \N__49818\
        );

    \I__9948\ : InMux
    port map (
            O => \N__49827\,
            I => \N__49815\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__49824\,
            I => \N__49812\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__49821\,
            I => \N__49809\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__49818\,
            I => \N__49806\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__49815\,
            I => \N__49799\
        );

    \I__9943\ : Span4Mux_v
    port map (
            O => \N__49812\,
            I => \N__49799\
        );

    \I__9942\ : Span4Mux_v
    port map (
            O => \N__49809\,
            I => \N__49799\
        );

    \I__9941\ : Odrv4
    port map (
            O => \N__49806\,
            I => \c0.n23912\
        );

    \I__9940\ : Odrv4
    port map (
            O => \N__49799\,
            I => \c0.n23912\
        );

    \I__9939\ : InMux
    port map (
            O => \N__49794\,
            I => \N__49788\
        );

    \I__9938\ : InMux
    port map (
            O => \N__49793\,
            I => \N__49788\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__49788\,
            I => \N__49783\
        );

    \I__9936\ : InMux
    port map (
            O => \N__49787\,
            I => \N__49780\
        );

    \I__9935\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49777\
        );

    \I__9934\ : Span4Mux_v
    port map (
            O => \N__49783\,
            I => \N__49774\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__49780\,
            I => \N__49771\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__49777\,
            I => \N__49768\
        );

    \I__9931\ : Span4Mux_h
    port map (
            O => \N__49774\,
            I => \N__49765\
        );

    \I__9930\ : Span4Mux_v
    port map (
            O => \N__49771\,
            I => \N__49762\
        );

    \I__9929\ : Odrv4
    port map (
            O => \N__49768\,
            I => \c0.n35\
        );

    \I__9928\ : Odrv4
    port map (
            O => \N__49765\,
            I => \c0.n35\
        );

    \I__9927\ : Odrv4
    port map (
            O => \N__49762\,
            I => \c0.n35\
        );

    \I__9926\ : CascadeMux
    port map (
            O => \N__49755\,
            I => \N__49752\
        );

    \I__9925\ : InMux
    port map (
            O => \N__49752\,
            I => \N__49749\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__49749\,
            I => \N__49746\
        );

    \I__9923\ : Span4Mux_h
    port map (
            O => \N__49746\,
            I => \N__49743\
        );

    \I__9922\ : Odrv4
    port map (
            O => \N__49743\,
            I => \c0.n22885\
        );

    \I__9921\ : InMux
    port map (
            O => \N__49740\,
            I => \N__49737\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__49737\,
            I => \N__49734\
        );

    \I__9919\ : Span4Mux_s1_v
    port map (
            O => \N__49734\,
            I => \N__49731\
        );

    \I__9918\ : Span4Mux_v
    port map (
            O => \N__49731\,
            I => \N__49727\
        );

    \I__9917\ : CascadeMux
    port map (
            O => \N__49730\,
            I => \N__49724\
        );

    \I__9916\ : Span4Mux_v
    port map (
            O => \N__49727\,
            I => \N__49719\
        );

    \I__9915\ : InMux
    port map (
            O => \N__49724\,
            I => \N__49713\
        );

    \I__9914\ : InMux
    port map (
            O => \N__49723\,
            I => \N__49713\
        );

    \I__9913\ : InMux
    port map (
            O => \N__49722\,
            I => \N__49710\
        );

    \I__9912\ : Span4Mux_v
    port map (
            O => \N__49719\,
            I => \N__49707\
        );

    \I__9911\ : InMux
    port map (
            O => \N__49718\,
            I => \N__49704\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__49713\,
            I => \N__49701\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__49710\,
            I => \N__49698\
        );

    \I__9908\ : Span4Mux_v
    port map (
            O => \N__49707\,
            I => \N__49693\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__49704\,
            I => \N__49693\
        );

    \I__9906\ : Span4Mux_v
    port map (
            O => \N__49701\,
            I => \N__49686\
        );

    \I__9905\ : Span4Mux_v
    port map (
            O => \N__49698\,
            I => \N__49686\
        );

    \I__9904\ : Span4Mux_h
    port map (
            O => \N__49693\,
            I => \N__49686\
        );

    \I__9903\ : Span4Mux_h
    port map (
            O => \N__49686\,
            I => \N__49681\
        );

    \I__9902\ : InMux
    port map (
            O => \N__49685\,
            I => \N__49678\
        );

    \I__9901\ : InMux
    port map (
            O => \N__49684\,
            I => \N__49675\
        );

    \I__9900\ : Span4Mux_h
    port map (
            O => \N__49681\,
            I => \N__49672\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__49678\,
            I => \N__49669\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__49675\,
            I => \r_Bit_Index_2\
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__49672\,
            I => \r_Bit_Index_2\
        );

    \I__9896\ : Odrv4
    port map (
            O => \N__49669\,
            I => \r_Bit_Index_2\
        );

    \I__9895\ : InMux
    port map (
            O => \N__49662\,
            I => \N__49659\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__49659\,
            I => \N__49653\
        );

    \I__9893\ : InMux
    port map (
            O => \N__49658\,
            I => \N__49650\
        );

    \I__9892\ : InMux
    port map (
            O => \N__49657\,
            I => \N__49645\
        );

    \I__9891\ : InMux
    port map (
            O => \N__49656\,
            I => \N__49642\
        );

    \I__9890\ : Span4Mux_s1_v
    port map (
            O => \N__49653\,
            I => \N__49639\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__49650\,
            I => \N__49635\
        );

    \I__9888\ : InMux
    port map (
            O => \N__49649\,
            I => \N__49629\
        );

    \I__9887\ : InMux
    port map (
            O => \N__49648\,
            I => \N__49629\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__49645\,
            I => \N__49626\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__49642\,
            I => \N__49623\
        );

    \I__9884\ : Sp12to4
    port map (
            O => \N__49639\,
            I => \N__49620\
        );

    \I__9883\ : CascadeMux
    port map (
            O => \N__49638\,
            I => \N__49617\
        );

    \I__9882\ : Span4Mux_v
    port map (
            O => \N__49635\,
            I => \N__49614\
        );

    \I__9881\ : InMux
    port map (
            O => \N__49634\,
            I => \N__49611\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__49629\,
            I => \N__49608\
        );

    \I__9879\ : Span4Mux_h
    port map (
            O => \N__49626\,
            I => \N__49603\
        );

    \I__9878\ : Span4Mux_h
    port map (
            O => \N__49623\,
            I => \N__49603\
        );

    \I__9877\ : Span12Mux_h
    port map (
            O => \N__49620\,
            I => \N__49600\
        );

    \I__9876\ : InMux
    port map (
            O => \N__49617\,
            I => \N__49597\
        );

    \I__9875\ : Span4Mux_h
    port map (
            O => \N__49614\,
            I => \N__49592\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__49611\,
            I => \N__49592\
        );

    \I__9873\ : Span4Mux_h
    port map (
            O => \N__49608\,
            I => \N__49589\
        );

    \I__9872\ : Span4Mux_h
    port map (
            O => \N__49603\,
            I => \N__49586\
        );

    \I__9871\ : Span12Mux_v
    port map (
            O => \N__49600\,
            I => \N__49583\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__49597\,
            I => \r_Bit_Index_1\
        );

    \I__9869\ : Odrv4
    port map (
            O => \N__49592\,
            I => \r_Bit_Index_1\
        );

    \I__9868\ : Odrv4
    port map (
            O => \N__49589\,
            I => \r_Bit_Index_1\
        );

    \I__9867\ : Odrv4
    port map (
            O => \N__49586\,
            I => \r_Bit_Index_1\
        );

    \I__9866\ : Odrv12
    port map (
            O => \N__49583\,
            I => \r_Bit_Index_1\
        );

    \I__9865\ : InMux
    port map (
            O => \N__49572\,
            I => \N__49569\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__49569\,
            I => \N__49566\
        );

    \I__9863\ : Span12Mux_h
    port map (
            O => \N__49566\,
            I => \N__49563\
        );

    \I__9862\ : Span12Mux_v
    port map (
            O => \N__49563\,
            I => \N__49560\
        );

    \I__9861\ : Odrv12
    port map (
            O => \N__49560\,
            I => n4
        );

    \I__9860\ : CascadeMux
    port map (
            O => \N__49557\,
            I => \c0.n20793_cascade_\
        );

    \I__9859\ : InMux
    port map (
            O => \N__49554\,
            I => \N__49545\
        );

    \I__9858\ : InMux
    port map (
            O => \N__49553\,
            I => \N__49545\
        );

    \I__9857\ : InMux
    port map (
            O => \N__49552\,
            I => \N__49545\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__49545\,
            I => \N__49542\
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__49542\,
            I => \c0.n12927\
        );

    \I__9854\ : CascadeMux
    port map (
            O => \N__49539\,
            I => \c0.n52_cascade_\
        );

    \I__9853\ : CascadeMux
    port map (
            O => \N__49536\,
            I => \c0.n47_adj_4537_cascade_\
        );

    \I__9852\ : InMux
    port map (
            O => \N__49533\,
            I => \N__49530\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__49530\,
            I => \N__49527\
        );

    \I__9850\ : Odrv4
    port map (
            O => \N__49527\,
            I => \c0.n24581\
        );

    \I__9849\ : CascadeMux
    port map (
            O => \N__49524\,
            I => \N__49520\
        );

    \I__9848\ : CascadeMux
    port map (
            O => \N__49523\,
            I => \N__49517\
        );

    \I__9847\ : InMux
    port map (
            O => \N__49520\,
            I => \N__49512\
        );

    \I__9846\ : InMux
    port map (
            O => \N__49517\,
            I => \N__49512\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__49512\,
            I => \c0.data_in_frame_29_1\
        );

    \I__9844\ : InMux
    port map (
            O => \N__49509\,
            I => \N__49503\
        );

    \I__9843\ : InMux
    port map (
            O => \N__49508\,
            I => \N__49503\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__49503\,
            I => \c0.data_in_frame_29_6\
        );

    \I__9841\ : InMux
    port map (
            O => \N__49500\,
            I => \N__49497\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__49497\,
            I => \c0.n20793\
        );

    \I__9839\ : CascadeMux
    port map (
            O => \N__49494\,
            I => \N__49491\
        );

    \I__9838\ : InMux
    port map (
            O => \N__49491\,
            I => \N__49488\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__49488\,
            I => \N__49485\
        );

    \I__9836\ : Span4Mux_h
    port map (
            O => \N__49485\,
            I => \N__49482\
        );

    \I__9835\ : Sp12to4
    port map (
            O => \N__49482\,
            I => \N__49479\
        );

    \I__9834\ : Odrv12
    port map (
            O => \N__49479\,
            I => \c0.n5_adj_4302\
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__49476\,
            I => \c0.n12_adj_4348_cascade_\
        );

    \I__9832\ : InMux
    port map (
            O => \N__49473\,
            I => \N__49470\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__49470\,
            I => \c0.n8_adj_4526\
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__49467\,
            I => \c0.n8_adj_4526_cascade_\
        );

    \I__9829\ : InMux
    port map (
            O => \N__49464\,
            I => \N__49461\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__49461\,
            I => \c0.n9_adj_4536\
        );

    \I__9827\ : InMux
    port map (
            O => \N__49458\,
            I => \N__49455\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__49455\,
            I => \c0.n14_adj_4528\
        );

    \I__9825\ : InMux
    port map (
            O => \N__49452\,
            I => \N__49449\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__49449\,
            I => \c0.n14_adj_4576\
        );

    \I__9823\ : InMux
    port map (
            O => \N__49446\,
            I => \N__49442\
        );

    \I__9822\ : InMux
    port map (
            O => \N__49445\,
            I => \N__49439\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__49442\,
            I => \c0.data_in_frame_29_5\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__49439\,
            I => \c0.data_in_frame_29_5\
        );

    \I__9819\ : CascadeMux
    port map (
            O => \N__49434\,
            I => \c0.n24098_cascade_\
        );

    \I__9818\ : InMux
    port map (
            O => \N__49431\,
            I => \N__49428\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__49428\,
            I => \c0.n10_adj_4484\
        );

    \I__9816\ : InMux
    port map (
            O => \N__49425\,
            I => \N__49419\
        );

    \I__9815\ : InMux
    port map (
            O => \N__49424\,
            I => \N__49416\
        );

    \I__9814\ : InMux
    port map (
            O => \N__49423\,
            I => \N__49413\
        );

    \I__9813\ : InMux
    port map (
            O => \N__49422\,
            I => \N__49410\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__49419\,
            I => \N__49407\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__49416\,
            I => \N__49402\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__49413\,
            I => \N__49402\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__49410\,
            I => \N__49397\
        );

    \I__9808\ : Span4Mux_h
    port map (
            O => \N__49407\,
            I => \N__49397\
        );

    \I__9807\ : Span4Mux_v
    port map (
            O => \N__49402\,
            I => \N__49394\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__49397\,
            I => data_in_3_0
        );

    \I__9805\ : Odrv4
    port map (
            O => \N__49394\,
            I => data_in_3_0
        );

    \I__9804\ : InMux
    port map (
            O => \N__49389\,
            I => \N__49386\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__49386\,
            I => \N__49382\
        );

    \I__9802\ : InMux
    port map (
            O => \N__49385\,
            I => \N__49379\
        );

    \I__9801\ : Span4Mux_v
    port map (
            O => \N__49382\,
            I => \N__49373\
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__49379\,
            I => \N__49373\
        );

    \I__9799\ : InMux
    port map (
            O => \N__49378\,
            I => \N__49370\
        );

    \I__9798\ : Span4Mux_v
    port map (
            O => \N__49373\,
            I => \N__49366\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__49370\,
            I => \N__49363\
        );

    \I__9796\ : InMux
    port map (
            O => \N__49369\,
            I => \N__49360\
        );

    \I__9795\ : Span4Mux_v
    port map (
            O => \N__49366\,
            I => \N__49353\
        );

    \I__9794\ : Span4Mux_h
    port map (
            O => \N__49363\,
            I => \N__49353\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__49360\,
            I => \N__49353\
        );

    \I__9792\ : Odrv4
    port map (
            O => \N__49353\,
            I => n12981
        );

    \I__9791\ : InMux
    port map (
            O => \N__49350\,
            I => \N__49344\
        );

    \I__9790\ : InMux
    port map (
            O => \N__49349\,
            I => \N__49344\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__49344\,
            I => \N__49341\
        );

    \I__9788\ : Span4Mux_h
    port map (
            O => \N__49341\,
            I => \N__49338\
        );

    \I__9787\ : Span4Mux_h
    port map (
            O => \N__49338\,
            I => \N__49335\
        );

    \I__9786\ : Odrv4
    port map (
            O => \N__49335\,
            I => n4_adj_4762
        );

    \I__9785\ : InMux
    port map (
            O => \N__49332\,
            I => \N__49329\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__49329\,
            I => \N__49326\
        );

    \I__9783\ : Odrv4
    port map (
            O => \N__49326\,
            I => \c0.n22716\
        );

    \I__9782\ : CascadeMux
    port map (
            O => \N__49323\,
            I => \c0.n22716_cascade_\
        );

    \I__9781\ : InMux
    port map (
            O => \N__49320\,
            I => \N__49317\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__49317\,
            I => \c0.n8_adj_4248\
        );

    \I__9779\ : CascadeMux
    port map (
            O => \N__49314\,
            I => \N__49311\
        );

    \I__9778\ : InMux
    port map (
            O => \N__49311\,
            I => \N__49307\
        );

    \I__9777\ : InMux
    port map (
            O => \N__49310\,
            I => \N__49304\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__49307\,
            I => \N__49299\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__49304\,
            I => \N__49296\
        );

    \I__9774\ : InMux
    port map (
            O => \N__49303\,
            I => \N__49293\
        );

    \I__9773\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49290\
        );

    \I__9772\ : Span4Mux_h
    port map (
            O => \N__49299\,
            I => \N__49287\
        );

    \I__9771\ : Span4Mux_h
    port map (
            O => \N__49296\,
            I => \N__49284\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__49293\,
            I => \N__49281\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__49290\,
            I => data_in_3_1
        );

    \I__9768\ : Odrv4
    port map (
            O => \N__49287\,
            I => data_in_3_1
        );

    \I__9767\ : Odrv4
    port map (
            O => \N__49284\,
            I => data_in_3_1
        );

    \I__9766\ : Odrv12
    port map (
            O => \N__49281\,
            I => data_in_3_1
        );

    \I__9765\ : InMux
    port map (
            O => \N__49272\,
            I => \N__49269\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__49269\,
            I => \N__49265\
        );

    \I__9763\ : CascadeMux
    port map (
            O => \N__49268\,
            I => \N__49261\
        );

    \I__9762\ : Span4Mux_v
    port map (
            O => \N__49265\,
            I => \N__49257\
        );

    \I__9761\ : InMux
    port map (
            O => \N__49264\,
            I => \N__49254\
        );

    \I__9760\ : InMux
    port map (
            O => \N__49261\,
            I => \N__49249\
        );

    \I__9759\ : InMux
    port map (
            O => \N__49260\,
            I => \N__49249\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__49257\,
            I => data_in_1_2
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__49254\,
            I => data_in_1_2
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__49249\,
            I => data_in_1_2
        );

    \I__9755\ : InMux
    port map (
            O => \N__49242\,
            I => \N__49239\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__49239\,
            I => \N__49234\
        );

    \I__9753\ : InMux
    port map (
            O => \N__49238\,
            I => \N__49231\
        );

    \I__9752\ : InMux
    port map (
            O => \N__49237\,
            I => \N__49228\
        );

    \I__9751\ : Span4Mux_h
    port map (
            O => \N__49234\,
            I => \N__49225\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__49231\,
            I => \N__49222\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__49228\,
            I => data_in_0_2
        );

    \I__9748\ : Odrv4
    port map (
            O => \N__49225\,
            I => data_in_0_2
        );

    \I__9747\ : Odrv12
    port map (
            O => \N__49222\,
            I => data_in_0_2
        );

    \I__9746\ : CascadeMux
    port map (
            O => \N__49215\,
            I => \N__49212\
        );

    \I__9745\ : InMux
    port map (
            O => \N__49212\,
            I => \N__49209\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__49209\,
            I => \c0.n10_adj_4732\
        );

    \I__9743\ : CascadeMux
    port map (
            O => \N__49206\,
            I => \c0.n26_adj_4733_cascade_\
        );

    \I__9742\ : CascadeMux
    port map (
            O => \N__49203\,
            I => \c0.n20409_cascade_\
        );

    \I__9741\ : InMux
    port map (
            O => \N__49200\,
            I => \N__49197\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__49197\,
            I => \N__49193\
        );

    \I__9739\ : InMux
    port map (
            O => \N__49196\,
            I => \N__49190\
        );

    \I__9738\ : Span4Mux_h
    port map (
            O => \N__49193\,
            I => \N__49187\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__49190\,
            I => \N__49181\
        );

    \I__9736\ : Span4Mux_h
    port map (
            O => \N__49187\,
            I => \N__49181\
        );

    \I__9735\ : InMux
    port map (
            O => \N__49186\,
            I => \N__49178\
        );

    \I__9734\ : Span4Mux_v
    port map (
            O => \N__49181\,
            I => \N__49175\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__49178\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__9732\ : Odrv4
    port map (
            O => \N__49175\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__9731\ : SRMux
    port map (
            O => \N__49170\,
            I => \N__49167\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__49167\,
            I => \N__49164\
        );

    \I__9729\ : Span4Mux_h
    port map (
            O => \N__49164\,
            I => \N__49161\
        );

    \I__9728\ : Span4Mux_v
    port map (
            O => \N__49161\,
            I => \N__49158\
        );

    \I__9727\ : Odrv4
    port map (
            O => \N__49158\,
            I => \c0.n21629\
        );

    \I__9726\ : InMux
    port map (
            O => \N__49155\,
            I => \N__49152\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__49152\,
            I => \N__49149\
        );

    \I__9724\ : Span4Mux_h
    port map (
            O => \N__49149\,
            I => \N__49146\
        );

    \I__9723\ : Odrv4
    port map (
            O => \N__49146\,
            I => \c0.n25_adj_4723\
        );

    \I__9722\ : InMux
    port map (
            O => \N__49143\,
            I => \N__49140\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__49140\,
            I => \N__49136\
        );

    \I__9720\ : CascadeMux
    port map (
            O => \N__49139\,
            I => \N__49133\
        );

    \I__9719\ : Span4Mux_v
    port map (
            O => \N__49136\,
            I => \N__49130\
        );

    \I__9718\ : InMux
    port map (
            O => \N__49133\,
            I => \N__49126\
        );

    \I__9717\ : Span4Mux_h
    port map (
            O => \N__49130\,
            I => \N__49123\
        );

    \I__9716\ : InMux
    port map (
            O => \N__49129\,
            I => \N__49120\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__49126\,
            I => \N__49117\
        );

    \I__9714\ : Sp12to4
    port map (
            O => \N__49123\,
            I => \N__49114\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__49120\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__9712\ : Odrv4
    port map (
            O => \N__49117\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__9711\ : Odrv12
    port map (
            O => \N__49114\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__9710\ : InMux
    port map (
            O => \N__49107\,
            I => \N__49104\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__49104\,
            I => \N__49099\
        );

    \I__9708\ : InMux
    port map (
            O => \N__49103\,
            I => \N__49096\
        );

    \I__9707\ : InMux
    port map (
            O => \N__49102\,
            I => \N__49093\
        );

    \I__9706\ : Span12Mux_h
    port map (
            O => \N__49099\,
            I => \N__49090\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__49096\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__49093\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__9703\ : Odrv12
    port map (
            O => \N__49090\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__9702\ : CascadeMux
    port map (
            O => \N__49083\,
            I => \N__49080\
        );

    \I__9701\ : InMux
    port map (
            O => \N__49080\,
            I => \N__49077\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__49077\,
            I => \N__49074\
        );

    \I__9699\ : Span4Mux_v
    port map (
            O => \N__49074\,
            I => \N__49070\
        );

    \I__9698\ : InMux
    port map (
            O => \N__49073\,
            I => \N__49066\
        );

    \I__9697\ : Span4Mux_h
    port map (
            O => \N__49070\,
            I => \N__49063\
        );

    \I__9696\ : InMux
    port map (
            O => \N__49069\,
            I => \N__49060\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__49066\,
            I => \N__49057\
        );

    \I__9694\ : Sp12to4
    port map (
            O => \N__49063\,
            I => \N__49054\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__49060\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__9692\ : Odrv4
    port map (
            O => \N__49057\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__9691\ : Odrv12
    port map (
            O => \N__49054\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__9690\ : InMux
    port map (
            O => \N__49047\,
            I => \N__49044\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__49044\,
            I => \N__49040\
        );

    \I__9688\ : InMux
    port map (
            O => \N__49043\,
            I => \N__49037\
        );

    \I__9687\ : Span4Mux_v
    port map (
            O => \N__49040\,
            I => \N__49033\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__49037\,
            I => \N__49030\
        );

    \I__9685\ : InMux
    port map (
            O => \N__49036\,
            I => \N__49027\
        );

    \I__9684\ : Span4Mux_v
    port map (
            O => \N__49033\,
            I => \N__49024\
        );

    \I__9683\ : Sp12to4
    port map (
            O => \N__49030\,
            I => \N__49019\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__49027\,
            I => \N__49019\
        );

    \I__9681\ : Sp12to4
    port map (
            O => \N__49024\,
            I => \N__49014\
        );

    \I__9680\ : Span12Mux_v
    port map (
            O => \N__49019\,
            I => \N__49014\
        );

    \I__9679\ : Odrv12
    port map (
            O => \N__49014\,
            I => \c0.n22049\
        );

    \I__9678\ : InMux
    port map (
            O => \N__49011\,
            I => \N__49008\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__49008\,
            I => \N__49004\
        );

    \I__9676\ : InMux
    port map (
            O => \N__49007\,
            I => \N__49000\
        );

    \I__9675\ : Span4Mux_h
    port map (
            O => \N__49004\,
            I => \N__48996\
        );

    \I__9674\ : InMux
    port map (
            O => \N__49003\,
            I => \N__48993\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__49000\,
            I => \N__48981\
        );

    \I__9672\ : InMux
    port map (
            O => \N__48999\,
            I => \N__48975\
        );

    \I__9671\ : Span4Mux_v
    port map (
            O => \N__48996\,
            I => \N__48970\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__48993\,
            I => \N__48970\
        );

    \I__9669\ : InMux
    port map (
            O => \N__48992\,
            I => \N__48966\
        );

    \I__9668\ : InMux
    port map (
            O => \N__48991\,
            I => \N__48963\
        );

    \I__9667\ : InMux
    port map (
            O => \N__48990\,
            I => \N__48957\
        );

    \I__9666\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48954\
        );

    \I__9665\ : InMux
    port map (
            O => \N__48988\,
            I => \N__48951\
        );

    \I__9664\ : InMux
    port map (
            O => \N__48987\,
            I => \N__48948\
        );

    \I__9663\ : InMux
    port map (
            O => \N__48986\,
            I => \N__48945\
        );

    \I__9662\ : InMux
    port map (
            O => \N__48985\,
            I => \N__48942\
        );

    \I__9661\ : InMux
    port map (
            O => \N__48984\,
            I => \N__48938\
        );

    \I__9660\ : Span4Mux_v
    port map (
            O => \N__48981\,
            I => \N__48935\
        );

    \I__9659\ : InMux
    port map (
            O => \N__48980\,
            I => \N__48932\
        );

    \I__9658\ : InMux
    port map (
            O => \N__48979\,
            I => \N__48929\
        );

    \I__9657\ : InMux
    port map (
            O => \N__48978\,
            I => \N__48925\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__48975\,
            I => \N__48922\
        );

    \I__9655\ : Span4Mux_v
    port map (
            O => \N__48970\,
            I => \N__48919\
        );

    \I__9654\ : InMux
    port map (
            O => \N__48969\,
            I => \N__48916\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__48966\,
            I => \N__48911\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__48963\,
            I => \N__48911\
        );

    \I__9651\ : InMux
    port map (
            O => \N__48962\,
            I => \N__48908\
        );

    \I__9650\ : InMux
    port map (
            O => \N__48961\,
            I => \N__48905\
        );

    \I__9649\ : InMux
    port map (
            O => \N__48960\,
            I => \N__48902\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__48957\,
            I => \N__48889\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__48954\,
            I => \N__48889\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__48951\,
            I => \N__48889\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__48948\,
            I => \N__48889\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__48945\,
            I => \N__48889\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__48942\,
            I => \N__48889\
        );

    \I__9642\ : InMux
    port map (
            O => \N__48941\,
            I => \N__48886\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__48938\,
            I => \N__48883\
        );

    \I__9640\ : Span4Mux_h
    port map (
            O => \N__48935\,
            I => \N__48879\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__48932\,
            I => \N__48874\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__48929\,
            I => \N__48874\
        );

    \I__9637\ : InMux
    port map (
            O => \N__48928\,
            I => \N__48871\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__48925\,
            I => \N__48867\
        );

    \I__9635\ : Span4Mux_h
    port map (
            O => \N__48922\,
            I => \N__48860\
        );

    \I__9634\ : Span4Mux_h
    port map (
            O => \N__48919\,
            I => \N__48860\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__48916\,
            I => \N__48860\
        );

    \I__9632\ : Span4Mux_h
    port map (
            O => \N__48911\,
            I => \N__48853\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__48908\,
            I => \N__48853\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__48905\,
            I => \N__48853\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__48902\,
            I => \N__48850\
        );

    \I__9628\ : Span4Mux_v
    port map (
            O => \N__48889\,
            I => \N__48845\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__48886\,
            I => \N__48845\
        );

    \I__9626\ : Span12Mux_h
    port map (
            O => \N__48883\,
            I => \N__48842\
        );

    \I__9625\ : InMux
    port map (
            O => \N__48882\,
            I => \N__48839\
        );

    \I__9624\ : Span4Mux_h
    port map (
            O => \N__48879\,
            I => \N__48834\
        );

    \I__9623\ : Span4Mux_h
    port map (
            O => \N__48874\,
            I => \N__48829\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__48871\,
            I => \N__48829\
        );

    \I__9621\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48826\
        );

    \I__9620\ : Span12Mux_v
    port map (
            O => \N__48867\,
            I => \N__48821\
        );

    \I__9619\ : Span4Mux_v
    port map (
            O => \N__48860\,
            I => \N__48814\
        );

    \I__9618\ : Span4Mux_v
    port map (
            O => \N__48853\,
            I => \N__48814\
        );

    \I__9617\ : Span4Mux_v
    port map (
            O => \N__48850\,
            I => \N__48814\
        );

    \I__9616\ : Span4Mux_h
    port map (
            O => \N__48845\,
            I => \N__48811\
        );

    \I__9615\ : Span12Mux_v
    port map (
            O => \N__48842\,
            I => \N__48806\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__48839\,
            I => \N__48806\
        );

    \I__9613\ : InMux
    port map (
            O => \N__48838\,
            I => \N__48803\
        );

    \I__9612\ : InMux
    port map (
            O => \N__48837\,
            I => \N__48800\
        );

    \I__9611\ : Span4Mux_v
    port map (
            O => \N__48834\,
            I => \N__48793\
        );

    \I__9610\ : Span4Mux_h
    port map (
            O => \N__48829\,
            I => \N__48793\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__48826\,
            I => \N__48793\
        );

    \I__9608\ : InMux
    port map (
            O => \N__48825\,
            I => \N__48790\
        );

    \I__9607\ : InMux
    port map (
            O => \N__48824\,
            I => \N__48787\
        );

    \I__9606\ : Odrv12
    port map (
            O => \N__48821\,
            I => \c0.n5\
        );

    \I__9605\ : Odrv4
    port map (
            O => \N__48814\,
            I => \c0.n5\
        );

    \I__9604\ : Odrv4
    port map (
            O => \N__48811\,
            I => \c0.n5\
        );

    \I__9603\ : Odrv12
    port map (
            O => \N__48806\,
            I => \c0.n5\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__48803\,
            I => \c0.n5\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__48800\,
            I => \c0.n5\
        );

    \I__9600\ : Odrv4
    port map (
            O => \N__48793\,
            I => \c0.n5\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__48790\,
            I => \c0.n5\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__48787\,
            I => \c0.n5\
        );

    \I__9597\ : InMux
    port map (
            O => \N__48768\,
            I => \N__48763\
        );

    \I__9596\ : InMux
    port map (
            O => \N__48767\,
            I => \N__48758\
        );

    \I__9595\ : InMux
    port map (
            O => \N__48766\,
            I => \N__48758\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__48763\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__48758\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__9592\ : SRMux
    port map (
            O => \N__48753\,
            I => \N__48750\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__48750\,
            I => \N__48747\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__48747\,
            I => \c0.n21647\
        );

    \I__9589\ : InMux
    port map (
            O => \N__48744\,
            I => \N__48740\
        );

    \I__9588\ : InMux
    port map (
            O => \N__48743\,
            I => \N__48736\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__48740\,
            I => \N__48733\
        );

    \I__9586\ : InMux
    port map (
            O => \N__48739\,
            I => \N__48728\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__48736\,
            I => \N__48723\
        );

    \I__9584\ : Span4Mux_v
    port map (
            O => \N__48733\,
            I => \N__48723\
        );

    \I__9583\ : InMux
    port map (
            O => \N__48732\,
            I => \N__48718\
        );

    \I__9582\ : InMux
    port map (
            O => \N__48731\,
            I => \N__48718\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__48728\,
            I => data_in_frame_5_6
        );

    \I__9580\ : Odrv4
    port map (
            O => \N__48723\,
            I => data_in_frame_5_6
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__48718\,
            I => data_in_frame_5_6
        );

    \I__9578\ : CascadeMux
    port map (
            O => \N__48711\,
            I => \N__48707\
        );

    \I__9577\ : InMux
    port map (
            O => \N__48710\,
            I => \N__48704\
        );

    \I__9576\ : InMux
    port map (
            O => \N__48707\,
            I => \N__48701\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__48704\,
            I => \N__48698\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__48701\,
            I => \N__48692\
        );

    \I__9573\ : Span4Mux_v
    port map (
            O => \N__48698\,
            I => \N__48692\
        );

    \I__9572\ : InMux
    port map (
            O => \N__48697\,
            I => \N__48689\
        );

    \I__9571\ : Odrv4
    port map (
            O => \N__48692\,
            I => \c0.data_in_frame_7_7\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__48689\,
            I => \c0.data_in_frame_7_7\
        );

    \I__9569\ : CascadeMux
    port map (
            O => \N__48684\,
            I => \N__48681\
        );

    \I__9568\ : InMux
    port map (
            O => \N__48681\,
            I => \N__48676\
        );

    \I__9567\ : InMux
    port map (
            O => \N__48680\,
            I => \N__48673\
        );

    \I__9566\ : InMux
    port map (
            O => \N__48679\,
            I => \N__48670\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__48676\,
            I => \N__48667\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__48673\,
            I => \N__48663\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__48670\,
            I => \N__48660\
        );

    \I__9562\ : Span4Mux_v
    port map (
            O => \N__48667\,
            I => \N__48657\
        );

    \I__9561\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48654\
        );

    \I__9560\ : Span12Mux_h
    port map (
            O => \N__48663\,
            I => \N__48651\
        );

    \I__9559\ : Span4Mux_v
    port map (
            O => \N__48660\,
            I => \N__48648\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__48657\,
            I => \N__48645\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__48654\,
            I => data_in_3_3
        );

    \I__9556\ : Odrv12
    port map (
            O => \N__48651\,
            I => data_in_3_3
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__48648\,
            I => data_in_3_3
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__48645\,
            I => data_in_3_3
        );

    \I__9553\ : InMux
    port map (
            O => \N__48636\,
            I => \N__48633\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__48633\,
            I => \N__48629\
        );

    \I__9551\ : InMux
    port map (
            O => \N__48632\,
            I => \N__48625\
        );

    \I__9550\ : Span4Mux_v
    port map (
            O => \N__48629\,
            I => \N__48622\
        );

    \I__9549\ : InMux
    port map (
            O => \N__48628\,
            I => \N__48619\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__48625\,
            I => \N__48616\
        );

    \I__9547\ : Span4Mux_h
    port map (
            O => \N__48622\,
            I => \N__48613\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__48619\,
            I => data_in_0_7
        );

    \I__9545\ : Odrv4
    port map (
            O => \N__48616\,
            I => data_in_0_7
        );

    \I__9544\ : Odrv4
    port map (
            O => \N__48613\,
            I => data_in_0_7
        );

    \I__9543\ : InMux
    port map (
            O => \N__48606\,
            I => \N__48603\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__48603\,
            I => \N__48600\
        );

    \I__9541\ : Span4Mux_v
    port map (
            O => \N__48600\,
            I => \N__48597\
        );

    \I__9540\ : Odrv4
    port map (
            O => \N__48597\,
            I => \c0.n14\
        );

    \I__9539\ : InMux
    port map (
            O => \N__48594\,
            I => \N__48591\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__48591\,
            I => \c0.n20_adj_4729\
        );

    \I__9537\ : CascadeMux
    port map (
            O => \N__48588\,
            I => \N__48585\
        );

    \I__9536\ : InMux
    port map (
            O => \N__48585\,
            I => \N__48582\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__48582\,
            I => \c0.n6_adj_4704\
        );

    \I__9534\ : CascadeMux
    port map (
            O => \N__48579\,
            I => \c0.n14016_cascade_\
        );

    \I__9533\ : CascadeMux
    port map (
            O => \N__48576\,
            I => \c0.n20_cascade_\
        );

    \I__9532\ : CascadeMux
    port map (
            O => \N__48573\,
            I => \c0.n6_adj_4254_cascade_\
        );

    \I__9531\ : InMux
    port map (
            O => \N__48570\,
            I => \N__48567\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__48567\,
            I => \N__48564\
        );

    \I__9529\ : Span4Mux_h
    port map (
            O => \N__48564\,
            I => \N__48561\
        );

    \I__9528\ : Odrv4
    port map (
            O => \N__48561\,
            I => \c0.n28_adj_4731\
        );

    \I__9527\ : CascadeMux
    port map (
            O => \N__48558\,
            I => \c0.n14_adj_4607_cascade_\
        );

    \I__9526\ : InMux
    port map (
            O => \N__48555\,
            I => \N__48549\
        );

    \I__9525\ : InMux
    port map (
            O => \N__48554\,
            I => \N__48549\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__48549\,
            I => \c0.n22626\
        );

    \I__9523\ : CascadeMux
    port map (
            O => \N__48546\,
            I => \c0.data_out_frame_0__7__N_2626_cascade_\
        );

    \I__9522\ : InMux
    port map (
            O => \N__48543\,
            I => \N__48537\
        );

    \I__9521\ : InMux
    port map (
            O => \N__48542\,
            I => \N__48537\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__48537\,
            I => \c0.n30_adj_4585\
        );

    \I__9519\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48531\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__48531\,
            I => \c0.n20_adj_4642\
        );

    \I__9517\ : CascadeMux
    port map (
            O => \N__48528\,
            I => \N__48525\
        );

    \I__9516\ : InMux
    port map (
            O => \N__48525\,
            I => \N__48522\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__48522\,
            I => \c0.n4_adj_4266\
        );

    \I__9514\ : CascadeMux
    port map (
            O => \N__48519\,
            I => \N__48516\
        );

    \I__9513\ : InMux
    port map (
            O => \N__48516\,
            I => \N__48512\
        );

    \I__9512\ : CascadeMux
    port map (
            O => \N__48515\,
            I => \N__48507\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__48512\,
            I => \N__48504\
        );

    \I__9510\ : InMux
    port map (
            O => \N__48511\,
            I => \N__48501\
        );

    \I__9509\ : InMux
    port map (
            O => \N__48510\,
            I => \N__48496\
        );

    \I__9508\ : InMux
    port map (
            O => \N__48507\,
            I => \N__48496\
        );

    \I__9507\ : Span4Mux_v
    port map (
            O => \N__48504\,
            I => \N__48493\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__48501\,
            I => \N__48486\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__48496\,
            I => \N__48486\
        );

    \I__9504\ : Sp12to4
    port map (
            O => \N__48493\,
            I => \N__48486\
        );

    \I__9503\ : Odrv12
    port map (
            O => \N__48486\,
            I => \c0.n5024\
        );

    \I__9502\ : InMux
    port map (
            O => \N__48483\,
            I => \N__48479\
        );

    \I__9501\ : InMux
    port map (
            O => \N__48482\,
            I => \N__48476\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__48479\,
            I => \N__48472\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__48476\,
            I => \N__48469\
        );

    \I__9498\ : InMux
    port map (
            O => \N__48475\,
            I => \N__48466\
        );

    \I__9497\ : Span4Mux_v
    port map (
            O => \N__48472\,
            I => \N__48463\
        );

    \I__9496\ : Span4Mux_h
    port map (
            O => \N__48469\,
            I => \N__48460\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__48466\,
            I => \N__48457\
        );

    \I__9494\ : Odrv4
    port map (
            O => \N__48463\,
            I => \c0.n12992\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__48460\,
            I => \c0.n12992\
        );

    \I__9492\ : Odrv12
    port map (
            O => \N__48457\,
            I => \c0.n12992\
        );

    \I__9491\ : InMux
    port map (
            O => \N__48450\,
            I => \N__48447\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__48447\,
            I => \N__48444\
        );

    \I__9489\ : Span4Mux_h
    port map (
            O => \N__48444\,
            I => \N__48440\
        );

    \I__9488\ : InMux
    port map (
            O => \N__48443\,
            I => \N__48437\
        );

    \I__9487\ : Odrv4
    port map (
            O => \N__48440\,
            I => \c0.n13052\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__48437\,
            I => \c0.n13052\
        );

    \I__9485\ : CascadeMux
    port map (
            O => \N__48432\,
            I => \N__48429\
        );

    \I__9484\ : InMux
    port map (
            O => \N__48429\,
            I => \N__48426\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__48426\,
            I => \N__48423\
        );

    \I__9482\ : Odrv4
    port map (
            O => \N__48423\,
            I => \c0.n24736\
        );

    \I__9481\ : InMux
    port map (
            O => \N__48420\,
            I => \N__48417\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__48417\,
            I => \N__48413\
        );

    \I__9479\ : InMux
    port map (
            O => \N__48416\,
            I => \N__48409\
        );

    \I__9478\ : Span4Mux_v
    port map (
            O => \N__48413\,
            I => \N__48406\
        );

    \I__9477\ : InMux
    port map (
            O => \N__48412\,
            I => \N__48403\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__48409\,
            I => \N__48400\
        );

    \I__9475\ : Span4Mux_h
    port map (
            O => \N__48406\,
            I => \N__48397\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__48403\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__9473\ : Odrv4
    port map (
            O => \N__48400\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__9472\ : Odrv4
    port map (
            O => \N__48397\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__9471\ : SRMux
    port map (
            O => \N__48390\,
            I => \N__48387\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__48387\,
            I => \N__48384\
        );

    \I__9469\ : Odrv4
    port map (
            O => \N__48384\,
            I => \c0.n21651\
        );

    \I__9468\ : CascadeMux
    port map (
            O => \N__48381\,
            I => \N__48369\
        );

    \I__9467\ : CascadeMux
    port map (
            O => \N__48380\,
            I => \N__48366\
        );

    \I__9466\ : InMux
    port map (
            O => \N__48379\,
            I => \N__48359\
        );

    \I__9465\ : CascadeMux
    port map (
            O => \N__48378\,
            I => \N__48356\
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__48377\,
            I => \N__48353\
        );

    \I__9463\ : InMux
    port map (
            O => \N__48376\,
            I => \N__48350\
        );

    \I__9462\ : InMux
    port map (
            O => \N__48375\,
            I => \N__48338\
        );

    \I__9461\ : InMux
    port map (
            O => \N__48374\,
            I => \N__48338\
        );

    \I__9460\ : InMux
    port map (
            O => \N__48373\,
            I => \N__48338\
        );

    \I__9459\ : InMux
    port map (
            O => \N__48372\,
            I => \N__48335\
        );

    \I__9458\ : InMux
    port map (
            O => \N__48369\,
            I => \N__48330\
        );

    \I__9457\ : InMux
    port map (
            O => \N__48366\,
            I => \N__48330\
        );

    \I__9456\ : InMux
    port map (
            O => \N__48365\,
            I => \N__48325\
        );

    \I__9455\ : InMux
    port map (
            O => \N__48364\,
            I => \N__48325\
        );

    \I__9454\ : InMux
    port map (
            O => \N__48363\,
            I => \N__48316\
        );

    \I__9453\ : InMux
    port map (
            O => \N__48362\,
            I => \N__48313\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__48359\,
            I => \N__48310\
        );

    \I__9451\ : InMux
    port map (
            O => \N__48356\,
            I => \N__48305\
        );

    \I__9450\ : InMux
    port map (
            O => \N__48353\,
            I => \N__48305\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__48350\,
            I => \N__48302\
        );

    \I__9448\ : InMux
    port map (
            O => \N__48349\,
            I => \N__48295\
        );

    \I__9447\ : InMux
    port map (
            O => \N__48348\,
            I => \N__48295\
        );

    \I__9446\ : InMux
    port map (
            O => \N__48347\,
            I => \N__48295\
        );

    \I__9445\ : InMux
    port map (
            O => \N__48346\,
            I => \N__48288\
        );

    \I__9444\ : InMux
    port map (
            O => \N__48345\,
            I => \N__48288\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__48338\,
            I => \N__48283\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__48335\,
            I => \N__48283\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__48330\,
            I => \N__48278\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__48325\,
            I => \N__48278\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__48324\,
            I => \N__48275\
        );

    \I__9438\ : CascadeMux
    port map (
            O => \N__48323\,
            I => \N__48272\
        );

    \I__9437\ : InMux
    port map (
            O => \N__48322\,
            I => \N__48260\
        );

    \I__9436\ : InMux
    port map (
            O => \N__48321\,
            I => \N__48260\
        );

    \I__9435\ : InMux
    port map (
            O => \N__48320\,
            I => \N__48260\
        );

    \I__9434\ : InMux
    port map (
            O => \N__48319\,
            I => \N__48260\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__48316\,
            I => \N__48257\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__48313\,
            I => \N__48227\
        );

    \I__9431\ : Span4Mux_h
    port map (
            O => \N__48310\,
            I => \N__48227\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__48305\,
            I => \N__48227\
        );

    \I__9429\ : Span4Mux_v
    port map (
            O => \N__48302\,
            I => \N__48227\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__48295\,
            I => \N__48227\
        );

    \I__9427\ : InMux
    port map (
            O => \N__48294\,
            I => \N__48222\
        );

    \I__9426\ : InMux
    port map (
            O => \N__48293\,
            I => \N__48222\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__48288\,
            I => \N__48215\
        );

    \I__9424\ : Span4Mux_v
    port map (
            O => \N__48283\,
            I => \N__48215\
        );

    \I__9423\ : Span4Mux_v
    port map (
            O => \N__48278\,
            I => \N__48215\
        );

    \I__9422\ : InMux
    port map (
            O => \N__48275\,
            I => \N__48210\
        );

    \I__9421\ : InMux
    port map (
            O => \N__48272\,
            I => \N__48210\
        );

    \I__9420\ : InMux
    port map (
            O => \N__48271\,
            I => \N__48197\
        );

    \I__9419\ : InMux
    port map (
            O => \N__48270\,
            I => \N__48194\
        );

    \I__9418\ : CascadeMux
    port map (
            O => \N__48269\,
            I => \N__48191\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__48260\,
            I => \N__48182\
        );

    \I__9416\ : Span4Mux_v
    port map (
            O => \N__48257\,
            I => \N__48179\
        );

    \I__9415\ : InMux
    port map (
            O => \N__48256\,
            I => \N__48176\
        );

    \I__9414\ : InMux
    port map (
            O => \N__48255\,
            I => \N__48169\
        );

    \I__9413\ : InMux
    port map (
            O => \N__48254\,
            I => \N__48169\
        );

    \I__9412\ : InMux
    port map (
            O => \N__48253\,
            I => \N__48169\
        );

    \I__9411\ : InMux
    port map (
            O => \N__48252\,
            I => \N__48162\
        );

    \I__9410\ : InMux
    port map (
            O => \N__48251\,
            I => \N__48162\
        );

    \I__9409\ : InMux
    port map (
            O => \N__48250\,
            I => \N__48162\
        );

    \I__9408\ : InMux
    port map (
            O => \N__48249\,
            I => \N__48159\
        );

    \I__9407\ : InMux
    port map (
            O => \N__48248\,
            I => \N__48154\
        );

    \I__9406\ : InMux
    port map (
            O => \N__48247\,
            I => \N__48154\
        );

    \I__9405\ : InMux
    port map (
            O => \N__48246\,
            I => \N__48143\
        );

    \I__9404\ : InMux
    port map (
            O => \N__48245\,
            I => \N__48143\
        );

    \I__9403\ : InMux
    port map (
            O => \N__48244\,
            I => \N__48143\
        );

    \I__9402\ : InMux
    port map (
            O => \N__48243\,
            I => \N__48143\
        );

    \I__9401\ : InMux
    port map (
            O => \N__48242\,
            I => \N__48143\
        );

    \I__9400\ : CascadeMux
    port map (
            O => \N__48241\,
            I => \N__48138\
        );

    \I__9399\ : CascadeMux
    port map (
            O => \N__48240\,
            I => \N__48135\
        );

    \I__9398\ : InMux
    port map (
            O => \N__48239\,
            I => \N__48126\
        );

    \I__9397\ : InMux
    port map (
            O => \N__48238\,
            I => \N__48126\
        );

    \I__9396\ : Span4Mux_v
    port map (
            O => \N__48227\,
            I => \N__48117\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__48222\,
            I => \N__48117\
        );

    \I__9394\ : Span4Mux_h
    port map (
            O => \N__48215\,
            I => \N__48117\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__48210\,
            I => \N__48117\
        );

    \I__9392\ : InMux
    port map (
            O => \N__48209\,
            I => \N__48108\
        );

    \I__9391\ : InMux
    port map (
            O => \N__48208\,
            I => \N__48108\
        );

    \I__9390\ : InMux
    port map (
            O => \N__48207\,
            I => \N__48108\
        );

    \I__9389\ : InMux
    port map (
            O => \N__48206\,
            I => \N__48108\
        );

    \I__9388\ : InMux
    port map (
            O => \N__48205\,
            I => \N__48099\
        );

    \I__9387\ : InMux
    port map (
            O => \N__48204\,
            I => \N__48099\
        );

    \I__9386\ : InMux
    port map (
            O => \N__48203\,
            I => \N__48099\
        );

    \I__9385\ : InMux
    port map (
            O => \N__48202\,
            I => \N__48099\
        );

    \I__9384\ : InMux
    port map (
            O => \N__48201\,
            I => \N__48094\
        );

    \I__9383\ : InMux
    port map (
            O => \N__48200\,
            I => \N__48094\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__48197\,
            I => \N__48091\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__48194\,
            I => \N__48088\
        );

    \I__9380\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48078\
        );

    \I__9379\ : InMux
    port map (
            O => \N__48190\,
            I => \N__48078\
        );

    \I__9378\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48078\
        );

    \I__9377\ : InMux
    port map (
            O => \N__48188\,
            I => \N__48072\
        );

    \I__9376\ : InMux
    port map (
            O => \N__48187\,
            I => \N__48072\
        );

    \I__9375\ : InMux
    port map (
            O => \N__48186\,
            I => \N__48069\
        );

    \I__9374\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48064\
        );

    \I__9373\ : Span4Mux_v
    port map (
            O => \N__48182\,
            I => \N__48047\
        );

    \I__9372\ : Span4Mux_h
    port map (
            O => \N__48179\,
            I => \N__48047\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__48176\,
            I => \N__48047\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__48169\,
            I => \N__48047\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__48162\,
            I => \N__48047\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__48159\,
            I => \N__48047\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__48154\,
            I => \N__48047\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__48143\,
            I => \N__48047\
        );

    \I__9365\ : InMux
    port map (
            O => \N__48142\,
            I => \N__48036\
        );

    \I__9364\ : InMux
    port map (
            O => \N__48141\,
            I => \N__48036\
        );

    \I__9363\ : InMux
    port map (
            O => \N__48138\,
            I => \N__48036\
        );

    \I__9362\ : InMux
    port map (
            O => \N__48135\,
            I => \N__48036\
        );

    \I__9361\ : InMux
    port map (
            O => \N__48134\,
            I => \N__48036\
        );

    \I__9360\ : InMux
    port map (
            O => \N__48133\,
            I => \N__48029\
        );

    \I__9359\ : InMux
    port map (
            O => \N__48132\,
            I => \N__48029\
        );

    \I__9358\ : InMux
    port map (
            O => \N__48131\,
            I => \N__48029\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__48126\,
            I => \N__48024\
        );

    \I__9356\ : Span4Mux_v
    port map (
            O => \N__48117\,
            I => \N__48024\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__48108\,
            I => \N__48013\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__48099\,
            I => \N__48013\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__48094\,
            I => \N__48013\
        );

    \I__9352\ : Span4Mux_h
    port map (
            O => \N__48091\,
            I => \N__48013\
        );

    \I__9351\ : Span4Mux_v
    port map (
            O => \N__48088\,
            I => \N__48013\
        );

    \I__9350\ : InMux
    port map (
            O => \N__48087\,
            I => \N__48006\
        );

    \I__9349\ : InMux
    port map (
            O => \N__48086\,
            I => \N__48006\
        );

    \I__9348\ : InMux
    port map (
            O => \N__48085\,
            I => \N__48006\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__48078\,
            I => \N__48003\
        );

    \I__9346\ : InMux
    port map (
            O => \N__48077\,
            I => \N__48000\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__48072\,
            I => \N__47995\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__48069\,
            I => \N__47995\
        );

    \I__9343\ : InMux
    port map (
            O => \N__48068\,
            I => \N__47991\
        );

    \I__9342\ : InMux
    port map (
            O => \N__48067\,
            I => \N__47988\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__48064\,
            I => \N__47983\
        );

    \I__9340\ : Span4Mux_v
    port map (
            O => \N__48047\,
            I => \N__47983\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__48036\,
            I => \N__47974\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__48029\,
            I => \N__47974\
        );

    \I__9337\ : Span4Mux_h
    port map (
            O => \N__48024\,
            I => \N__47974\
        );

    \I__9336\ : Span4Mux_v
    port map (
            O => \N__48013\,
            I => \N__47974\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__48006\,
            I => \N__47969\
        );

    \I__9334\ : Span4Mux_h
    port map (
            O => \N__48003\,
            I => \N__47969\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__48000\,
            I => \N__47964\
        );

    \I__9332\ : Span4Mux_v
    port map (
            O => \N__47995\,
            I => \N__47964\
        );

    \I__9331\ : InMux
    port map (
            O => \N__47994\,
            I => \N__47961\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__47991\,
            I => \N__47956\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__47988\,
            I => \N__47956\
        );

    \I__9328\ : Sp12to4
    port map (
            O => \N__47983\,
            I => \N__47953\
        );

    \I__9327\ : Span4Mux_v
    port map (
            O => \N__47974\,
            I => \N__47950\
        );

    \I__9326\ : Span4Mux_h
    port map (
            O => \N__47969\,
            I => \N__47947\
        );

    \I__9325\ : Sp12to4
    port map (
            O => \N__47964\,
            I => \N__47944\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__47961\,
            I => \N__47939\
        );

    \I__9323\ : Span12Mux_v
    port map (
            O => \N__47956\,
            I => \N__47939\
        );

    \I__9322\ : Span12Mux_h
    port map (
            O => \N__47953\,
            I => \N__47936\
        );

    \I__9321\ : Span4Mux_v
    port map (
            O => \N__47950\,
            I => \N__47933\
        );

    \I__9320\ : Span4Mux_v
    port map (
            O => \N__47947\,
            I => \N__47930\
        );

    \I__9319\ : Span12Mux_h
    port map (
            O => \N__47944\,
            I => \N__47927\
        );

    \I__9318\ : Span12Mux_v
    port map (
            O => \N__47939\,
            I => \N__47922\
        );

    \I__9317\ : Span12Mux_v
    port map (
            O => \N__47936\,
            I => \N__47922\
        );

    \I__9316\ : Span4Mux_v
    port map (
            O => \N__47933\,
            I => \N__47919\
        );

    \I__9315\ : Odrv4
    port map (
            O => \N__47930\,
            I => \FRAME_MATCHER_state_31_N_2975_2\
        );

    \I__9314\ : Odrv12
    port map (
            O => \N__47927\,
            I => \FRAME_MATCHER_state_31_N_2975_2\
        );

    \I__9313\ : Odrv12
    port map (
            O => \N__47922\,
            I => \FRAME_MATCHER_state_31_N_2975_2\
        );

    \I__9312\ : Odrv4
    port map (
            O => \N__47919\,
            I => \FRAME_MATCHER_state_31_N_2975_2\
        );

    \I__9311\ : CascadeMux
    port map (
            O => \N__47910\,
            I => \c0.n22_adj_4643_cascade_\
        );

    \I__9310\ : CascadeMux
    port map (
            O => \N__47907\,
            I => \c0.n10_adj_4639_cascade_\
        );

    \I__9309\ : InMux
    port map (
            O => \N__47904\,
            I => \N__47901\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__47901\,
            I => \c0.n13_adj_4640\
        );

    \I__9307\ : CascadeMux
    port map (
            O => \N__47898\,
            I => \c0.n22134_cascade_\
        );

    \I__9306\ : CascadeMux
    port map (
            O => \N__47895\,
            I => \N__47890\
        );

    \I__9305\ : InMux
    port map (
            O => \N__47894\,
            I => \N__47887\
        );

    \I__9304\ : InMux
    port map (
            O => \N__47893\,
            I => \N__47884\
        );

    \I__9303\ : InMux
    port map (
            O => \N__47890\,
            I => \N__47880\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__47887\,
            I => \N__47873\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__47884\,
            I => \N__47873\
        );

    \I__9300\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47870\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__47880\,
            I => \N__47867\
        );

    \I__9298\ : InMux
    port map (
            O => \N__47879\,
            I => \N__47862\
        );

    \I__9297\ : InMux
    port map (
            O => \N__47878\,
            I => \N__47862\
        );

    \I__9296\ : Span4Mux_h
    port map (
            O => \N__47873\,
            I => \N__47859\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__47870\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__9294\ : Odrv12
    port map (
            O => \N__47867\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__47862\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__9292\ : Odrv4
    port map (
            O => \N__47859\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__9291\ : SRMux
    port map (
            O => \N__47850\,
            I => \N__47847\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__47847\,
            I => \N__47844\
        );

    \I__9289\ : Odrv4
    port map (
            O => \N__47844\,
            I => \c0.n21633\
        );

    \I__9288\ : InMux
    port map (
            O => \N__47841\,
            I => \N__47838\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__47838\,
            I => \N__47833\
        );

    \I__9286\ : InMux
    port map (
            O => \N__47837\,
            I => \N__47830\
        );

    \I__9285\ : InMux
    port map (
            O => \N__47836\,
            I => \N__47824\
        );

    \I__9284\ : Span4Mux_v
    port map (
            O => \N__47833\,
            I => \N__47819\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__47830\,
            I => \N__47819\
        );

    \I__9282\ : InMux
    port map (
            O => \N__47829\,
            I => \N__47809\
        );

    \I__9281\ : InMux
    port map (
            O => \N__47828\,
            I => \N__47809\
        );

    \I__9280\ : InMux
    port map (
            O => \N__47827\,
            I => \N__47806\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__47824\,
            I => \N__47803\
        );

    \I__9278\ : Span4Mux_h
    port map (
            O => \N__47819\,
            I => \N__47800\
        );

    \I__9277\ : InMux
    port map (
            O => \N__47818\,
            I => \N__47791\
        );

    \I__9276\ : InMux
    port map (
            O => \N__47817\,
            I => \N__47791\
        );

    \I__9275\ : InMux
    port map (
            O => \N__47816\,
            I => \N__47791\
        );

    \I__9274\ : InMux
    port map (
            O => \N__47815\,
            I => \N__47791\
        );

    \I__9273\ : InMux
    port map (
            O => \N__47814\,
            I => \N__47784\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__47809\,
            I => \N__47781\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__47806\,
            I => \N__47778\
        );

    \I__9270\ : Span12Mux_v
    port map (
            O => \N__47803\,
            I => \N__47775\
        );

    \I__9269\ : Span4Mux_v
    port map (
            O => \N__47800\,
            I => \N__47770\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__47791\,
            I => \N__47770\
        );

    \I__9267\ : InMux
    port map (
            O => \N__47790\,
            I => \N__47763\
        );

    \I__9266\ : InMux
    port map (
            O => \N__47789\,
            I => \N__47763\
        );

    \I__9265\ : InMux
    port map (
            O => \N__47788\,
            I => \N__47763\
        );

    \I__9264\ : InMux
    port map (
            O => \N__47787\,
            I => \N__47760\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__47784\,
            I => \N__47757\
        );

    \I__9262\ : Span4Mux_h
    port map (
            O => \N__47781\,
            I => \N__47752\
        );

    \I__9261\ : Span4Mux_v
    port map (
            O => \N__47778\,
            I => \N__47752\
        );

    \I__9260\ : Odrv12
    port map (
            O => \N__47775\,
            I => \c0.n6\
        );

    \I__9259\ : Odrv4
    port map (
            O => \N__47770\,
            I => \c0.n6\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__47763\,
            I => \c0.n6\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__47760\,
            I => \c0.n6\
        );

    \I__9256\ : Odrv4
    port map (
            O => \N__47757\,
            I => \c0.n6\
        );

    \I__9255\ : Odrv4
    port map (
            O => \N__47752\,
            I => \c0.n6\
        );

    \I__9254\ : InMux
    port map (
            O => \N__47739\,
            I => \N__47736\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__47736\,
            I => \c0.n18_adj_4485\
        );

    \I__9252\ : CascadeMux
    port map (
            O => \N__47733\,
            I => \N__47717\
        );

    \I__9251\ : InMux
    port map (
            O => \N__47732\,
            I => \N__47712\
        );

    \I__9250\ : InMux
    port map (
            O => \N__47731\,
            I => \N__47700\
        );

    \I__9249\ : InMux
    port map (
            O => \N__47730\,
            I => \N__47700\
        );

    \I__9248\ : InMux
    port map (
            O => \N__47729\,
            I => \N__47700\
        );

    \I__9247\ : InMux
    port map (
            O => \N__47728\,
            I => \N__47700\
        );

    \I__9246\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47700\
        );

    \I__9245\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47697\
        );

    \I__9244\ : InMux
    port map (
            O => \N__47725\,
            I => \N__47691\
        );

    \I__9243\ : InMux
    port map (
            O => \N__47724\,
            I => \N__47691\
        );

    \I__9242\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47688\
        );

    \I__9241\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47683\
        );

    \I__9240\ : InMux
    port map (
            O => \N__47721\,
            I => \N__47683\
        );

    \I__9239\ : InMux
    port map (
            O => \N__47720\,
            I => \N__47680\
        );

    \I__9238\ : InMux
    port map (
            O => \N__47717\,
            I => \N__47673\
        );

    \I__9237\ : InMux
    port map (
            O => \N__47716\,
            I => \N__47673\
        );

    \I__9236\ : InMux
    port map (
            O => \N__47715\,
            I => \N__47673\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__47712\,
            I => \N__47670\
        );

    \I__9234\ : InMux
    port map (
            O => \N__47711\,
            I => \N__47667\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__47700\,
            I => \N__47662\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__47697\,
            I => \N__47662\
        );

    \I__9231\ : InMux
    port map (
            O => \N__47696\,
            I => \N__47659\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__47691\,
            I => \N__47649\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__47688\,
            I => \N__47642\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__47683\,
            I => \N__47642\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__47680\,
            I => \N__47637\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__47673\,
            I => \N__47637\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__47670\,
            I => \N__47628\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__47667\,
            I => \N__47628\
        );

    \I__9223\ : Span4Mux_v
    port map (
            O => \N__47662\,
            I => \N__47628\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__47659\,
            I => \N__47628\
        );

    \I__9221\ : InMux
    port map (
            O => \N__47658\,
            I => \N__47623\
        );

    \I__9220\ : InMux
    port map (
            O => \N__47657\,
            I => \N__47623\
        );

    \I__9219\ : InMux
    port map (
            O => \N__47656\,
            I => \N__47616\
        );

    \I__9218\ : InMux
    port map (
            O => \N__47655\,
            I => \N__47616\
        );

    \I__9217\ : InMux
    port map (
            O => \N__47654\,
            I => \N__47616\
        );

    \I__9216\ : InMux
    port map (
            O => \N__47653\,
            I => \N__47613\
        );

    \I__9215\ : CascadeMux
    port map (
            O => \N__47652\,
            I => \N__47607\
        );

    \I__9214\ : Span4Mux_v
    port map (
            O => \N__47649\,
            I => \N__47604\
        );

    \I__9213\ : InMux
    port map (
            O => \N__47648\,
            I => \N__47599\
        );

    \I__9212\ : InMux
    port map (
            O => \N__47647\,
            I => \N__47599\
        );

    \I__9211\ : Span4Mux_v
    port map (
            O => \N__47642\,
            I => \N__47594\
        );

    \I__9210\ : Span4Mux_h
    port map (
            O => \N__47637\,
            I => \N__47585\
        );

    \I__9209\ : Span4Mux_v
    port map (
            O => \N__47628\,
            I => \N__47585\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__47623\,
            I => \N__47585\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__47616\,
            I => \N__47585\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__47613\,
            I => \N__47582\
        );

    \I__9205\ : InMux
    port map (
            O => \N__47612\,
            I => \N__47579\
        );

    \I__9204\ : InMux
    port map (
            O => \N__47611\,
            I => \N__47576\
        );

    \I__9203\ : InMux
    port map (
            O => \N__47610\,
            I => \N__47571\
        );

    \I__9202\ : InMux
    port map (
            O => \N__47607\,
            I => \N__47571\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__47604\,
            I => \N__47566\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__47599\,
            I => \N__47566\
        );

    \I__9199\ : InMux
    port map (
            O => \N__47598\,
            I => \N__47563\
        );

    \I__9198\ : InMux
    port map (
            O => \N__47597\,
            I => \N__47560\
        );

    \I__9197\ : Sp12to4
    port map (
            O => \N__47594\,
            I => \N__47557\
        );

    \I__9196\ : Span4Mux_h
    port map (
            O => \N__47585\,
            I => \N__47554\
        );

    \I__9195\ : Span12Mux_v
    port map (
            O => \N__47582\,
            I => \N__47545\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__47579\,
            I => \N__47545\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__47576\,
            I => \N__47545\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__47571\,
            I => \N__47545\
        );

    \I__9191\ : Sp12to4
    port map (
            O => \N__47566\,
            I => \N__47538\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__47563\,
            I => \N__47538\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__47560\,
            I => \N__47538\
        );

    \I__9188\ : Span12Mux_h
    port map (
            O => \N__47557\,
            I => \N__47535\
        );

    \I__9187\ : Span4Mux_h
    port map (
            O => \N__47554\,
            I => \N__47532\
        );

    \I__9186\ : Span12Mux_h
    port map (
            O => \N__47545\,
            I => \N__47527\
        );

    \I__9185\ : Span12Mux_s11_v
    port map (
            O => \N__47538\,
            I => \N__47527\
        );

    \I__9184\ : Odrv12
    port map (
            O => \N__47535\,
            I => count_enable
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__47532\,
            I => count_enable
        );

    \I__9182\ : Odrv12
    port map (
            O => \N__47527\,
            I => count_enable
        );

    \I__9181\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47517\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__47517\,
            I => \N__47514\
        );

    \I__9179\ : Span4Mux_h
    port map (
            O => \N__47514\,
            I => \N__47511\
        );

    \I__9178\ : Span4Mux_v
    port map (
            O => \N__47511\,
            I => \N__47508\
        );

    \I__9177\ : Span4Mux_v
    port map (
            O => \N__47508\,
            I => \N__47505\
        );

    \I__9176\ : Odrv4
    port map (
            O => \N__47505\,
            I => n2343
        );

    \I__9175\ : CascadeMux
    port map (
            O => \N__47502\,
            I => \N__47498\
        );

    \I__9174\ : CascadeMux
    port map (
            O => \N__47501\,
            I => \N__47494\
        );

    \I__9173\ : InMux
    port map (
            O => \N__47498\,
            I => \N__47489\
        );

    \I__9172\ : InMux
    port map (
            O => \N__47497\,
            I => \N__47489\
        );

    \I__9171\ : InMux
    port map (
            O => \N__47494\,
            I => \N__47486\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__47489\,
            I => \N__47481\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__47486\,
            I => \N__47478\
        );

    \I__9168\ : InMux
    port map (
            O => \N__47485\,
            I => \N__47475\
        );

    \I__9167\ : InMux
    port map (
            O => \N__47484\,
            I => \N__47472\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__47481\,
            I => \N__47469\
        );

    \I__9165\ : Sp12to4
    port map (
            O => \N__47478\,
            I => \N__47465\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__47475\,
            I => \N__47462\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__47472\,
            I => \N__47457\
        );

    \I__9162\ : Span4Mux_v
    port map (
            O => \N__47469\,
            I => \N__47457\
        );

    \I__9161\ : InMux
    port map (
            O => \N__47468\,
            I => \N__47453\
        );

    \I__9160\ : Span12Mux_v
    port map (
            O => \N__47465\,
            I => \N__47450\
        );

    \I__9159\ : Span12Mux_h
    port map (
            O => \N__47462\,
            I => \N__47447\
        );

    \I__9158\ : Span4Mux_v
    port map (
            O => \N__47457\,
            I => \N__47444\
        );

    \I__9157\ : InMux
    port map (
            O => \N__47456\,
            I => \N__47441\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__47453\,
            I => encoder0_position_14
        );

    \I__9155\ : Odrv12
    port map (
            O => \N__47450\,
            I => encoder0_position_14
        );

    \I__9154\ : Odrv12
    port map (
            O => \N__47447\,
            I => encoder0_position_14
        );

    \I__9153\ : Odrv4
    port map (
            O => \N__47444\,
            I => encoder0_position_14
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__47441\,
            I => encoder0_position_14
        );

    \I__9151\ : InMux
    port map (
            O => \N__47430\,
            I => \N__47426\
        );

    \I__9150\ : InMux
    port map (
            O => \N__47429\,
            I => \N__47423\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__47426\,
            I => \N__47420\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__47423\,
            I => \N__47415\
        );

    \I__9147\ : Span4Mux_v
    port map (
            O => \N__47420\,
            I => \N__47415\
        );

    \I__9146\ : Span4Mux_h
    port map (
            O => \N__47415\,
            I => \N__47412\
        );

    \I__9145\ : Odrv4
    port map (
            O => \N__47412\,
            I => n4_adj_4761
        );

    \I__9144\ : CascadeMux
    port map (
            O => \N__47409\,
            I => \N__47405\
        );

    \I__9143\ : CascadeMux
    port map (
            O => \N__47408\,
            I => \N__47402\
        );

    \I__9142\ : InMux
    port map (
            O => \N__47405\,
            I => \N__47399\
        );

    \I__9141\ : InMux
    port map (
            O => \N__47402\,
            I => \N__47396\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__47399\,
            I => \N__47393\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__47396\,
            I => \c0.data_in_frame_29_3\
        );

    \I__9138\ : Odrv4
    port map (
            O => \N__47393\,
            I => \c0.data_in_frame_29_3\
        );

    \I__9137\ : InMux
    port map (
            O => \N__47388\,
            I => \N__47385\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__47385\,
            I => \N__47382\
        );

    \I__9135\ : Span4Mux_v
    port map (
            O => \N__47382\,
            I => \N__47379\
        );

    \I__9134\ : Odrv4
    port map (
            O => \N__47379\,
            I => \c0.n17_adj_4483\
        );

    \I__9133\ : CascadeMux
    port map (
            O => \N__47376\,
            I => \c0.n26_adj_4480_cascade_\
        );

    \I__9132\ : InMux
    port map (
            O => \N__47373\,
            I => \N__47370\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__47370\,
            I => \N__47367\
        );

    \I__9130\ : Span4Mux_h
    port map (
            O => \N__47367\,
            I => \N__47363\
        );

    \I__9129\ : InMux
    port map (
            O => \N__47366\,
            I => \N__47360\
        );

    \I__9128\ : Odrv4
    port map (
            O => \N__47363\,
            I => \c0.n63_adj_4249\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__47360\,
            I => \c0.n63_adj_4249\
        );

    \I__9126\ : CascadeMux
    port map (
            O => \N__47355\,
            I => \c0.n34_adj_4546_cascade_\
        );

    \I__9125\ : CascadeMux
    port map (
            O => \N__47352\,
            I => \N__47344\
        );

    \I__9124\ : InMux
    port map (
            O => \N__47351\,
            I => \N__47336\
        );

    \I__9123\ : InMux
    port map (
            O => \N__47350\,
            I => \N__47336\
        );

    \I__9122\ : InMux
    port map (
            O => \N__47349\,
            I => \N__47336\
        );

    \I__9121\ : InMux
    port map (
            O => \N__47348\,
            I => \N__47333\
        );

    \I__9120\ : InMux
    port map (
            O => \N__47347\,
            I => \N__47326\
        );

    \I__9119\ : InMux
    port map (
            O => \N__47344\,
            I => \N__47326\
        );

    \I__9118\ : InMux
    port map (
            O => \N__47343\,
            I => \N__47326\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__47336\,
            I => n24622
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__47333\,
            I => n24622
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__47326\,
            I => n24622
        );

    \I__9114\ : CascadeMux
    port map (
            O => \N__47319\,
            I => \n24622_cascade_\
        );

    \I__9113\ : CascadeMux
    port map (
            O => \N__47316\,
            I => \N__47313\
        );

    \I__9112\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47309\
        );

    \I__9111\ : InMux
    port map (
            O => \N__47312\,
            I => \N__47306\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__47309\,
            I => \N__47302\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__47306\,
            I => \N__47299\
        );

    \I__9108\ : CascadeMux
    port map (
            O => \N__47305\,
            I => \N__47295\
        );

    \I__9107\ : Span4Mux_h
    port map (
            O => \N__47302\,
            I => \N__47290\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__47299\,
            I => \N__47287\
        );

    \I__9105\ : InMux
    port map (
            O => \N__47298\,
            I => \N__47278\
        );

    \I__9104\ : InMux
    port map (
            O => \N__47295\,
            I => \N__47278\
        );

    \I__9103\ : InMux
    port map (
            O => \N__47294\,
            I => \N__47278\
        );

    \I__9102\ : InMux
    port map (
            O => \N__47293\,
            I => \N__47278\
        );

    \I__9101\ : Span4Mux_h
    port map (
            O => \N__47290\,
            I => \N__47271\
        );

    \I__9100\ : Span4Mux_v
    port map (
            O => \N__47287\,
            I => \N__47271\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__47278\,
            I => \N__47268\
        );

    \I__9098\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47265\
        );

    \I__9097\ : InMux
    port map (
            O => \N__47276\,
            I => \N__47262\
        );

    \I__9096\ : Span4Mux_v
    port map (
            O => \N__47271\,
            I => \N__47259\
        );

    \I__9095\ : Span12Mux_s11_v
    port map (
            O => \N__47268\,
            I => \N__47256\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__47265\,
            I => control_mode_2
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__47262\,
            I => control_mode_2
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__47259\,
            I => control_mode_2
        );

    \I__9091\ : Odrv12
    port map (
            O => \N__47256\,
            I => control_mode_2
        );

    \I__9090\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47244\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__47244\,
            I => \c0.n24539\
        );

    \I__9088\ : InMux
    port map (
            O => \N__47241\,
            I => \N__47238\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__47238\,
            I => \c0.n24733\
        );

    \I__9086\ : InMux
    port map (
            O => \N__47235\,
            I => \N__47228\
        );

    \I__9085\ : InMux
    port map (
            O => \N__47234\,
            I => \N__47224\
        );

    \I__9084\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47221\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__47232\,
            I => \N__47218\
        );

    \I__9082\ : InMux
    port map (
            O => \N__47231\,
            I => \N__47215\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__47228\,
            I => \N__47212\
        );

    \I__9080\ : InMux
    port map (
            O => \N__47227\,
            I => \N__47209\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__47224\,
            I => \N__47206\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__47221\,
            I => \N__47203\
        );

    \I__9077\ : InMux
    port map (
            O => \N__47218\,
            I => \N__47200\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__47215\,
            I => \N__47197\
        );

    \I__9075\ : Span4Mux_v
    port map (
            O => \N__47212\,
            I => \N__47194\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__47209\,
            I => \N__47191\
        );

    \I__9073\ : Span4Mux_v
    port map (
            O => \N__47206\,
            I => \N__47188\
        );

    \I__9072\ : Span4Mux_v
    port map (
            O => \N__47203\,
            I => \N__47183\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__47200\,
            I => \N__47183\
        );

    \I__9070\ : Span4Mux_v
    port map (
            O => \N__47197\,
            I => \N__47180\
        );

    \I__9069\ : Span4Mux_v
    port map (
            O => \N__47194\,
            I => \N__47174\
        );

    \I__9068\ : Span4Mux_v
    port map (
            O => \N__47191\,
            I => \N__47174\
        );

    \I__9067\ : Span4Mux_h
    port map (
            O => \N__47188\,
            I => \N__47167\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__47183\,
            I => \N__47167\
        );

    \I__9065\ : Span4Mux_h
    port map (
            O => \N__47180\,
            I => \N__47167\
        );

    \I__9064\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47164\
        );

    \I__9063\ : Sp12to4
    port map (
            O => \N__47174\,
            I => \N__47159\
        );

    \I__9062\ : Sp12to4
    port map (
            O => \N__47167\,
            I => \N__47159\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__47164\,
            I => \r_Bit_Index_0\
        );

    \I__9060\ : Odrv12
    port map (
            O => \N__47159\,
            I => \r_Bit_Index_0\
        );

    \I__9059\ : CascadeMux
    port map (
            O => \N__47154\,
            I => \c0.rx.n17834_cascade_\
        );

    \I__9058\ : InMux
    port map (
            O => \N__47151\,
            I => \N__47146\
        );

    \I__9057\ : InMux
    port map (
            O => \N__47150\,
            I => \N__47143\
        );

    \I__9056\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47139\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__47146\,
            I => \N__47136\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__47143\,
            I => \N__47133\
        );

    \I__9053\ : InMux
    port map (
            O => \N__47142\,
            I => \N__47130\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__47139\,
            I => \N__47127\
        );

    \I__9051\ : Span4Mux_h
    port map (
            O => \N__47136\,
            I => \N__47124\
        );

    \I__9050\ : Span4Mux_h
    port map (
            O => \N__47133\,
            I => \N__47121\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__47130\,
            I => \N__47118\
        );

    \I__9048\ : Span4Mux_v
    port map (
            O => \N__47127\,
            I => \N__47115\
        );

    \I__9047\ : Span4Mux_h
    port map (
            O => \N__47124\,
            I => \N__47112\
        );

    \I__9046\ : Odrv4
    port map (
            O => \N__47121\,
            I => n14484
        );

    \I__9045\ : Odrv4
    port map (
            O => \N__47118\,
            I => n14484
        );

    \I__9044\ : Odrv4
    port map (
            O => \N__47115\,
            I => n14484
        );

    \I__9043\ : Odrv4
    port map (
            O => \N__47112\,
            I => n14484
        );

    \I__9042\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47099\
        );

    \I__9041\ : InMux
    port map (
            O => \N__47102\,
            I => \N__47095\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__47092\
        );

    \I__9039\ : InMux
    port map (
            O => \N__47098\,
            I => \N__47089\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__47095\,
            I => \N__47086\
        );

    \I__9037\ : Span4Mux_v
    port map (
            O => \N__47092\,
            I => \N__47083\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__47089\,
            I => \N__47080\
        );

    \I__9035\ : Span4Mux_h
    port map (
            O => \N__47086\,
            I => \N__47077\
        );

    \I__9034\ : Span4Mux_h
    port map (
            O => \N__47083\,
            I => \N__47072\
        );

    \I__9033\ : Span4Mux_v
    port map (
            O => \N__47080\,
            I => \N__47072\
        );

    \I__9032\ : Span4Mux_v
    port map (
            O => \N__47077\,
            I => \N__47067\
        );

    \I__9031\ : Span4Mux_h
    port map (
            O => \N__47072\,
            I => \N__47067\
        );

    \I__9030\ : Odrv4
    port map (
            O => \N__47067\,
            I => n14988
        );

    \I__9029\ : InMux
    port map (
            O => \N__47064\,
            I => \N__47061\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__47061\,
            I => \N__47058\
        );

    \I__9027\ : Span4Mux_h
    port map (
            O => \N__47058\,
            I => \N__47054\
        );

    \I__9026\ : InMux
    port map (
            O => \N__47057\,
            I => \N__47048\
        );

    \I__9025\ : Span4Mux_h
    port map (
            O => \N__47054\,
            I => \N__47045\
        );

    \I__9024\ : InMux
    port map (
            O => \N__47053\,
            I => \N__47040\
        );

    \I__9023\ : InMux
    port map (
            O => \N__47052\,
            I => \N__47040\
        );

    \I__9022\ : InMux
    port map (
            O => \N__47051\,
            I => \N__47037\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__47048\,
            I => control_mode_5
        );

    \I__9020\ : Odrv4
    port map (
            O => \N__47045\,
            I => control_mode_5
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__47040\,
            I => control_mode_5
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__47037\,
            I => control_mode_5
        );

    \I__9017\ : InMux
    port map (
            O => \N__47028\,
            I => \N__47024\
        );

    \I__9016\ : CascadeMux
    port map (
            O => \N__47027\,
            I => \N__47021\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__47024\,
            I => \N__47018\
        );

    \I__9014\ : InMux
    port map (
            O => \N__47021\,
            I => \N__47015\
        );

    \I__9013\ : Span4Mux_h
    port map (
            O => \N__47018\,
            I => \N__47008\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__47015\,
            I => \N__47004\
        );

    \I__9011\ : InMux
    port map (
            O => \N__47014\,
            I => \N__47001\
        );

    \I__9010\ : InMux
    port map (
            O => \N__47013\,
            I => \N__46994\
        );

    \I__9009\ : InMux
    port map (
            O => \N__47012\,
            I => \N__46994\
        );

    \I__9008\ : InMux
    port map (
            O => \N__47011\,
            I => \N__46994\
        );

    \I__9007\ : Span4Mux_v
    port map (
            O => \N__47008\,
            I => \N__46991\
        );

    \I__9006\ : InMux
    port map (
            O => \N__47007\,
            I => \N__46988\
        );

    \I__9005\ : Span4Mux_h
    port map (
            O => \N__47004\,
            I => \N__46985\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__47001\,
            I => \N__46982\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__46994\,
            I => \N__46979\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__46991\,
            I => \N__46976\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__46988\,
            I => \N__46969\
        );

    \I__9000\ : Span4Mux_h
    port map (
            O => \N__46985\,
            I => \N__46969\
        );

    \I__8999\ : Span4Mux_v
    port map (
            O => \N__46982\,
            I => \N__46969\
        );

    \I__8998\ : Odrv12
    port map (
            O => \N__46979\,
            I => control_mode_1
        );

    \I__8997\ : Odrv4
    port map (
            O => \N__46976\,
            I => control_mode_1
        );

    \I__8996\ : Odrv4
    port map (
            O => \N__46969\,
            I => control_mode_1
        );

    \I__8995\ : CascadeMux
    port map (
            O => \N__46962\,
            I => \N__46959\
        );

    \I__8994\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46956\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__46956\,
            I => \N__46950\
        );

    \I__8992\ : InMux
    port map (
            O => \N__46955\,
            I => \N__46946\
        );

    \I__8991\ : InMux
    port map (
            O => \N__46954\,
            I => \N__46943\
        );

    \I__8990\ : InMux
    port map (
            O => \N__46953\,
            I => \N__46940\
        );

    \I__8989\ : Span12Mux_h
    port map (
            O => \N__46950\,
            I => \N__46937\
        );

    \I__8988\ : InMux
    port map (
            O => \N__46949\,
            I => \N__46934\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__46946\,
            I => \N__46929\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__46943\,
            I => \N__46929\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__46940\,
            I => control_mode_3
        );

    \I__8984\ : Odrv12
    port map (
            O => \N__46937\,
            I => control_mode_3
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__46934\,
            I => control_mode_3
        );

    \I__8982\ : Odrv12
    port map (
            O => \N__46929\,
            I => control_mode_3
        );

    \I__8981\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46915\
        );

    \I__8980\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46910\
        );

    \I__8979\ : InMux
    port map (
            O => \N__46918\,
            I => \N__46910\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__46915\,
            I => \N__46907\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__46910\,
            I => \N__46903\
        );

    \I__8976\ : Span4Mux_h
    port map (
            O => \N__46907\,
            I => \N__46900\
        );

    \I__8975\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46897\
        );

    \I__8974\ : Span4Mux_h
    port map (
            O => \N__46903\,
            I => \N__46894\
        );

    \I__8973\ : Odrv4
    port map (
            O => \N__46900\,
            I => data_in_2_3
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__46897\,
            I => data_in_2_3
        );

    \I__8971\ : Odrv4
    port map (
            O => \N__46894\,
            I => data_in_2_3
        );

    \I__8970\ : CascadeMux
    port map (
            O => \N__46887\,
            I => \c0.n82_cascade_\
        );

    \I__8969\ : InMux
    port map (
            O => \N__46884\,
            I => \N__46880\
        );

    \I__8968\ : InMux
    port map (
            O => \N__46883\,
            I => \N__46874\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__46880\,
            I => \N__46870\
        );

    \I__8966\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46867\
        );

    \I__8965\ : InMux
    port map (
            O => \N__46878\,
            I => \N__46864\
        );

    \I__8964\ : InMux
    port map (
            O => \N__46877\,
            I => \N__46861\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__46874\,
            I => \N__46858\
        );

    \I__8962\ : CascadeMux
    port map (
            O => \N__46873\,
            I => \N__46855\
        );

    \I__8961\ : Span4Mux_v
    port map (
            O => \N__46870\,
            I => \N__46851\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__46867\,
            I => \N__46846\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__46864\,
            I => \N__46846\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__46861\,
            I => \N__46841\
        );

    \I__8957\ : Span4Mux_v
    port map (
            O => \N__46858\,
            I => \N__46841\
        );

    \I__8956\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46836\
        );

    \I__8955\ : InMux
    port map (
            O => \N__46854\,
            I => \N__46836\
        );

    \I__8954\ : Odrv4
    port map (
            O => \N__46851\,
            I => \c0.n10467\
        );

    \I__8953\ : Odrv4
    port map (
            O => \N__46846\,
            I => \c0.n10467\
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__46841\,
            I => \c0.n10467\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__46836\,
            I => \c0.n10467\
        );

    \I__8950\ : CascadeMux
    port map (
            O => \N__46827\,
            I => \N__46819\
        );

    \I__8949\ : CascadeMux
    port map (
            O => \N__46826\,
            I => \N__46816\
        );

    \I__8948\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46808\
        );

    \I__8947\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46808\
        );

    \I__8946\ : InMux
    port map (
            O => \N__46823\,
            I => \N__46808\
        );

    \I__8945\ : InMux
    port map (
            O => \N__46822\,
            I => \N__46801\
        );

    \I__8944\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46801\
        );

    \I__8943\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46801\
        );

    \I__8942\ : InMux
    port map (
            O => \N__46815\,
            I => \N__46797\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__46808\,
            I => \N__46792\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__46801\,
            I => \N__46792\
        );

    \I__8939\ : InMux
    port map (
            O => \N__46800\,
            I => \N__46786\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__46797\,
            I => \N__46783\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__46792\,
            I => \N__46780\
        );

    \I__8936\ : InMux
    port map (
            O => \N__46791\,
            I => \N__46773\
        );

    \I__8935\ : InMux
    port map (
            O => \N__46790\,
            I => \N__46773\
        );

    \I__8934\ : InMux
    port map (
            O => \N__46789\,
            I => \N__46773\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__46786\,
            I => \N__46770\
        );

    \I__8932\ : Span4Mux_h
    port map (
            O => \N__46783\,
            I => \N__46767\
        );

    \I__8931\ : Span4Mux_h
    port map (
            O => \N__46780\,
            I => \N__46762\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46762\
        );

    \I__8929\ : Span4Mux_v
    port map (
            O => \N__46770\,
            I => \N__46759\
        );

    \I__8928\ : Odrv4
    port map (
            O => \N__46767\,
            I => \c0.n10500\
        );

    \I__8927\ : Odrv4
    port map (
            O => \N__46762\,
            I => \c0.n10500\
        );

    \I__8926\ : Odrv4
    port map (
            O => \N__46759\,
            I => \c0.n10500\
        );

    \I__8925\ : InMux
    port map (
            O => \N__46752\,
            I => \N__46749\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__46749\,
            I => \N__46746\
        );

    \I__8923\ : Span4Mux_h
    port map (
            O => \N__46746\,
            I => \N__46737\
        );

    \I__8922\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46732\
        );

    \I__8921\ : InMux
    port map (
            O => \N__46744\,
            I => \N__46732\
        );

    \I__8920\ : InMux
    port map (
            O => \N__46743\,
            I => \N__46723\
        );

    \I__8919\ : InMux
    port map (
            O => \N__46742\,
            I => \N__46723\
        );

    \I__8918\ : InMux
    port map (
            O => \N__46741\,
            I => \N__46723\
        );

    \I__8917\ : InMux
    port map (
            O => \N__46740\,
            I => \N__46723\
        );

    \I__8916\ : Odrv4
    port map (
            O => \N__46737\,
            I => \c0.n21349\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__46732\,
            I => \c0.n21349\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__46723\,
            I => \c0.n21349\
        );

    \I__8913\ : InMux
    port map (
            O => \N__46716\,
            I => \N__46713\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__46713\,
            I => \c0.n4_adj_4271\
        );

    \I__8911\ : InMux
    port map (
            O => \N__46710\,
            I => \N__46707\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__46707\,
            I => \c0.data_out_frame_29__6__N_1538\
        );

    \I__8909\ : InMux
    port map (
            O => \N__46704\,
            I => \N__46700\
        );

    \I__8908\ : InMux
    port map (
            O => \N__46703\,
            I => \N__46697\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__46700\,
            I => \N__46691\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__46697\,
            I => \N__46691\
        );

    \I__8905\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46688\
        );

    \I__8904\ : Span4Mux_v
    port map (
            O => \N__46691\,
            I => \N__46683\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__46688\,
            I => \N__46683\
        );

    \I__8902\ : Odrv4
    port map (
            O => \N__46683\,
            I => \c0.n21327\
        );

    \I__8901\ : CascadeMux
    port map (
            O => \N__46680\,
            I => \c0.n4_adj_4271_cascade_\
        );

    \I__8900\ : InMux
    port map (
            O => \N__46677\,
            I => \N__46674\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__46674\,
            I => \c0.data_out_frame_29__3__N_1730\
        );

    \I__8898\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46667\
        );

    \I__8897\ : InMux
    port map (
            O => \N__46670\,
            I => \N__46664\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__46667\,
            I => \N__46661\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__46664\,
            I => \data_out_frame_29__3__N_1661\
        );

    \I__8894\ : Odrv4
    port map (
            O => \N__46661\,
            I => \data_out_frame_29__3__N_1661\
        );

    \I__8893\ : InMux
    port map (
            O => \N__46656\,
            I => \N__46653\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__46653\,
            I => \N__46649\
        );

    \I__8891\ : InMux
    port map (
            O => \N__46652\,
            I => \N__46646\
        );

    \I__8890\ : Span4Mux_v
    port map (
            O => \N__46649\,
            I => \N__46643\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__46646\,
            I => \N__46640\
        );

    \I__8888\ : Odrv4
    port map (
            O => \N__46643\,
            I => \c0.rx.n12909\
        );

    \I__8887\ : Odrv4
    port map (
            O => \N__46640\,
            I => \c0.rx.n12909\
        );

    \I__8886\ : CascadeMux
    port map (
            O => \N__46635\,
            I => \c0.n22112_cascade_\
        );

    \I__8885\ : InMux
    port map (
            O => \N__46632\,
            I => \N__46628\
        );

    \I__8884\ : InMux
    port map (
            O => \N__46631\,
            I => \N__46625\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__46628\,
            I => \N__46620\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__46625\,
            I => \N__46620\
        );

    \I__8881\ : Span4Mux_v
    port map (
            O => \N__46620\,
            I => \N__46617\
        );

    \I__8880\ : Odrv4
    port map (
            O => \N__46617\,
            I => \c0.n21355\
        );

    \I__8879\ : InMux
    port map (
            O => \N__46614\,
            I => \N__46611\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__46611\,
            I => \N__46603\
        );

    \I__8877\ : InMux
    port map (
            O => \N__46610\,
            I => \N__46600\
        );

    \I__8876\ : InMux
    port map (
            O => \N__46609\,
            I => \N__46594\
        );

    \I__8875\ : InMux
    port map (
            O => \N__46608\,
            I => \N__46594\
        );

    \I__8874\ : InMux
    port map (
            O => \N__46607\,
            I => \N__46591\
        );

    \I__8873\ : InMux
    port map (
            O => \N__46606\,
            I => \N__46587\
        );

    \I__8872\ : Sp12to4
    port map (
            O => \N__46603\,
            I => \N__46582\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__46600\,
            I => \N__46582\
        );

    \I__8870\ : InMux
    port map (
            O => \N__46599\,
            I => \N__46579\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__46594\,
            I => \N__46576\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__46591\,
            I => \N__46573\
        );

    \I__8867\ : InMux
    port map (
            O => \N__46590\,
            I => \N__46570\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__46587\,
            I => \c0.n12604\
        );

    \I__8865\ : Odrv12
    port map (
            O => \N__46582\,
            I => \c0.n12604\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__46579\,
            I => \c0.n12604\
        );

    \I__8863\ : Odrv4
    port map (
            O => \N__46576\,
            I => \c0.n12604\
        );

    \I__8862\ : Odrv4
    port map (
            O => \N__46573\,
            I => \c0.n12604\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__46570\,
            I => \c0.n12604\
        );

    \I__8860\ : InMux
    port map (
            O => \N__46557\,
            I => \N__46554\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__46554\,
            I => \N__46550\
        );

    \I__8858\ : InMux
    port map (
            O => \N__46553\,
            I => \N__46547\
        );

    \I__8857\ : Odrv12
    port map (
            O => \N__46550\,
            I => \c0.n20786\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__46547\,
            I => \c0.n20786\
        );

    \I__8855\ : CascadeMux
    port map (
            O => \N__46542\,
            I => \c0.n20786_cascade_\
        );

    \I__8854\ : InMux
    port map (
            O => \N__46539\,
            I => \N__46536\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__46536\,
            I => \c0.n9_adj_4494\
        );

    \I__8852\ : InMux
    port map (
            O => \N__46533\,
            I => \N__46529\
        );

    \I__8851\ : InMux
    port map (
            O => \N__46532\,
            I => \N__46526\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__46529\,
            I => \N__46523\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__46526\,
            I => \N__46519\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__46523\,
            I => \N__46516\
        );

    \I__8847\ : InMux
    port map (
            O => \N__46522\,
            I => \N__46513\
        );

    \I__8846\ : Span4Mux_h
    port map (
            O => \N__46519\,
            I => \N__46510\
        );

    \I__8845\ : Span4Mux_h
    port map (
            O => \N__46516\,
            I => \N__46505\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__46513\,
            I => \N__46505\
        );

    \I__8843\ : Odrv4
    port map (
            O => \N__46510\,
            I => \c0.n10497\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__46505\,
            I => \c0.n10497\
        );

    \I__8841\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46493\
        );

    \I__8840\ : InMux
    port map (
            O => \N__46499\,
            I => \N__46493\
        );

    \I__8839\ : InMux
    port map (
            O => \N__46498\,
            I => \N__46490\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__46493\,
            I => \c0.n21433\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__46490\,
            I => \c0.n21433\
        );

    \I__8836\ : CascadeMux
    port map (
            O => \N__46485\,
            I => \N__46479\
        );

    \I__8835\ : InMux
    port map (
            O => \N__46484\,
            I => \N__46475\
        );

    \I__8834\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46466\
        );

    \I__8833\ : InMux
    port map (
            O => \N__46482\,
            I => \N__46466\
        );

    \I__8832\ : InMux
    port map (
            O => \N__46479\,
            I => \N__46466\
        );

    \I__8831\ : InMux
    port map (
            O => \N__46478\,
            I => \N__46466\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__46475\,
            I => \c0.n21311\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__46466\,
            I => \c0.n21311\
        );

    \I__8828\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46457\
        );

    \I__8827\ : InMux
    port map (
            O => \N__46460\,
            I => \N__46454\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__46457\,
            I => \c0.n12590\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__46454\,
            I => \c0.n12590\
        );

    \I__8824\ : InMux
    port map (
            O => \N__46449\,
            I => \N__46445\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__46448\,
            I => \N__46441\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__46445\,
            I => \N__46437\
        );

    \I__8821\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46434\
        );

    \I__8820\ : InMux
    port map (
            O => \N__46441\,
            I => \N__46431\
        );

    \I__8819\ : InMux
    port map (
            O => \N__46440\,
            I => \N__46428\
        );

    \I__8818\ : Span4Mux_h
    port map (
            O => \N__46437\,
            I => \N__46425\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__46434\,
            I => \N__46422\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__46431\,
            I => \N__46417\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__46428\,
            I => \N__46417\
        );

    \I__8814\ : Span4Mux_h
    port map (
            O => \N__46425\,
            I => \N__46414\
        );

    \I__8813\ : Span4Mux_v
    port map (
            O => \N__46422\,
            I => \N__46411\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__46417\,
            I => \N__46408\
        );

    \I__8811\ : Span4Mux_v
    port map (
            O => \N__46414\,
            I => \N__46405\
        );

    \I__8810\ : Span4Mux_h
    port map (
            O => \N__46411\,
            I => \N__46402\
        );

    \I__8809\ : Odrv4
    port map (
            O => \N__46408\,
            I => \c0.n21399\
        );

    \I__8808\ : Odrv4
    port map (
            O => \N__46405\,
            I => \c0.n21399\
        );

    \I__8807\ : Odrv4
    port map (
            O => \N__46402\,
            I => \c0.n21399\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__46395\,
            I => \N__46392\
        );

    \I__8805\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46388\
        );

    \I__8804\ : InMux
    port map (
            O => \N__46391\,
            I => \N__46385\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__46388\,
            I => \N__46382\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__46385\,
            I => \N__46379\
        );

    \I__8801\ : Span4Mux_v
    port map (
            O => \N__46382\,
            I => \N__46373\
        );

    \I__8800\ : Span4Mux_v
    port map (
            O => \N__46379\,
            I => \N__46373\
        );

    \I__8799\ : InMux
    port map (
            O => \N__46378\,
            I => \N__46370\
        );

    \I__8798\ : Span4Mux_h
    port map (
            O => \N__46373\,
            I => \N__46365\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__46370\,
            I => \N__46365\
        );

    \I__8796\ : Odrv4
    port map (
            O => \N__46365\,
            I => \c0.n22553\
        );

    \I__8795\ : CascadeMux
    port map (
            O => \N__46362\,
            I => \N__46358\
        );

    \I__8794\ : CascadeMux
    port map (
            O => \N__46361\,
            I => \N__46353\
        );

    \I__8793\ : InMux
    port map (
            O => \N__46358\,
            I => \N__46350\
        );

    \I__8792\ : InMux
    port map (
            O => \N__46357\,
            I => \N__46345\
        );

    \I__8791\ : InMux
    port map (
            O => \N__46356\,
            I => \N__46342\
        );

    \I__8790\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46339\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__46350\,
            I => \N__46336\
        );

    \I__8788\ : InMux
    port map (
            O => \N__46349\,
            I => \N__46333\
        );

    \I__8787\ : InMux
    port map (
            O => \N__46348\,
            I => \N__46330\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__46345\,
            I => \N__46326\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__46342\,
            I => \N__46323\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__46339\,
            I => \N__46320\
        );

    \I__8783\ : Span4Mux_v
    port map (
            O => \N__46336\,
            I => \N__46315\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__46333\,
            I => \N__46315\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__46330\,
            I => \N__46311\
        );

    \I__8780\ : InMux
    port map (
            O => \N__46329\,
            I => \N__46308\
        );

    \I__8779\ : Span4Mux_v
    port map (
            O => \N__46326\,
            I => \N__46305\
        );

    \I__8778\ : Span4Mux_h
    port map (
            O => \N__46323\,
            I => \N__46302\
        );

    \I__8777\ : Span4Mux_v
    port map (
            O => \N__46320\,
            I => \N__46297\
        );

    \I__8776\ : Span4Mux_h
    port map (
            O => \N__46315\,
            I => \N__46297\
        );

    \I__8775\ : InMux
    port map (
            O => \N__46314\,
            I => \N__46294\
        );

    \I__8774\ : Span4Mux_v
    port map (
            O => \N__46311\,
            I => \N__46289\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__46308\,
            I => \N__46289\
        );

    \I__8772\ : Span4Mux_v
    port map (
            O => \N__46305\,
            I => \N__46286\
        );

    \I__8771\ : Span4Mux_v
    port map (
            O => \N__46302\,
            I => \N__46281\
        );

    \I__8770\ : Span4Mux_h
    port map (
            O => \N__46297\,
            I => \N__46281\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__46294\,
            I => encoder1_position_2
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__46289\,
            I => encoder1_position_2
        );

    \I__8767\ : Odrv4
    port map (
            O => \N__46286\,
            I => encoder1_position_2
        );

    \I__8766\ : Odrv4
    port map (
            O => \N__46281\,
            I => encoder1_position_2
        );

    \I__8765\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46265\
        );

    \I__8764\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46265\
        );

    \I__8763\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46261\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__46265\,
            I => \N__46258\
        );

    \I__8761\ : CascadeMux
    port map (
            O => \N__46264\,
            I => \N__46255\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__46261\,
            I => \N__46251\
        );

    \I__8759\ : Span4Mux_h
    port map (
            O => \N__46258\,
            I => \N__46248\
        );

    \I__8758\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46244\
        );

    \I__8757\ : InMux
    port map (
            O => \N__46254\,
            I => \N__46241\
        );

    \I__8756\ : Span4Mux_h
    port map (
            O => \N__46251\,
            I => \N__46236\
        );

    \I__8755\ : Span4Mux_h
    port map (
            O => \N__46248\,
            I => \N__46236\
        );

    \I__8754\ : InMux
    port map (
            O => \N__46247\,
            I => \N__46233\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__46244\,
            I => \N__46228\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__46241\,
            I => \N__46228\
        );

    \I__8751\ : Odrv4
    port map (
            O => \N__46236\,
            I => \c0.n21416\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__46233\,
            I => \c0.n21416\
        );

    \I__8749\ : Odrv4
    port map (
            O => \N__46228\,
            I => \c0.n21416\
        );

    \I__8748\ : InMux
    port map (
            O => \N__46221\,
            I => \N__46217\
        );

    \I__8747\ : InMux
    port map (
            O => \N__46220\,
            I => \N__46214\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__46217\,
            I => \N__46210\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__46214\,
            I => \N__46207\
        );

    \I__8744\ : InMux
    port map (
            O => \N__46213\,
            I => \N__46204\
        );

    \I__8743\ : Span4Mux_h
    port map (
            O => \N__46210\,
            I => \N__46199\
        );

    \I__8742\ : Span4Mux_v
    port map (
            O => \N__46207\,
            I => \N__46199\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__46204\,
            I => \N__46196\
        );

    \I__8740\ : Sp12to4
    port map (
            O => \N__46199\,
            I => \N__46191\
        );

    \I__8739\ : Span12Mux_s11_h
    port map (
            O => \N__46196\,
            I => \N__46191\
        );

    \I__8738\ : Odrv12
    port map (
            O => \N__46191\,
            I => \c0.n10531\
        );

    \I__8737\ : InMux
    port map (
            O => \N__46188\,
            I => \N__46185\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__46185\,
            I => \N__46180\
        );

    \I__8735\ : InMux
    port map (
            O => \N__46184\,
            I => \N__46174\
        );

    \I__8734\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46174\
        );

    \I__8733\ : Span4Mux_h
    port map (
            O => \N__46180\,
            I => \N__46171\
        );

    \I__8732\ : InMux
    port map (
            O => \N__46179\,
            I => \N__46168\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__46174\,
            I => \N__46165\
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__46171\,
            I => \c0.n20511\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__46168\,
            I => \c0.n20511\
        );

    \I__8728\ : Odrv12
    port map (
            O => \N__46165\,
            I => \c0.n20511\
        );

    \I__8727\ : CascadeMux
    port map (
            O => \N__46158\,
            I => \c0.n10531_cascade_\
        );

    \I__8726\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46152\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__46152\,
            I => \N__46148\
        );

    \I__8724\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46145\
        );

    \I__8723\ : Odrv4
    port map (
            O => \N__46148\,
            I => \c0.n21451\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__46145\,
            I => \c0.n21451\
        );

    \I__8721\ : CascadeMux
    port map (
            O => \N__46140\,
            I => \N__46136\
        );

    \I__8720\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46129\
        );

    \I__8719\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46122\
        );

    \I__8718\ : InMux
    port map (
            O => \N__46135\,
            I => \N__46122\
        );

    \I__8717\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46122\
        );

    \I__8716\ : InMux
    port map (
            O => \N__46133\,
            I => \N__46119\
        );

    \I__8715\ : InMux
    port map (
            O => \N__46132\,
            I => \N__46116\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__46129\,
            I => \N__46113\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__46122\,
            I => \N__46106\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__46119\,
            I => \N__46106\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__46116\,
            I => \N__46106\
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__46113\,
            I => \c0.n21437\
        );

    \I__8709\ : Odrv12
    port map (
            O => \N__46106\,
            I => \c0.n21437\
        );

    \I__8708\ : CascadeMux
    port map (
            O => \N__46101\,
            I => \c0.n21451_cascade_\
        );

    \I__8707\ : InMux
    port map (
            O => \N__46098\,
            I => \N__46080\
        );

    \I__8706\ : InMux
    port map (
            O => \N__46097\,
            I => \N__46071\
        );

    \I__8705\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46071\
        );

    \I__8704\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46071\
        );

    \I__8703\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46064\
        );

    \I__8702\ : InMux
    port map (
            O => \N__46093\,
            I => \N__46064\
        );

    \I__8701\ : InMux
    port map (
            O => \N__46092\,
            I => \N__46064\
        );

    \I__8700\ : InMux
    port map (
            O => \N__46091\,
            I => \N__46052\
        );

    \I__8699\ : InMux
    port map (
            O => \N__46090\,
            I => \N__46044\
        );

    \I__8698\ : InMux
    port map (
            O => \N__46089\,
            I => \N__46041\
        );

    \I__8697\ : InMux
    port map (
            O => \N__46088\,
            I => \N__46032\
        );

    \I__8696\ : InMux
    port map (
            O => \N__46087\,
            I => \N__46032\
        );

    \I__8695\ : InMux
    port map (
            O => \N__46086\,
            I => \N__46032\
        );

    \I__8694\ : InMux
    port map (
            O => \N__46085\,
            I => \N__46032\
        );

    \I__8693\ : InMux
    port map (
            O => \N__46084\,
            I => \N__46027\
        );

    \I__8692\ : InMux
    port map (
            O => \N__46083\,
            I => \N__46015\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__46080\,
            I => \N__46012\
        );

    \I__8690\ : InMux
    port map (
            O => \N__46079\,
            I => \N__46005\
        );

    \I__8689\ : InMux
    port map (
            O => \N__46078\,
            I => \N__46005\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__46071\,
            I => \N__46002\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__46064\,
            I => \N__45999\
        );

    \I__8686\ : InMux
    port map (
            O => \N__46063\,
            I => \N__45972\
        );

    \I__8685\ : InMux
    port map (
            O => \N__46062\,
            I => \N__45972\
        );

    \I__8684\ : InMux
    port map (
            O => \N__46061\,
            I => \N__45972\
        );

    \I__8683\ : InMux
    port map (
            O => \N__46060\,
            I => \N__45972\
        );

    \I__8682\ : InMux
    port map (
            O => \N__46059\,
            I => \N__45972\
        );

    \I__8681\ : InMux
    port map (
            O => \N__46058\,
            I => \N__45963\
        );

    \I__8680\ : InMux
    port map (
            O => \N__46057\,
            I => \N__45963\
        );

    \I__8679\ : InMux
    port map (
            O => \N__46056\,
            I => \N__45963\
        );

    \I__8678\ : InMux
    port map (
            O => \N__46055\,
            I => \N__45963\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__46052\,
            I => \N__45960\
        );

    \I__8676\ : InMux
    port map (
            O => \N__46051\,
            I => \N__45949\
        );

    \I__8675\ : InMux
    port map (
            O => \N__46050\,
            I => \N__45949\
        );

    \I__8674\ : InMux
    port map (
            O => \N__46049\,
            I => \N__45949\
        );

    \I__8673\ : InMux
    port map (
            O => \N__46048\,
            I => \N__45949\
        );

    \I__8672\ : InMux
    port map (
            O => \N__46047\,
            I => \N__45949\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__46044\,
            I => \N__45946\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__46041\,
            I => \N__45940\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__46032\,
            I => \N__45940\
        );

    \I__8668\ : InMux
    port map (
            O => \N__46031\,
            I => \N__45937\
        );

    \I__8667\ : InMux
    port map (
            O => \N__46030\,
            I => \N__45933\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__46027\,
            I => \N__45930\
        );

    \I__8665\ : InMux
    port map (
            O => \N__46026\,
            I => \N__45927\
        );

    \I__8664\ : InMux
    port map (
            O => \N__46025\,
            I => \N__45922\
        );

    \I__8663\ : InMux
    port map (
            O => \N__46024\,
            I => \N__45922\
        );

    \I__8662\ : InMux
    port map (
            O => \N__46023\,
            I => \N__45919\
        );

    \I__8661\ : InMux
    port map (
            O => \N__46022\,
            I => \N__45914\
        );

    \I__8660\ : InMux
    port map (
            O => \N__46021\,
            I => \N__45914\
        );

    \I__8659\ : InMux
    port map (
            O => \N__46020\,
            I => \N__45907\
        );

    \I__8658\ : InMux
    port map (
            O => \N__46019\,
            I => \N__45907\
        );

    \I__8657\ : InMux
    port map (
            O => \N__46018\,
            I => \N__45907\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__46015\,
            I => \N__45902\
        );

    \I__8655\ : Span4Mux_h
    port map (
            O => \N__46012\,
            I => \N__45902\
        );

    \I__8654\ : InMux
    port map (
            O => \N__46011\,
            I => \N__45897\
        );

    \I__8653\ : InMux
    port map (
            O => \N__46010\,
            I => \N__45897\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__46005\,
            I => \N__45890\
        );

    \I__8651\ : Span4Mux_h
    port map (
            O => \N__46002\,
            I => \N__45890\
        );

    \I__8650\ : Span4Mux_h
    port map (
            O => \N__45999\,
            I => \N__45890\
        );

    \I__8649\ : CascadeMux
    port map (
            O => \N__45998\,
            I => \N__45886\
        );

    \I__8648\ : CascadeMux
    port map (
            O => \N__45997\,
            I => \N__45883\
        );

    \I__8647\ : InMux
    port map (
            O => \N__45996\,
            I => \N__45864\
        );

    \I__8646\ : InMux
    port map (
            O => \N__45995\,
            I => \N__45864\
        );

    \I__8645\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45864\
        );

    \I__8644\ : InMux
    port map (
            O => \N__45993\,
            I => \N__45859\
        );

    \I__8643\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45859\
        );

    \I__8642\ : InMux
    port map (
            O => \N__45991\,
            I => \N__45852\
        );

    \I__8641\ : InMux
    port map (
            O => \N__45990\,
            I => \N__45852\
        );

    \I__8640\ : InMux
    port map (
            O => \N__45989\,
            I => \N__45852\
        );

    \I__8639\ : InMux
    port map (
            O => \N__45988\,
            I => \N__45839\
        );

    \I__8638\ : InMux
    port map (
            O => \N__45987\,
            I => \N__45839\
        );

    \I__8637\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45839\
        );

    \I__8636\ : InMux
    port map (
            O => \N__45985\,
            I => \N__45839\
        );

    \I__8635\ : InMux
    port map (
            O => \N__45984\,
            I => \N__45839\
        );

    \I__8634\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45839\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__45972\,
            I => \N__45832\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__45963\,
            I => \N__45832\
        );

    \I__8631\ : Span4Mux_v
    port map (
            O => \N__45960\,
            I => \N__45832\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__45949\,
            I => \N__45827\
        );

    \I__8629\ : Span4Mux_v
    port map (
            O => \N__45946\,
            I => \N__45827\
        );

    \I__8628\ : InMux
    port map (
            O => \N__45945\,
            I => \N__45824\
        );

    \I__8627\ : Span4Mux_v
    port map (
            O => \N__45940\,
            I => \N__45821\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__45937\,
            I => \N__45818\
        );

    \I__8625\ : InMux
    port map (
            O => \N__45936\,
            I => \N__45815\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__45933\,
            I => \N__45812\
        );

    \I__8623\ : Span4Mux_v
    port map (
            O => \N__45930\,
            I => \N__45809\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__45927\,
            I => \N__45796\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__45922\,
            I => \N__45796\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__45919\,
            I => \N__45796\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__45914\,
            I => \N__45796\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__45907\,
            I => \N__45796\
        );

    \I__8617\ : Span4Mux_v
    port map (
            O => \N__45902\,
            I => \N__45796\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__45897\,
            I => \N__45791\
        );

    \I__8615\ : Span4Mux_v
    port map (
            O => \N__45890\,
            I => \N__45791\
        );

    \I__8614\ : InMux
    port map (
            O => \N__45889\,
            I => \N__45788\
        );

    \I__8613\ : InMux
    port map (
            O => \N__45886\,
            I => \N__45785\
        );

    \I__8612\ : InMux
    port map (
            O => \N__45883\,
            I => \N__45782\
        );

    \I__8611\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45775\
        );

    \I__8610\ : InMux
    port map (
            O => \N__45881\,
            I => \N__45775\
        );

    \I__8609\ : InMux
    port map (
            O => \N__45880\,
            I => \N__45775\
        );

    \I__8608\ : InMux
    port map (
            O => \N__45879\,
            I => \N__45766\
        );

    \I__8607\ : InMux
    port map (
            O => \N__45878\,
            I => \N__45766\
        );

    \I__8606\ : InMux
    port map (
            O => \N__45877\,
            I => \N__45766\
        );

    \I__8605\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45766\
        );

    \I__8604\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45755\
        );

    \I__8603\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45755\
        );

    \I__8602\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45755\
        );

    \I__8601\ : InMux
    port map (
            O => \N__45872\,
            I => \N__45755\
        );

    \I__8600\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45755\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__45864\,
            I => \N__45752\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__45859\,
            I => \N__45741\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__45852\,
            I => \N__45741\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__45839\,
            I => \N__45741\
        );

    \I__8595\ : Span4Mux_h
    port map (
            O => \N__45832\,
            I => \N__45741\
        );

    \I__8594\ : Span4Mux_h
    port map (
            O => \N__45827\,
            I => \N__45741\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__45824\,
            I => \N__45734\
        );

    \I__8592\ : Sp12to4
    port map (
            O => \N__45821\,
            I => \N__45734\
        );

    \I__8591\ : Span12Mux_v
    port map (
            O => \N__45818\,
            I => \N__45734\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__45815\,
            I => \N__45723\
        );

    \I__8589\ : Span4Mux_v
    port map (
            O => \N__45812\,
            I => \N__45723\
        );

    \I__8588\ : Span4Mux_h
    port map (
            O => \N__45809\,
            I => \N__45723\
        );

    \I__8587\ : Span4Mux_v
    port map (
            O => \N__45796\,
            I => \N__45723\
        );

    \I__8586\ : Span4Mux_v
    port map (
            O => \N__45791\,
            I => \N__45723\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__45788\,
            I => \N__45718\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__45785\,
            I => \N__45718\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__45782\,
            I => n13058
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__45775\,
            I => n13058
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__45766\,
            I => n13058
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__45755\,
            I => n13058
        );

    \I__8579\ : Odrv12
    port map (
            O => \N__45752\,
            I => n13058
        );

    \I__8578\ : Odrv4
    port map (
            O => \N__45741\,
            I => n13058
        );

    \I__8577\ : Odrv12
    port map (
            O => \N__45734\,
            I => n13058
        );

    \I__8576\ : Odrv4
    port map (
            O => \N__45723\,
            I => n13058
        );

    \I__8575\ : Odrv4
    port map (
            O => \N__45718\,
            I => n13058
        );

    \I__8574\ : InMux
    port map (
            O => \N__45699\,
            I => \N__45696\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__45696\,
            I => \N__45693\
        );

    \I__8572\ : Span4Mux_v
    port map (
            O => \N__45693\,
            I => \N__45689\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__45692\,
            I => \N__45686\
        );

    \I__8570\ : Span4Mux_h
    port map (
            O => \N__45689\,
            I => \N__45683\
        );

    \I__8569\ : InMux
    port map (
            O => \N__45686\,
            I => \N__45680\
        );

    \I__8568\ : Span4Mux_v
    port map (
            O => \N__45683\,
            I => \N__45677\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__45680\,
            I => data_out_frame_8_6
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__45677\,
            I => data_out_frame_8_6
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__45672\,
            I => \N__45669\
        );

    \I__8564\ : InMux
    port map (
            O => \N__45669\,
            I => \N__45666\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__45666\,
            I => \N__45663\
        );

    \I__8562\ : Span4Mux_h
    port map (
            O => \N__45663\,
            I => \N__45660\
        );

    \I__8561\ : Span4Mux_v
    port map (
            O => \N__45660\,
            I => \N__45657\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__45657\,
            I => \N__45652\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__45656\,
            I => \N__45649\
        );

    \I__8558\ : InMux
    port map (
            O => \N__45655\,
            I => \N__45645\
        );

    \I__8557\ : Span4Mux_v
    port map (
            O => \N__45652\,
            I => \N__45642\
        );

    \I__8556\ : InMux
    port map (
            O => \N__45649\,
            I => \N__45639\
        );

    \I__8555\ : InMux
    port map (
            O => \N__45648\,
            I => \N__45636\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__45645\,
            I => encoder0_position_21
        );

    \I__8553\ : Odrv4
    port map (
            O => \N__45642\,
            I => encoder0_position_21
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__45639\,
            I => encoder0_position_21
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__45636\,
            I => encoder0_position_21
        );

    \I__8550\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45623\
        );

    \I__8549\ : InMux
    port map (
            O => \N__45626\,
            I => \N__45620\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__45623\,
            I => \c0.n22252\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__45620\,
            I => \c0.n22252\
        );

    \I__8546\ : CascadeMux
    port map (
            O => \N__45615\,
            I => \N__45609\
        );

    \I__8545\ : CascadeMux
    port map (
            O => \N__45614\,
            I => \N__45606\
        );

    \I__8544\ : CascadeMux
    port map (
            O => \N__45613\,
            I => \N__45603\
        );

    \I__8543\ : InMux
    port map (
            O => \N__45612\,
            I => \N__45599\
        );

    \I__8542\ : InMux
    port map (
            O => \N__45609\,
            I => \N__45595\
        );

    \I__8541\ : InMux
    port map (
            O => \N__45606\,
            I => \N__45592\
        );

    \I__8540\ : InMux
    port map (
            O => \N__45603\,
            I => \N__45588\
        );

    \I__8539\ : InMux
    port map (
            O => \N__45602\,
            I => \N__45584\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__45599\,
            I => \N__45581\
        );

    \I__8537\ : InMux
    port map (
            O => \N__45598\,
            I => \N__45578\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__45595\,
            I => \N__45573\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__45592\,
            I => \N__45573\
        );

    \I__8534\ : InMux
    port map (
            O => \N__45591\,
            I => \N__45570\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__45588\,
            I => \N__45567\
        );

    \I__8532\ : InMux
    port map (
            O => \N__45587\,
            I => \N__45564\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__45584\,
            I => \N__45561\
        );

    \I__8530\ : Span4Mux_v
    port map (
            O => \N__45581\,
            I => \N__45556\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__45578\,
            I => \N__45556\
        );

    \I__8528\ : Span4Mux_h
    port map (
            O => \N__45573\,
            I => \N__45549\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__45570\,
            I => \N__45549\
        );

    \I__8526\ : Span4Mux_h
    port map (
            O => \N__45567\,
            I => \N__45549\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__45564\,
            I => encoder0_position_27
        );

    \I__8524\ : Odrv12
    port map (
            O => \N__45561\,
            I => encoder0_position_27
        );

    \I__8523\ : Odrv4
    port map (
            O => \N__45556\,
            I => encoder0_position_27
        );

    \I__8522\ : Odrv4
    port map (
            O => \N__45549\,
            I => encoder0_position_27
        );

    \I__8521\ : InMux
    port map (
            O => \N__45540\,
            I => \N__45537\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__45537\,
            I => \N__45534\
        );

    \I__8519\ : Span4Mux_v
    port map (
            O => \N__45534\,
            I => \N__45530\
        );

    \I__8518\ : InMux
    port map (
            O => \N__45533\,
            I => \N__45527\
        );

    \I__8517\ : Span4Mux_h
    port map (
            O => \N__45530\,
            I => \N__45524\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__45527\,
            I => data_out_frame_6_3
        );

    \I__8515\ : Odrv4
    port map (
            O => \N__45524\,
            I => data_out_frame_6_3
        );

    \I__8514\ : InMux
    port map (
            O => \N__45519\,
            I => \N__45514\
        );

    \I__8513\ : InMux
    port map (
            O => \N__45518\,
            I => \N__45511\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__45517\,
            I => \N__45508\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__45514\,
            I => \N__45502\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__45511\,
            I => \N__45499\
        );

    \I__8509\ : InMux
    port map (
            O => \N__45508\,
            I => \N__45494\
        );

    \I__8508\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45494\
        );

    \I__8507\ : InMux
    port map (
            O => \N__45506\,
            I => \N__45490\
        );

    \I__8506\ : InMux
    port map (
            O => \N__45505\,
            I => \N__45487\
        );

    \I__8505\ : Span4Mux_v
    port map (
            O => \N__45502\,
            I => \N__45480\
        );

    \I__8504\ : Span4Mux_h
    port map (
            O => \N__45499\,
            I => \N__45480\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__45494\,
            I => \N__45480\
        );

    \I__8502\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45476\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__45490\,
            I => \N__45473\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__45487\,
            I => \N__45470\
        );

    \I__8499\ : Span4Mux_v
    port map (
            O => \N__45480\,
            I => \N__45467\
        );

    \I__8498\ : InMux
    port map (
            O => \N__45479\,
            I => \N__45464\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__45476\,
            I => \N__45461\
        );

    \I__8496\ : Span12Mux_s7_v
    port map (
            O => \N__45473\,
            I => \N__45458\
        );

    \I__8495\ : Span4Mux_v
    port map (
            O => \N__45470\,
            I => \N__45453\
        );

    \I__8494\ : Span4Mux_h
    port map (
            O => \N__45467\,
            I => \N__45453\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__45464\,
            I => encoder1_position_3
        );

    \I__8492\ : Odrv4
    port map (
            O => \N__45461\,
            I => encoder1_position_3
        );

    \I__8491\ : Odrv12
    port map (
            O => \N__45458\,
            I => encoder1_position_3
        );

    \I__8490\ : Odrv4
    port map (
            O => \N__45453\,
            I => encoder1_position_3
        );

    \I__8489\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45441\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__45441\,
            I => \N__45433\
        );

    \I__8487\ : InMux
    port map (
            O => \N__45440\,
            I => \N__45430\
        );

    \I__8486\ : InMux
    port map (
            O => \N__45439\,
            I => \N__45425\
        );

    \I__8485\ : InMux
    port map (
            O => \N__45438\,
            I => \N__45425\
        );

    \I__8484\ : InMux
    port map (
            O => \N__45437\,
            I => \N__45422\
        );

    \I__8483\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45419\
        );

    \I__8482\ : Span4Mux_v
    port map (
            O => \N__45433\,
            I => \N__45416\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__45430\,
            I => \N__45411\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__45425\,
            I => \N__45411\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__45422\,
            I => \N__45408\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__45419\,
            I => \c0.n20455\
        );

    \I__8477\ : Odrv4
    port map (
            O => \N__45416\,
            I => \c0.n20455\
        );

    \I__8476\ : Odrv12
    port map (
            O => \N__45411\,
            I => \c0.n20455\
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__45408\,
            I => \c0.n20455\
        );

    \I__8474\ : InMux
    port map (
            O => \N__45399\,
            I => \N__45396\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__45396\,
            I => \N__45393\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__45393\,
            I => \N__45389\
        );

    \I__8471\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45386\
        );

    \I__8470\ : Span4Mux_h
    port map (
            O => \N__45389\,
            I => \N__45383\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__45386\,
            I => \N__45377\
        );

    \I__8468\ : Span4Mux_v
    port map (
            O => \N__45383\,
            I => \N__45374\
        );

    \I__8467\ : InMux
    port map (
            O => \N__45382\,
            I => \N__45371\
        );

    \I__8466\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45368\
        );

    \I__8465\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45365\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__45377\,
            I => \N__45362\
        );

    \I__8463\ : Sp12to4
    port map (
            O => \N__45374\,
            I => \N__45357\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__45371\,
            I => \N__45357\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__45368\,
            I => encoder0_position_5
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__45365\,
            I => encoder0_position_5
        );

    \I__8459\ : Odrv4
    port map (
            O => \N__45362\,
            I => encoder0_position_5
        );

    \I__8458\ : Odrv12
    port map (
            O => \N__45357\,
            I => encoder0_position_5
        );

    \I__8457\ : InMux
    port map (
            O => \N__45348\,
            I => \N__45345\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__45345\,
            I => \N__45341\
        );

    \I__8455\ : CascadeMux
    port map (
            O => \N__45344\,
            I => \N__45337\
        );

    \I__8454\ : Span4Mux_h
    port map (
            O => \N__45341\,
            I => \N__45333\
        );

    \I__8453\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45330\
        );

    \I__8452\ : InMux
    port map (
            O => \N__45337\,
            I => \N__45327\
        );

    \I__8451\ : InMux
    port map (
            O => \N__45336\,
            I => \N__45324\
        );

    \I__8450\ : Span4Mux_v
    port map (
            O => \N__45333\,
            I => \N__45316\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__45330\,
            I => \N__45316\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__45327\,
            I => \N__45311\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__45324\,
            I => \N__45311\
        );

    \I__8446\ : CascadeMux
    port map (
            O => \N__45323\,
            I => \N__45308\
        );

    \I__8445\ : InMux
    port map (
            O => \N__45322\,
            I => \N__45305\
        );

    \I__8444\ : InMux
    port map (
            O => \N__45321\,
            I => \N__45302\
        );

    \I__8443\ : Span4Mux_v
    port map (
            O => \N__45316\,
            I => \N__45297\
        );

    \I__8442\ : Span4Mux_h
    port map (
            O => \N__45311\,
            I => \N__45297\
        );

    \I__8441\ : InMux
    port map (
            O => \N__45308\,
            I => \N__45294\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__45305\,
            I => encoder0_position_20
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__45302\,
            I => encoder0_position_20
        );

    \I__8438\ : Odrv4
    port map (
            O => \N__45297\,
            I => encoder0_position_20
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__45294\,
            I => encoder0_position_20
        );

    \I__8436\ : CascadeMux
    port map (
            O => \N__45285\,
            I => \N__45282\
        );

    \I__8435\ : InMux
    port map (
            O => \N__45282\,
            I => \N__45279\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__45279\,
            I => \c0.n22689\
        );

    \I__8433\ : InMux
    port map (
            O => \N__45276\,
            I => \N__45273\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__45273\,
            I => \N__45270\
        );

    \I__8431\ : Odrv4
    port map (
            O => \N__45270\,
            I => \c0.n22641\
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__45267\,
            I => \N__45264\
        );

    \I__8429\ : InMux
    port map (
            O => \N__45264\,
            I => \N__45257\
        );

    \I__8428\ : InMux
    port map (
            O => \N__45263\,
            I => \N__45254\
        );

    \I__8427\ : InMux
    port map (
            O => \N__45262\,
            I => \N__45251\
        );

    \I__8426\ : InMux
    port map (
            O => \N__45261\,
            I => \N__45248\
        );

    \I__8425\ : InMux
    port map (
            O => \N__45260\,
            I => \N__45245\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__45257\,
            I => \N__45242\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__45254\,
            I => \N__45239\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__45251\,
            I => \N__45236\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__45248\,
            I => \N__45233\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__45245\,
            I => \N__45230\
        );

    \I__8419\ : Span4Mux_v
    port map (
            O => \N__45242\,
            I => \N__45219\
        );

    \I__8418\ : Span4Mux_v
    port map (
            O => \N__45239\,
            I => \N__45219\
        );

    \I__8417\ : Span4Mux_h
    port map (
            O => \N__45236\,
            I => \N__45219\
        );

    \I__8416\ : Span4Mux_v
    port map (
            O => \N__45233\,
            I => \N__45219\
        );

    \I__8415\ : Span4Mux_v
    port map (
            O => \N__45230\,
            I => \N__45216\
        );

    \I__8414\ : InMux
    port map (
            O => \N__45229\,
            I => \N__45213\
        );

    \I__8413\ : InMux
    port map (
            O => \N__45228\,
            I => \N__45210\
        );

    \I__8412\ : Span4Mux_h
    port map (
            O => \N__45219\,
            I => \N__45207\
        );

    \I__8411\ : Span4Mux_h
    port map (
            O => \N__45216\,
            I => \N__45204\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__45213\,
            I => \N__45201\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__45210\,
            I => encoder0_position_4
        );

    \I__8408\ : Odrv4
    port map (
            O => \N__45207\,
            I => encoder0_position_4
        );

    \I__8407\ : Odrv4
    port map (
            O => \N__45204\,
            I => encoder0_position_4
        );

    \I__8406\ : Odrv4
    port map (
            O => \N__45201\,
            I => encoder0_position_4
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__45192\,
            I => \c0.n22689_cascade_\
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__45189\,
            I => \N__45186\
        );

    \I__8403\ : InMux
    port map (
            O => \N__45186\,
            I => \N__45181\
        );

    \I__8402\ : InMux
    port map (
            O => \N__45185\,
            I => \N__45178\
        );

    \I__8401\ : InMux
    port map (
            O => \N__45184\,
            I => \N__45175\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__45181\,
            I => \N__45170\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__45178\,
            I => \N__45165\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__45175\,
            I => \N__45165\
        );

    \I__8397\ : InMux
    port map (
            O => \N__45174\,
            I => \N__45162\
        );

    \I__8396\ : InMux
    port map (
            O => \N__45173\,
            I => \N__45159\
        );

    \I__8395\ : Span4Mux_h
    port map (
            O => \N__45170\,
            I => \N__45155\
        );

    \I__8394\ : Span4Mux_v
    port map (
            O => \N__45165\,
            I => \N__45152\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45149\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__45159\,
            I => \N__45146\
        );

    \I__8391\ : InMux
    port map (
            O => \N__45158\,
            I => \N__45143\
        );

    \I__8390\ : Span4Mux_h
    port map (
            O => \N__45155\,
            I => \N__45140\
        );

    \I__8389\ : Span4Mux_v
    port map (
            O => \N__45152\,
            I => \N__45137\
        );

    \I__8388\ : Span12Mux_h
    port map (
            O => \N__45149\,
            I => \N__45132\
        );

    \I__8387\ : Span12Mux_v
    port map (
            O => \N__45146\,
            I => \N__45132\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__45143\,
            I => control_mode_0
        );

    \I__8385\ : Odrv4
    port map (
            O => \N__45140\,
            I => control_mode_0
        );

    \I__8384\ : Odrv4
    port map (
            O => \N__45137\,
            I => control_mode_0
        );

    \I__8383\ : Odrv12
    port map (
            O => \N__45132\,
            I => control_mode_0
        );

    \I__8382\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45120\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__45120\,
            I => \N__45117\
        );

    \I__8380\ : Span4Mux_h
    port map (
            O => \N__45117\,
            I => \N__45113\
        );

    \I__8379\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45110\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__45113\,
            I => \c0.n10455\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__45110\,
            I => \c0.n10455\
        );

    \I__8376\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45102\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__45102\,
            I => \N__45099\
        );

    \I__8374\ : Span4Mux_h
    port map (
            O => \N__45099\,
            I => \N__45095\
        );

    \I__8373\ : InMux
    port map (
            O => \N__45098\,
            I => \N__45092\
        );

    \I__8372\ : Odrv4
    port map (
            O => \N__45095\,
            I => \c0.n20312\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__45092\,
            I => \c0.n20312\
        );

    \I__8370\ : CascadeMux
    port map (
            O => \N__45087\,
            I => \c0.n20312_cascade_\
        );

    \I__8369\ : InMux
    port map (
            O => \N__45084\,
            I => \N__45081\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__45081\,
            I => \c0.n22522\
        );

    \I__8367\ : CascadeMux
    port map (
            O => \N__45078\,
            I => \c0.n6_adj_4674_cascade_\
        );

    \I__8366\ : InMux
    port map (
            O => \N__45075\,
            I => \N__45072\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__45072\,
            I => \N__45069\
        );

    \I__8364\ : Span4Mux_h
    port map (
            O => \N__45069\,
            I => \N__45066\
        );

    \I__8363\ : Span4Mux_h
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__8362\ : Odrv4
    port map (
            O => \N__45063\,
            I => \c0.data_out_frame_29_4\
        );

    \I__8361\ : CEMux
    port map (
            O => \N__45060\,
            I => \N__45056\
        );

    \I__8360\ : CEMux
    port map (
            O => \N__45059\,
            I => \N__45051\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__45056\,
            I => \N__45047\
        );

    \I__8358\ : CEMux
    port map (
            O => \N__45055\,
            I => \N__45044\
        );

    \I__8357\ : CEMux
    port map (
            O => \N__45054\,
            I => \N__45038\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__45051\,
            I => \N__45032\
        );

    \I__8355\ : CEMux
    port map (
            O => \N__45050\,
            I => \N__45029\
        );

    \I__8354\ : Span4Mux_h
    port map (
            O => \N__45047\,
            I => \N__45022\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__45044\,
            I => \N__45022\
        );

    \I__8352\ : CEMux
    port map (
            O => \N__45043\,
            I => \N__45019\
        );

    \I__8351\ : CEMux
    port map (
            O => \N__45042\,
            I => \N__45016\
        );

    \I__8350\ : CEMux
    port map (
            O => \N__45041\,
            I => \N__45013\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__45038\,
            I => \N__45010\
        );

    \I__8348\ : CEMux
    port map (
            O => \N__45037\,
            I => \N__45007\
        );

    \I__8347\ : CEMux
    port map (
            O => \N__45036\,
            I => \N__45004\
        );

    \I__8346\ : CEMux
    port map (
            O => \N__45035\,
            I => \N__45001\
        );

    \I__8345\ : Span4Mux_v
    port map (
            O => \N__45032\,
            I => \N__44996\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__45029\,
            I => \N__44996\
        );

    \I__8343\ : SRMux
    port map (
            O => \N__45028\,
            I => \N__44992\
        );

    \I__8342\ : SRMux
    port map (
            O => \N__45027\,
            I => \N__44989\
        );

    \I__8341\ : Span4Mux_h
    port map (
            O => \N__45022\,
            I => \N__44986\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__45019\,
            I => \N__44983\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__45016\,
            I => \N__44980\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__45013\,
            I => \N__44975\
        );

    \I__8337\ : Span4Mux_h
    port map (
            O => \N__45010\,
            I => \N__44975\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__45007\,
            I => \N__44972\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__45004\,
            I => \N__44967\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__45001\,
            I => \N__44967\
        );

    \I__8333\ : Span4Mux_h
    port map (
            O => \N__44996\,
            I => \N__44964\
        );

    \I__8332\ : SRMux
    port map (
            O => \N__44995\,
            I => \N__44961\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__44992\,
            I => \N__44956\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__44989\,
            I => \N__44956\
        );

    \I__8329\ : Span4Mux_v
    port map (
            O => \N__44986\,
            I => \N__44953\
        );

    \I__8328\ : Span4Mux_v
    port map (
            O => \N__44983\,
            I => \N__44948\
        );

    \I__8327\ : Span4Mux_v
    port map (
            O => \N__44980\,
            I => \N__44948\
        );

    \I__8326\ : Span4Mux_v
    port map (
            O => \N__44975\,
            I => \N__44945\
        );

    \I__8325\ : Span4Mux_h
    port map (
            O => \N__44972\,
            I => \N__44938\
        );

    \I__8324\ : Span4Mux_h
    port map (
            O => \N__44967\,
            I => \N__44938\
        );

    \I__8323\ : Span4Mux_h
    port map (
            O => \N__44964\,
            I => \N__44938\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__44961\,
            I => \N__44931\
        );

    \I__8321\ : Span4Mux_v
    port map (
            O => \N__44956\,
            I => \N__44931\
        );

    \I__8320\ : Span4Mux_h
    port map (
            O => \N__44953\,
            I => \N__44931\
        );

    \I__8319\ : Span4Mux_v
    port map (
            O => \N__44948\,
            I => \N__44926\
        );

    \I__8318\ : Span4Mux_v
    port map (
            O => \N__44945\,
            I => \N__44926\
        );

    \I__8317\ : Sp12to4
    port map (
            O => \N__44938\,
            I => \N__44923\
        );

    \I__8316\ : Span4Mux_v
    port map (
            O => \N__44931\,
            I => \N__44920\
        );

    \I__8315\ : Span4Mux_h
    port map (
            O => \N__44926\,
            I => \N__44917\
        );

    \I__8314\ : Odrv12
    port map (
            O => \N__44923\,
            I => \c0.n8162\
        );

    \I__8313\ : Odrv4
    port map (
            O => \N__44920\,
            I => \c0.n8162\
        );

    \I__8312\ : Odrv4
    port map (
            O => \N__44917\,
            I => \c0.n8162\
        );

    \I__8311\ : InMux
    port map (
            O => \N__44910\,
            I => \N__44907\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__44907\,
            I => \N__44904\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__44904\,
            I => \c0.n22580\
        );

    \I__8308\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44896\
        );

    \I__8307\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44891\
        );

    \I__8306\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44891\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__44896\,
            I => \N__44888\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__44891\,
            I => \N__44883\
        );

    \I__8303\ : Span4Mux_h
    port map (
            O => \N__44888\,
            I => \N__44883\
        );

    \I__8302\ : Odrv4
    port map (
            O => \N__44883\,
            I => \c0.n10477\
        );

    \I__8301\ : InMux
    port map (
            O => \N__44880\,
            I => \N__44877\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__44877\,
            I => \N__44874\
        );

    \I__8299\ : Odrv4
    port map (
            O => \N__44874\,
            I => n2339
        );

    \I__8298\ : CascadeMux
    port map (
            O => \N__44871\,
            I => \N__44868\
        );

    \I__8297\ : InMux
    port map (
            O => \N__44868\,
            I => \N__44865\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__44865\,
            I => \N__44858\
        );

    \I__8295\ : InMux
    port map (
            O => \N__44864\,
            I => \N__44855\
        );

    \I__8294\ : CascadeMux
    port map (
            O => \N__44863\,
            I => \N__44852\
        );

    \I__8293\ : InMux
    port map (
            O => \N__44862\,
            I => \N__44847\
        );

    \I__8292\ : InMux
    port map (
            O => \N__44861\,
            I => \N__44847\
        );

    \I__8291\ : Span4Mux_h
    port map (
            O => \N__44858\,
            I => \N__44841\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__44855\,
            I => \N__44841\
        );

    \I__8289\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44838\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__44847\,
            I => \N__44835\
        );

    \I__8287\ : CascadeMux
    port map (
            O => \N__44846\,
            I => \N__44832\
        );

    \I__8286\ : Span4Mux_v
    port map (
            O => \N__44841\,
            I => \N__44827\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__44838\,
            I => \N__44822\
        );

    \I__8284\ : Span4Mux_v
    port map (
            O => \N__44835\,
            I => \N__44822\
        );

    \I__8283\ : InMux
    port map (
            O => \N__44832\,
            I => \N__44815\
        );

    \I__8282\ : InMux
    port map (
            O => \N__44831\,
            I => \N__44815\
        );

    \I__8281\ : InMux
    port map (
            O => \N__44830\,
            I => \N__44815\
        );

    \I__8280\ : Odrv4
    port map (
            O => \N__44827\,
            I => encoder0_position_18
        );

    \I__8279\ : Odrv4
    port map (
            O => \N__44822\,
            I => encoder0_position_18
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__44815\,
            I => encoder0_position_18
        );

    \I__8277\ : InMux
    port map (
            O => \N__44808\,
            I => \N__44805\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__44805\,
            I => \c0.n22583\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__44802\,
            I => \N__44799\
        );

    \I__8274\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44793\
        );

    \I__8273\ : InMux
    port map (
            O => \N__44798\,
            I => \N__44793\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__44793\,
            I => \N__44790\
        );

    \I__8271\ : Sp12to4
    port map (
            O => \N__44790\,
            I => \N__44787\
        );

    \I__8270\ : Span12Mux_s9_v
    port map (
            O => \N__44787\,
            I => \N__44784\
        );

    \I__8269\ : Odrv12
    port map (
            O => \N__44784\,
            I => \c0.n22149\
        );

    \I__8268\ : CascadeMux
    port map (
            O => \N__44781\,
            I => \N__44778\
        );

    \I__8267\ : InMux
    port map (
            O => \N__44778\,
            I => \N__44775\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__44775\,
            I => \N__44770\
        );

    \I__8265\ : InMux
    port map (
            O => \N__44774\,
            I => \N__44766\
        );

    \I__8264\ : InMux
    port map (
            O => \N__44773\,
            I => \N__44763\
        );

    \I__8263\ : Span4Mux_v
    port map (
            O => \N__44770\,
            I => \N__44759\
        );

    \I__8262\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44756\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__44766\,
            I => \N__44750\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__44763\,
            I => \N__44750\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__44762\,
            I => \N__44747\
        );

    \I__8258\ : Span4Mux_v
    port map (
            O => \N__44759\,
            I => \N__44744\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__44756\,
            I => \N__44741\
        );

    \I__8256\ : InMux
    port map (
            O => \N__44755\,
            I => \N__44738\
        );

    \I__8255\ : Span4Mux_v
    port map (
            O => \N__44750\,
            I => \N__44735\
        );

    \I__8254\ : InMux
    port map (
            O => \N__44747\,
            I => \N__44732\
        );

    \I__8253\ : Span4Mux_h
    port map (
            O => \N__44744\,
            I => \N__44727\
        );

    \I__8252\ : Span4Mux_v
    port map (
            O => \N__44741\,
            I => \N__44727\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__44738\,
            I => encoder0_position_3
        );

    \I__8250\ : Odrv4
    port map (
            O => \N__44735\,
            I => encoder0_position_3
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__44732\,
            I => encoder0_position_3
        );

    \I__8248\ : Odrv4
    port map (
            O => \N__44727\,
            I => encoder0_position_3
        );

    \I__8247\ : CascadeMux
    port map (
            O => \N__44718\,
            I => \c0.n22583_cascade_\
        );

    \I__8246\ : CascadeMux
    port map (
            O => \N__44715\,
            I => \N__44712\
        );

    \I__8245\ : InMux
    port map (
            O => \N__44712\,
            I => \N__44709\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__44709\,
            I => \N__44704\
        );

    \I__8243\ : InMux
    port map (
            O => \N__44708\,
            I => \N__44700\
        );

    \I__8242\ : InMux
    port map (
            O => \N__44707\,
            I => \N__44696\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__44704\,
            I => \N__44693\
        );

    \I__8240\ : InMux
    port map (
            O => \N__44703\,
            I => \N__44690\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__44700\,
            I => \N__44687\
        );

    \I__8238\ : InMux
    port map (
            O => \N__44699\,
            I => \N__44680\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__44696\,
            I => \N__44677\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__44693\,
            I => \N__44674\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__44690\,
            I => \N__44671\
        );

    \I__8234\ : Span4Mux_v
    port map (
            O => \N__44687\,
            I => \N__44668\
        );

    \I__8233\ : InMux
    port map (
            O => \N__44686\,
            I => \N__44665\
        );

    \I__8232\ : InMux
    port map (
            O => \N__44685\,
            I => \N__44660\
        );

    \I__8231\ : InMux
    port map (
            O => \N__44684\,
            I => \N__44660\
        );

    \I__8230\ : InMux
    port map (
            O => \N__44683\,
            I => \N__44657\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__44680\,
            I => \N__44652\
        );

    \I__8228\ : Span4Mux_h
    port map (
            O => \N__44677\,
            I => \N__44652\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__44674\,
            I => \N__44645\
        );

    \I__8226\ : Span4Mux_v
    port map (
            O => \N__44671\,
            I => \N__44645\
        );

    \I__8225\ : Span4Mux_v
    port map (
            O => \N__44668\,
            I => \N__44645\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__44665\,
            I => \N__44642\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__44660\,
            I => encoder0_position_31
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__44657\,
            I => encoder0_position_31
        );

    \I__8221\ : Odrv4
    port map (
            O => \N__44652\,
            I => encoder0_position_31
        );

    \I__8220\ : Odrv4
    port map (
            O => \N__44645\,
            I => encoder0_position_31
        );

    \I__8219\ : Odrv4
    port map (
            O => \N__44642\,
            I => encoder0_position_31
        );

    \I__8218\ : CascadeMux
    port map (
            O => \N__44631\,
            I => \N__44628\
        );

    \I__8217\ : InMux
    port map (
            O => \N__44628\,
            I => \N__44623\
        );

    \I__8216\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44618\
        );

    \I__8215\ : InMux
    port map (
            O => \N__44626\,
            I => \N__44618\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__44623\,
            I => \N__44613\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__44618\,
            I => \N__44613\
        );

    \I__8212\ : Span4Mux_h
    port map (
            O => \N__44613\,
            I => \N__44610\
        );

    \I__8211\ : Odrv4
    port map (
            O => \N__44610\,
            I => \c0.n13872\
        );

    \I__8210\ : CascadeMux
    port map (
            O => \N__44607\,
            I => \N__44604\
        );

    \I__8209\ : InMux
    port map (
            O => \N__44604\,
            I => \N__44601\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__44601\,
            I => \N__44598\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__44598\,
            I => \N__44595\
        );

    \I__8206\ : Span4Mux_v
    port map (
            O => \N__44595\,
            I => \N__44592\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__44592\,
            I => n2337
        );

    \I__8204\ : InMux
    port map (
            O => \N__44589\,
            I => \N__44585\
        );

    \I__8203\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44582\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__44585\,
            I => \N__44577\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__44582\,
            I => \N__44577\
        );

    \I__8200\ : Span4Mux_v
    port map (
            O => \N__44577\,
            I => \N__44574\
        );

    \I__8199\ : Span4Mux_v
    port map (
            O => \N__44574\,
            I => \N__44571\
        );

    \I__8198\ : Span4Mux_v
    port map (
            O => \N__44571\,
            I => \N__44568\
        );

    \I__8197\ : Odrv4
    port map (
            O => \N__44568\,
            I => n17571
        );

    \I__8196\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44562\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__44562\,
            I => \N__44559\
        );

    \I__8194\ : Span4Mux_h
    port map (
            O => \N__44559\,
            I => \N__44554\
        );

    \I__8193\ : InMux
    port map (
            O => \N__44558\,
            I => \N__44549\
        );

    \I__8192\ : InMux
    port map (
            O => \N__44557\,
            I => \N__44549\
        );

    \I__8191\ : Sp12to4
    port map (
            O => \N__44554\,
            I => \N__44545\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__44549\,
            I => \N__44542\
        );

    \I__8189\ : InMux
    port map (
            O => \N__44548\,
            I => \N__44539\
        );

    \I__8188\ : Span12Mux_v
    port map (
            O => \N__44545\,
            I => \N__44536\
        );

    \I__8187\ : Span4Mux_h
    port map (
            O => \N__44542\,
            I => \N__44533\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__44539\,
            I => data_in_1_6
        );

    \I__8185\ : Odrv12
    port map (
            O => \N__44536\,
            I => data_in_1_6
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__44533\,
            I => data_in_1_6
        );

    \I__8183\ : InMux
    port map (
            O => \N__44526\,
            I => \N__44522\
        );

    \I__8182\ : InMux
    port map (
            O => \N__44525\,
            I => \N__44519\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__44522\,
            I => \N__44514\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__44519\,
            I => \N__44514\
        );

    \I__8179\ : Span4Mux_v
    port map (
            O => \N__44514\,
            I => \N__44510\
        );

    \I__8178\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44507\
        );

    \I__8177\ : Span4Mux_v
    port map (
            O => \N__44510\,
            I => \N__44504\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__44507\,
            I => data_in_0_6
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__44504\,
            I => data_in_0_6
        );

    \I__8174\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44496\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__44496\,
            I => \N__44493\
        );

    \I__8172\ : Span4Mux_v
    port map (
            O => \N__44493\,
            I => \N__44489\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__44492\,
            I => \N__44486\
        );

    \I__8170\ : Span4Mux_h
    port map (
            O => \N__44489\,
            I => \N__44482\
        );

    \I__8169\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44479\
        );

    \I__8168\ : CascadeMux
    port map (
            O => \N__44485\,
            I => \N__44476\
        );

    \I__8167\ : Sp12to4
    port map (
            O => \N__44482\,
            I => \N__44473\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__44479\,
            I => \N__44470\
        );

    \I__8165\ : InMux
    port map (
            O => \N__44476\,
            I => \N__44467\
        );

    \I__8164\ : Span12Mux_h
    port map (
            O => \N__44473\,
            I => \N__44459\
        );

    \I__8163\ : Sp12to4
    port map (
            O => \N__44470\,
            I => \N__44459\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__44467\,
            I => \N__44459\
        );

    \I__8161\ : InMux
    port map (
            O => \N__44466\,
            I => \N__44456\
        );

    \I__8160\ : Span12Mux_v
    port map (
            O => \N__44459\,
            I => \N__44453\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__44456\,
            I => data_in_3_6
        );

    \I__8158\ : Odrv12
    port map (
            O => \N__44453\,
            I => data_in_3_6
        );

    \I__8157\ : CascadeMux
    port map (
            O => \N__44448\,
            I => \N__44445\
        );

    \I__8156\ : InMux
    port map (
            O => \N__44445\,
            I => \N__44442\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__44442\,
            I => \c0.n20_adj_4726\
        );

    \I__8154\ : InMux
    port map (
            O => \N__44439\,
            I => \N__44436\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__44436\,
            I => \c0.n27_adj_4735\
        );

    \I__8152\ : InMux
    port map (
            O => \N__44433\,
            I => \N__44429\
        );

    \I__8151\ : CascadeMux
    port map (
            O => \N__44432\,
            I => \N__44426\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__44429\,
            I => \N__44423\
        );

    \I__8149\ : InMux
    port map (
            O => \N__44426\,
            I => \N__44420\
        );

    \I__8148\ : Span4Mux_v
    port map (
            O => \N__44423\,
            I => \N__44417\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__44420\,
            I => \N__44414\
        );

    \I__8146\ : Odrv4
    port map (
            O => \N__44417\,
            I => \c0.data_out_frame_29__7__N_735\
        );

    \I__8145\ : Odrv12
    port map (
            O => \N__44414\,
            I => \c0.data_out_frame_29__7__N_735\
        );

    \I__8144\ : InMux
    port map (
            O => \N__44409\,
            I => \N__44406\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__44406\,
            I => \N__44402\
        );

    \I__8142\ : InMux
    port map (
            O => \N__44405\,
            I => \N__44399\
        );

    \I__8141\ : Span4Mux_h
    port map (
            O => \N__44402\,
            I => \N__44396\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__44399\,
            I => \N__44393\
        );

    \I__8139\ : Span4Mux_v
    port map (
            O => \N__44396\,
            I => \N__44390\
        );

    \I__8138\ : Span4Mux_v
    port map (
            O => \N__44393\,
            I => \N__44387\
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__44390\,
            I => \c0.n13665\
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__44387\,
            I => \c0.n13665\
        );

    \I__8135\ : InMux
    port map (
            O => \N__44382\,
            I => \N__44379\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__44379\,
            I => \N__44376\
        );

    \I__8133\ : Span4Mux_h
    port map (
            O => \N__44376\,
            I => \N__44373\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__44373\,
            I => \c0.n22754\
        );

    \I__8131\ : InMux
    port map (
            O => \N__44370\,
            I => \N__44367\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__44367\,
            I => \N__44364\
        );

    \I__8129\ : Span4Mux_h
    port map (
            O => \N__44364\,
            I => \N__44360\
        );

    \I__8128\ : InMux
    port map (
            O => \N__44363\,
            I => \N__44357\
        );

    \I__8127\ : Odrv4
    port map (
            O => \N__44360\,
            I => \c0.n13558\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__44357\,
            I => \c0.n13558\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__44352\,
            I => \c0.n22754_cascade_\
        );

    \I__8124\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44346\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__44346\,
            I => \N__44342\
        );

    \I__8122\ : InMux
    port map (
            O => \N__44345\,
            I => \N__44339\
        );

    \I__8121\ : Span4Mux_v
    port map (
            O => \N__44342\,
            I => \N__44336\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__44339\,
            I => \c0.n22243\
        );

    \I__8119\ : Odrv4
    port map (
            O => \N__44336\,
            I => \c0.n22243\
        );

    \I__8118\ : CascadeMux
    port map (
            O => \N__44331\,
            I => \N__44328\
        );

    \I__8117\ : InMux
    port map (
            O => \N__44328\,
            I => \N__44322\
        );

    \I__8116\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44315\
        );

    \I__8115\ : InMux
    port map (
            O => \N__44326\,
            I => \N__44315\
        );

    \I__8114\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44315\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__44322\,
            I => \N__44311\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__44315\,
            I => \N__44308\
        );

    \I__8111\ : InMux
    port map (
            O => \N__44314\,
            I => \N__44305\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__44311\,
            I => \N__44302\
        );

    \I__8109\ : Span4Mux_v
    port map (
            O => \N__44308\,
            I => \N__44299\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__44305\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__8107\ : Odrv4
    port map (
            O => \N__44302\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__44299\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__8105\ : SRMux
    port map (
            O => \N__44292\,
            I => \N__44289\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__44289\,
            I => \N__44286\
        );

    \I__8103\ : Span4Mux_h
    port map (
            O => \N__44286\,
            I => \N__44283\
        );

    \I__8102\ : Span4Mux_v
    port map (
            O => \N__44283\,
            I => \N__44280\
        );

    \I__8101\ : Odrv4
    port map (
            O => \N__44280\,
            I => \c0.n8_adj_4553\
        );

    \I__8100\ : InMux
    port map (
            O => \N__44277\,
            I => \N__44273\
        );

    \I__8099\ : InMux
    port map (
            O => \N__44276\,
            I => \N__44270\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__44273\,
            I => \N__44266\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__44270\,
            I => \N__44263\
        );

    \I__8096\ : InMux
    port map (
            O => \N__44269\,
            I => \N__44259\
        );

    \I__8095\ : Span4Mux_h
    port map (
            O => \N__44266\,
            I => \N__44256\
        );

    \I__8094\ : Span4Mux_v
    port map (
            O => \N__44263\,
            I => \N__44253\
        );

    \I__8093\ : InMux
    port map (
            O => \N__44262\,
            I => \N__44250\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__44259\,
            I => \N__44247\
        );

    \I__8091\ : Odrv4
    port map (
            O => \N__44256\,
            I => \c0.n4_adj_4212\
        );

    \I__8090\ : Odrv4
    port map (
            O => \N__44253\,
            I => \c0.n4_adj_4212\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__44250\,
            I => \c0.n4_adj_4212\
        );

    \I__8088\ : Odrv12
    port map (
            O => \N__44247\,
            I => \c0.n4_adj_4212\
        );

    \I__8087\ : CascadeMux
    port map (
            O => \N__44238\,
            I => \c0.n22098_cascade_\
        );

    \I__8086\ : InMux
    port map (
            O => \N__44235\,
            I => \N__44232\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__44232\,
            I => \c0.n4_adj_4306\
        );

    \I__8084\ : CascadeMux
    port map (
            O => \N__44229\,
            I => \c0.n63_adj_4305_cascade_\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__44226\,
            I => \N__44222\
        );

    \I__8082\ : InMux
    port map (
            O => \N__44225\,
            I => \N__44214\
        );

    \I__8081\ : InMux
    port map (
            O => \N__44222\,
            I => \N__44205\
        );

    \I__8080\ : InMux
    port map (
            O => \N__44221\,
            I => \N__44205\
        );

    \I__8079\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44205\
        );

    \I__8078\ : InMux
    port map (
            O => \N__44219\,
            I => \N__44205\
        );

    \I__8077\ : CascadeMux
    port map (
            O => \N__44218\,
            I => \N__44202\
        );

    \I__8076\ : CascadeMux
    port map (
            O => \N__44217\,
            I => \N__44198\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__44214\,
            I => \N__44191\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__44205\,
            I => \N__44188\
        );

    \I__8073\ : InMux
    port map (
            O => \N__44202\,
            I => \N__44179\
        );

    \I__8072\ : InMux
    port map (
            O => \N__44201\,
            I => \N__44179\
        );

    \I__8071\ : InMux
    port map (
            O => \N__44198\,
            I => \N__44179\
        );

    \I__8070\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44179\
        );

    \I__8069\ : InMux
    port map (
            O => \N__44196\,
            I => \N__44176\
        );

    \I__8068\ : InMux
    port map (
            O => \N__44195\,
            I => \N__44173\
        );

    \I__8067\ : InMux
    port map (
            O => \N__44194\,
            I => \N__44170\
        );

    \I__8066\ : Span4Mux_v
    port map (
            O => \N__44191\,
            I => \N__44159\
        );

    \I__8065\ : Span4Mux_h
    port map (
            O => \N__44188\,
            I => \N__44159\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__44179\,
            I => \N__44159\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__44176\,
            I => \N__44159\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__44173\,
            I => \N__44159\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__44170\,
            I => \N__44155\
        );

    \I__8060\ : Span4Mux_h
    port map (
            O => \N__44159\,
            I => \N__44152\
        );

    \I__8059\ : InMux
    port map (
            O => \N__44158\,
            I => \N__44149\
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__44155\,
            I => \c0.n13001\
        );

    \I__8057\ : Odrv4
    port map (
            O => \N__44152\,
            I => \c0.n13001\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__44149\,
            I => \c0.n13001\
        );

    \I__8055\ : CascadeMux
    port map (
            O => \N__44142\,
            I => \N__44138\
        );

    \I__8054\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44135\
        );

    \I__8053\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44132\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__44135\,
            I => \N__44128\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__44132\,
            I => \N__44125\
        );

    \I__8050\ : InMux
    port map (
            O => \N__44131\,
            I => \N__44122\
        );

    \I__8049\ : Span4Mux_h
    port map (
            O => \N__44128\,
            I => \N__44119\
        );

    \I__8048\ : Span4Mux_h
    port map (
            O => \N__44125\,
            I => \N__44116\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__44122\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__8046\ : Odrv4
    port map (
            O => \N__44119\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__8045\ : Odrv4
    port map (
            O => \N__44116\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__8044\ : InMux
    port map (
            O => \N__44109\,
            I => \N__44105\
        );

    \I__8043\ : InMux
    port map (
            O => \N__44108\,
            I => \N__44100\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__44105\,
            I => \N__44097\
        );

    \I__8041\ : InMux
    port map (
            O => \N__44104\,
            I => \N__44094\
        );

    \I__8040\ : InMux
    port map (
            O => \N__44103\,
            I => \N__44091\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__44100\,
            I => \N__44088\
        );

    \I__8038\ : Span4Mux_v
    port map (
            O => \N__44097\,
            I => \N__44079\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__44094\,
            I => \N__44079\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__44091\,
            I => \N__44079\
        );

    \I__8035\ : Span4Mux_h
    port map (
            O => \N__44088\,
            I => \N__44076\
        );

    \I__8034\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44073\
        );

    \I__8033\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44070\
        );

    \I__8032\ : Span4Mux_h
    port map (
            O => \N__44079\,
            I => \N__44067\
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__44076\,
            I => \c0.n9248\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__44073\,
            I => \c0.n9248\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__44070\,
            I => \c0.n9248\
        );

    \I__8028\ : Odrv4
    port map (
            O => \N__44067\,
            I => \c0.n9248\
        );

    \I__8027\ : InMux
    port map (
            O => \N__44058\,
            I => \N__44053\
        );

    \I__8026\ : InMux
    port map (
            O => \N__44057\,
            I => \N__44050\
        );

    \I__8025\ : InMux
    port map (
            O => \N__44056\,
            I => \N__44047\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__44053\,
            I => \N__44040\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__44050\,
            I => \N__44040\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__44047\,
            I => \N__44037\
        );

    \I__8021\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44034\
        );

    \I__8020\ : InMux
    port map (
            O => \N__44045\,
            I => \N__44031\
        );

    \I__8019\ : Span4Mux_h
    port map (
            O => \N__44040\,
            I => \N__44028\
        );

    \I__8018\ : Span4Mux_h
    port map (
            O => \N__44037\,
            I => \N__44025\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__44034\,
            I => \N__44022\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__44031\,
            I => \c0.n13055\
        );

    \I__8015\ : Odrv4
    port map (
            O => \N__44028\,
            I => \c0.n13055\
        );

    \I__8014\ : Odrv4
    port map (
            O => \N__44025\,
            I => \c0.n13055\
        );

    \I__8013\ : Odrv4
    port map (
            O => \N__44022\,
            I => \c0.n13055\
        );

    \I__8012\ : InMux
    port map (
            O => \N__44013\,
            I => \N__44008\
        );

    \I__8011\ : CascadeMux
    port map (
            O => \N__44012\,
            I => \N__44005\
        );

    \I__8010\ : CascadeMux
    port map (
            O => \N__44011\,
            I => \N__43999\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__44008\,
            I => \N__43994\
        );

    \I__8008\ : InMux
    port map (
            O => \N__44005\,
            I => \N__43991\
        );

    \I__8007\ : InMux
    port map (
            O => \N__44004\,
            I => \N__43986\
        );

    \I__8006\ : InMux
    port map (
            O => \N__44003\,
            I => \N__43986\
        );

    \I__8005\ : InMux
    port map (
            O => \N__44002\,
            I => \N__43983\
        );

    \I__8004\ : InMux
    port map (
            O => \N__43999\,
            I => \N__43980\
        );

    \I__8003\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43977\
        );

    \I__8002\ : CascadeMux
    port map (
            O => \N__43997\,
            I => \N__43974\
        );

    \I__8001\ : Span4Mux_v
    port map (
            O => \N__43994\,
            I => \N__43969\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__43991\,
            I => \N__43969\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__43986\,
            I => \N__43964\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__43983\,
            I => \N__43959\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__43980\,
            I => \N__43959\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__43977\,
            I => \N__43956\
        );

    \I__7995\ : InMux
    port map (
            O => \N__43974\,
            I => \N__43953\
        );

    \I__7994\ : Span4Mux_h
    port map (
            O => \N__43969\,
            I => \N__43950\
        );

    \I__7993\ : InMux
    port map (
            O => \N__43968\,
            I => \N__43947\
        );

    \I__7992\ : InMux
    port map (
            O => \N__43967\,
            I => \N__43944\
        );

    \I__7991\ : Span4Mux_v
    port map (
            O => \N__43964\,
            I => \N__43939\
        );

    \I__7990\ : Span4Mux_v
    port map (
            O => \N__43959\,
            I => \N__43939\
        );

    \I__7989\ : Odrv4
    port map (
            O => \N__43956\,
            I => \c0.data_out_frame_29_7_N_1482_0\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__43953\,
            I => \c0.data_out_frame_29_7_N_1482_0\
        );

    \I__7987\ : Odrv4
    port map (
            O => \N__43950\,
            I => \c0.data_out_frame_29_7_N_1482_0\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__43947\,
            I => \c0.data_out_frame_29_7_N_1482_0\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__43944\,
            I => \c0.data_out_frame_29_7_N_1482_0\
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__43939\,
            I => \c0.data_out_frame_29_7_N_1482_0\
        );

    \I__7983\ : InMux
    port map (
            O => \N__43926\,
            I => \N__43918\
        );

    \I__7982\ : InMux
    port map (
            O => \N__43925\,
            I => \N__43918\
        );

    \I__7981\ : InMux
    port map (
            O => \N__43924\,
            I => \N__43915\
        );

    \I__7980\ : InMux
    port map (
            O => \N__43923\,
            I => \N__43912\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__43918\,
            I => \N__43908\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__43915\,
            I => \N__43905\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__43912\,
            I => \N__43902\
        );

    \I__7976\ : InMux
    port map (
            O => \N__43911\,
            I => \N__43896\
        );

    \I__7975\ : Span4Mux_h
    port map (
            O => \N__43908\,
            I => \N__43891\
        );

    \I__7974\ : Span4Mux_v
    port map (
            O => \N__43905\,
            I => \N__43891\
        );

    \I__7973\ : Span4Mux_h
    port map (
            O => \N__43902\,
            I => \N__43888\
        );

    \I__7972\ : InMux
    port map (
            O => \N__43901\,
            I => \N__43885\
        );

    \I__7971\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43880\
        );

    \I__7970\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43880\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__43896\,
            I => \data_out_frame_29_7_N_2878_2\
        );

    \I__7968\ : Odrv4
    port map (
            O => \N__43891\,
            I => \data_out_frame_29_7_N_2878_2\
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__43888\,
            I => \data_out_frame_29_7_N_2878_2\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__43885\,
            I => \data_out_frame_29_7_N_2878_2\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__43880\,
            I => \data_out_frame_29_7_N_2878_2\
        );

    \I__7964\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43866\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43862\
        );

    \I__7962\ : InMux
    port map (
            O => \N__43865\,
            I => \N__43859\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__43862\,
            I => \N__43856\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__43859\,
            I => \N__43853\
        );

    \I__7959\ : Span4Mux_h
    port map (
            O => \N__43856\,
            I => \N__43850\
        );

    \I__7958\ : Span4Mux_v
    port map (
            O => \N__43853\,
            I => \N__43847\
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__43850\,
            I => \c0.n9_adj_4549\
        );

    \I__7956\ : Odrv4
    port map (
            O => \N__43847\,
            I => \c0.n9_adj_4549\
        );

    \I__7955\ : CascadeMux
    port map (
            O => \N__43842\,
            I => \N__43839\
        );

    \I__7954\ : InMux
    port map (
            O => \N__43839\,
            I => \N__43831\
        );

    \I__7953\ : CascadeMux
    port map (
            O => \N__43838\,
            I => \N__43826\
        );

    \I__7952\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43821\
        );

    \I__7951\ : InMux
    port map (
            O => \N__43836\,
            I => \N__43817\
        );

    \I__7950\ : CascadeMux
    port map (
            O => \N__43835\,
            I => \N__43813\
        );

    \I__7949\ : CascadeMux
    port map (
            O => \N__43834\,
            I => \N__43810\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__43831\,
            I => \N__43806\
        );

    \I__7947\ : InMux
    port map (
            O => \N__43830\,
            I => \N__43803\
        );

    \I__7946\ : InMux
    port map (
            O => \N__43829\,
            I => \N__43800\
        );

    \I__7945\ : InMux
    port map (
            O => \N__43826\,
            I => \N__43797\
        );

    \I__7944\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43793\
        );

    \I__7943\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43790\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__43821\,
            I => \N__43787\
        );

    \I__7941\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43784\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__43817\,
            I => \N__43781\
        );

    \I__7939\ : InMux
    port map (
            O => \N__43816\,
            I => \N__43778\
        );

    \I__7938\ : InMux
    port map (
            O => \N__43813\,
            I => \N__43773\
        );

    \I__7937\ : InMux
    port map (
            O => \N__43810\,
            I => \N__43773\
        );

    \I__7936\ : InMux
    port map (
            O => \N__43809\,
            I => \N__43770\
        );

    \I__7935\ : Span4Mux_v
    port map (
            O => \N__43806\,
            I => \N__43765\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__43803\,
            I => \N__43765\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__43800\,
            I => \N__43760\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__43797\,
            I => \N__43760\
        );

    \I__7931\ : InMux
    port map (
            O => \N__43796\,
            I => \N__43757\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__43793\,
            I => \N__43754\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__43790\,
            I => \N__43737\
        );

    \I__7928\ : Span4Mux_h
    port map (
            O => \N__43787\,
            I => \N__43737\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__43784\,
            I => \N__43737\
        );

    \I__7926\ : Span4Mux_v
    port map (
            O => \N__43781\,
            I => \N__43737\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__43778\,
            I => \N__43737\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__43773\,
            I => \N__43737\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__43770\,
            I => \N__43737\
        );

    \I__7922\ : Span4Mux_h
    port map (
            O => \N__43765\,
            I => \N__43734\
        );

    \I__7921\ : Span4Mux_h
    port map (
            O => \N__43760\,
            I => \N__43727\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__43757\,
            I => \N__43727\
        );

    \I__7919\ : Span4Mux_v
    port map (
            O => \N__43754\,
            I => \N__43727\
        );

    \I__7918\ : InMux
    port map (
            O => \N__43753\,
            I => \N__43722\
        );

    \I__7917\ : InMux
    port map (
            O => \N__43752\,
            I => \N__43722\
        );

    \I__7916\ : Span4Mux_v
    port map (
            O => \N__43737\,
            I => \N__43719\
        );

    \I__7915\ : Odrv4
    port map (
            O => \N__43734\,
            I => n63
        );

    \I__7914\ : Odrv4
    port map (
            O => \N__43727\,
            I => n63
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__43722\,
            I => n63
        );

    \I__7912\ : Odrv4
    port map (
            O => \N__43719\,
            I => n63
        );

    \I__7911\ : InMux
    port map (
            O => \N__43710\,
            I => \N__43705\
        );

    \I__7910\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43702\
        );

    \I__7909\ : CascadeMux
    port map (
            O => \N__43708\,
            I => \N__43699\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__43705\,
            I => \N__43693\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__43702\,
            I => \N__43693\
        );

    \I__7906\ : InMux
    port map (
            O => \N__43699\,
            I => \N__43690\
        );

    \I__7905\ : InMux
    port map (
            O => \N__43698\,
            I => \N__43687\
        );

    \I__7904\ : Span4Mux_v
    port map (
            O => \N__43693\,
            I => \N__43682\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__43690\,
            I => \N__43682\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__43687\,
            I => \N__43679\
        );

    \I__7901\ : Span4Mux_h
    port map (
            O => \N__43682\,
            I => \N__43676\
        );

    \I__7900\ : Odrv4
    port map (
            O => \N__43679\,
            I => \c0.n3844\
        );

    \I__7899\ : Odrv4
    port map (
            O => \N__43676\,
            I => \c0.n3844\
        );

    \I__7898\ : InMux
    port map (
            O => \N__43671\,
            I => \N__43668\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__43668\,
            I => \N__43664\
        );

    \I__7896\ : InMux
    port map (
            O => \N__43667\,
            I => \N__43661\
        );

    \I__7895\ : Span4Mux_v
    port map (
            O => \N__43664\,
            I => \N__43656\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__43661\,
            I => \N__43656\
        );

    \I__7893\ : Span4Mux_h
    port map (
            O => \N__43656\,
            I => \N__43651\
        );

    \I__7892\ : InMux
    port map (
            O => \N__43655\,
            I => \N__43648\
        );

    \I__7891\ : InMux
    port map (
            O => \N__43654\,
            I => \N__43645\
        );

    \I__7890\ : Odrv4
    port map (
            O => \N__43651\,
            I => \c0.n58_adj_4706\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__43648\,
            I => \c0.n58_adj_4706\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__43645\,
            I => \c0.n58_adj_4706\
        );

    \I__7887\ : CascadeMux
    port map (
            O => \N__43638\,
            I => \c0.n24591_cascade_\
        );

    \I__7886\ : InMux
    port map (
            O => \N__43635\,
            I => \N__43632\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__43632\,
            I => \N__43629\
        );

    \I__7884\ : Span4Mux_h
    port map (
            O => \N__43629\,
            I => \N__43626\
        );

    \I__7883\ : Odrv4
    port map (
            O => \N__43626\,
            I => \c0.n6_adj_4728\
        );

    \I__7882\ : InMux
    port map (
            O => \N__43623\,
            I => \N__43620\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__43620\,
            I => \N__43617\
        );

    \I__7880\ : Span12Mux_v
    port map (
            O => \N__43617\,
            I => \N__43614\
        );

    \I__7879\ : Odrv12
    port map (
            O => \N__43614\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__7878\ : InMux
    port map (
            O => \N__43611\,
            I => \N__43606\
        );

    \I__7877\ : InMux
    port map (
            O => \N__43610\,
            I => \N__43599\
        );

    \I__7876\ : InMux
    port map (
            O => \N__43609\,
            I => \N__43599\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__43606\,
            I => \N__43595\
        );

    \I__7874\ : InMux
    port map (
            O => \N__43605\,
            I => \N__43592\
        );

    \I__7873\ : InMux
    port map (
            O => \N__43604\,
            I => \N__43589\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__43599\,
            I => \N__43586\
        );

    \I__7871\ : InMux
    port map (
            O => \N__43598\,
            I => \N__43583\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__43595\,
            I => \N__43580\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__43592\,
            I => \N__43575\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__43589\,
            I => \N__43575\
        );

    \I__7867\ : Span4Mux_h
    port map (
            O => \N__43586\,
            I => \N__43572\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__43583\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__7865\ : Odrv4
    port map (
            O => \N__43580\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__7864\ : Odrv4
    port map (
            O => \N__43575\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__7863\ : Odrv4
    port map (
            O => \N__43572\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__7862\ : SRMux
    port map (
            O => \N__43563\,
            I => \N__43560\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__43560\,
            I => \N__43557\
        );

    \I__7860\ : Span12Mux_s9_v
    port map (
            O => \N__43557\,
            I => \N__43554\
        );

    \I__7859\ : Odrv12
    port map (
            O => \N__43554\,
            I => \c0.n21659\
        );

    \I__7858\ : InMux
    port map (
            O => \N__43551\,
            I => \N__43548\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__43548\,
            I => \c0.n4_adj_4721\
        );

    \I__7856\ : CascadeMux
    port map (
            O => \N__43545\,
            I => \N__43542\
        );

    \I__7855\ : InMux
    port map (
            O => \N__43542\,
            I => \N__43539\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__43539\,
            I => \N__43536\
        );

    \I__7853\ : Odrv12
    port map (
            O => \N__43536\,
            I => \c0.n937\
        );

    \I__7852\ : InMux
    port map (
            O => \N__43533\,
            I => \N__43527\
        );

    \I__7851\ : InMux
    port map (
            O => \N__43532\,
            I => \N__43523\
        );

    \I__7850\ : InMux
    port map (
            O => \N__43531\,
            I => \N__43520\
        );

    \I__7849\ : InMux
    port map (
            O => \N__43530\,
            I => \N__43517\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__43527\,
            I => \N__43510\
        );

    \I__7847\ : InMux
    port map (
            O => \N__43526\,
            I => \N__43507\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__43523\,
            I => \N__43500\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__43520\,
            I => \N__43500\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__43517\,
            I => \N__43500\
        );

    \I__7843\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43497\
        );

    \I__7842\ : InMux
    port map (
            O => \N__43515\,
            I => \N__43494\
        );

    \I__7841\ : InMux
    port map (
            O => \N__43514\,
            I => \N__43488\
        );

    \I__7840\ : InMux
    port map (
            O => \N__43513\,
            I => \N__43485\
        );

    \I__7839\ : Span4Mux_v
    port map (
            O => \N__43510\,
            I => \N__43478\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__43507\,
            I => \N__43478\
        );

    \I__7837\ : Span4Mux_v
    port map (
            O => \N__43500\,
            I => \N__43478\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__43497\,
            I => \N__43473\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__43494\,
            I => \N__43473\
        );

    \I__7834\ : InMux
    port map (
            O => \N__43493\,
            I => \N__43468\
        );

    \I__7833\ : InMux
    port map (
            O => \N__43492\,
            I => \N__43468\
        );

    \I__7832\ : InMux
    port map (
            O => \N__43491\,
            I => \N__43465\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__43488\,
            I => \c0.data_out_frame_29_7_N_1482_1\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__43485\,
            I => \c0.data_out_frame_29_7_N_1482_1\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__43478\,
            I => \c0.data_out_frame_29_7_N_1482_1\
        );

    \I__7828\ : Odrv4
    port map (
            O => \N__43473\,
            I => \c0.data_out_frame_29_7_N_1482_1\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__43468\,
            I => \c0.data_out_frame_29_7_N_1482_1\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__43465\,
            I => \c0.data_out_frame_29_7_N_1482_1\
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__43452\,
            I => \N__43449\
        );

    \I__7824\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43446\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__43446\,
            I => \N__43442\
        );

    \I__7822\ : InMux
    port map (
            O => \N__43445\,
            I => \N__43439\
        );

    \I__7821\ : Span4Mux_h
    port map (
            O => \N__43442\,
            I => \N__43436\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__43439\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__7819\ : Odrv4
    port map (
            O => \N__43436\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__7818\ : CascadeMux
    port map (
            O => \N__43431\,
            I => \N__43428\
        );

    \I__7817\ : InMux
    port map (
            O => \N__43428\,
            I => \N__43425\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__43425\,
            I => \N__43422\
        );

    \I__7815\ : Span4Mux_h
    port map (
            O => \N__43422\,
            I => \N__43419\
        );

    \I__7814\ : Odrv4
    port map (
            O => \N__43419\,
            I => \c0.n74_adj_4525\
        );

    \I__7813\ : InMux
    port map (
            O => \N__43416\,
            I => \N__43412\
        );

    \I__7812\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43409\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__43412\,
            I => \N__43403\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__43409\,
            I => \N__43403\
        );

    \I__7809\ : InMux
    port map (
            O => \N__43408\,
            I => \N__43400\
        );

    \I__7808\ : Span4Mux_h
    port map (
            O => \N__43403\,
            I => \N__43397\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__43400\,
            I => \N__43390\
        );

    \I__7806\ : Span4Mux_v
    port map (
            O => \N__43397\,
            I => \N__43390\
        );

    \I__7805\ : InMux
    port map (
            O => \N__43396\,
            I => \N__43387\
        );

    \I__7804\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43384\
        );

    \I__7803\ : Span4Mux_v
    port map (
            O => \N__43390\,
            I => \N__43381\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__43387\,
            I => \N__43378\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__43384\,
            I => control_mode_6
        );

    \I__7800\ : Odrv4
    port map (
            O => \N__43381\,
            I => control_mode_6
        );

    \I__7799\ : Odrv4
    port map (
            O => \N__43378\,
            I => control_mode_6
        );

    \I__7798\ : InMux
    port map (
            O => \N__43371\,
            I => \N__43368\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__43368\,
            I => \N__43364\
        );

    \I__7796\ : InMux
    port map (
            O => \N__43367\,
            I => \N__43360\
        );

    \I__7795\ : Span4Mux_v
    port map (
            O => \N__43364\,
            I => \N__43357\
        );

    \I__7794\ : InMux
    port map (
            O => \N__43363\,
            I => \N__43354\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__43360\,
            I => data_in_1_1
        );

    \I__7792\ : Odrv4
    port map (
            O => \N__43357\,
            I => data_in_1_1
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__43354\,
            I => data_in_1_1
        );

    \I__7790\ : InMux
    port map (
            O => \N__43347\,
            I => \N__43342\
        );

    \I__7789\ : InMux
    port map (
            O => \N__43346\,
            I => \N__43339\
        );

    \I__7788\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43336\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__43342\,
            I => data_in_0_1
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__43339\,
            I => data_in_0_1
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__43336\,
            I => data_in_0_1
        );

    \I__7784\ : InMux
    port map (
            O => \N__43329\,
            I => \N__43325\
        );

    \I__7783\ : CascadeMux
    port map (
            O => \N__43328\,
            I => \N__43322\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__43325\,
            I => \N__43319\
        );

    \I__7781\ : InMux
    port map (
            O => \N__43322\,
            I => \N__43314\
        );

    \I__7780\ : Span4Mux_h
    port map (
            O => \N__43319\,
            I => \N__43311\
        );

    \I__7779\ : InMux
    port map (
            O => \N__43318\,
            I => \N__43308\
        );

    \I__7778\ : InMux
    port map (
            O => \N__43317\,
            I => \N__43305\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__43314\,
            I => data_in_3_2
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__43311\,
            I => data_in_3_2
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__43308\,
            I => data_in_3_2
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__43305\,
            I => data_in_3_2
        );

    \I__7773\ : CascadeMux
    port map (
            O => \N__43296\,
            I => \N__43293\
        );

    \I__7772\ : InMux
    port map (
            O => \N__43293\,
            I => \N__43289\
        );

    \I__7771\ : InMux
    port map (
            O => \N__43292\,
            I => \N__43286\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__43289\,
            I => \N__43282\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__43286\,
            I => \N__43279\
        );

    \I__7768\ : InMux
    port map (
            O => \N__43285\,
            I => \N__43276\
        );

    \I__7767\ : Span4Mux_v
    port map (
            O => \N__43282\,
            I => \N__43271\
        );

    \I__7766\ : Span4Mux_v
    port map (
            O => \N__43279\,
            I => \N__43268\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__43276\,
            I => \N__43265\
        );

    \I__7764\ : InMux
    port map (
            O => \N__43275\,
            I => \N__43262\
        );

    \I__7763\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43259\
        );

    \I__7762\ : Span4Mux_v
    port map (
            O => \N__43271\,
            I => \N__43256\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__43268\,
            I => \N__43253\
        );

    \I__7760\ : Span12Mux_h
    port map (
            O => \N__43265\,
            I => \N__43248\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__43262\,
            I => \N__43248\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__43259\,
            I => control_mode_4
        );

    \I__7757\ : Odrv4
    port map (
            O => \N__43256\,
            I => control_mode_4
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__43253\,
            I => control_mode_4
        );

    \I__7755\ : Odrv12
    port map (
            O => \N__43248\,
            I => control_mode_4
        );

    \I__7754\ : InMux
    port map (
            O => \N__43239\,
            I => \N__43235\
        );

    \I__7753\ : InMux
    port map (
            O => \N__43238\,
            I => \N__43224\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__43235\,
            I => \N__43213\
        );

    \I__7751\ : InMux
    port map (
            O => \N__43234\,
            I => \N__43210\
        );

    \I__7750\ : InMux
    port map (
            O => \N__43233\,
            I => \N__43207\
        );

    \I__7749\ : InMux
    port map (
            O => \N__43232\,
            I => \N__43193\
        );

    \I__7748\ : InMux
    port map (
            O => \N__43231\,
            I => \N__43193\
        );

    \I__7747\ : InMux
    port map (
            O => \N__43230\,
            I => \N__43193\
        );

    \I__7746\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43193\
        );

    \I__7745\ : InMux
    port map (
            O => \N__43228\,
            I => \N__43193\
        );

    \I__7744\ : InMux
    port map (
            O => \N__43227\,
            I => \N__43193\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__43224\,
            I => \N__43190\
        );

    \I__7742\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43187\
        );

    \I__7741\ : InMux
    port map (
            O => \N__43222\,
            I => \N__43183\
        );

    \I__7740\ : InMux
    port map (
            O => \N__43221\,
            I => \N__43172\
        );

    \I__7739\ : InMux
    port map (
            O => \N__43220\,
            I => \N__43168\
        );

    \I__7738\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43165\
        );

    \I__7737\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43161\
        );

    \I__7736\ : InMux
    port map (
            O => \N__43217\,
            I => \N__43157\
        );

    \I__7735\ : InMux
    port map (
            O => \N__43216\,
            I => \N__43154\
        );

    \I__7734\ : Span4Mux_v
    port map (
            O => \N__43213\,
            I => \N__43149\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__43210\,
            I => \N__43149\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__43207\,
            I => \N__43146\
        );

    \I__7731\ : InMux
    port map (
            O => \N__43206\,
            I => \N__43143\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__43193\,
            I => \N__43138\
        );

    \I__7729\ : Span4Mux_v
    port map (
            O => \N__43190\,
            I => \N__43138\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__43187\,
            I => \N__43135\
        );

    \I__7727\ : InMux
    port map (
            O => \N__43186\,
            I => \N__43132\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__43183\,
            I => \N__43129\
        );

    \I__7725\ : InMux
    port map (
            O => \N__43182\,
            I => \N__43126\
        );

    \I__7724\ : InMux
    port map (
            O => \N__43181\,
            I => \N__43122\
        );

    \I__7723\ : InMux
    port map (
            O => \N__43180\,
            I => \N__43119\
        );

    \I__7722\ : InMux
    port map (
            O => \N__43179\,
            I => \N__43114\
        );

    \I__7721\ : InMux
    port map (
            O => \N__43178\,
            I => \N__43114\
        );

    \I__7720\ : InMux
    port map (
            O => \N__43177\,
            I => \N__43109\
        );

    \I__7719\ : InMux
    port map (
            O => \N__43176\,
            I => \N__43109\
        );

    \I__7718\ : InMux
    port map (
            O => \N__43175\,
            I => \N__43106\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__43172\,
            I => \N__43103\
        );

    \I__7716\ : InMux
    port map (
            O => \N__43171\,
            I => \N__43100\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__43168\,
            I => \N__43097\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__43165\,
            I => \N__43094\
        );

    \I__7713\ : InMux
    port map (
            O => \N__43164\,
            I => \N__43091\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__43161\,
            I => \N__43088\
        );

    \I__7711\ : InMux
    port map (
            O => \N__43160\,
            I => \N__43081\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__43157\,
            I => \N__43068\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__43154\,
            I => \N__43068\
        );

    \I__7708\ : Span4Mux_h
    port map (
            O => \N__43149\,
            I => \N__43068\
        );

    \I__7707\ : Span4Mux_v
    port map (
            O => \N__43146\,
            I => \N__43068\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__43143\,
            I => \N__43068\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__43138\,
            I => \N__43068\
        );

    \I__7704\ : Span4Mux_v
    port map (
            O => \N__43135\,
            I => \N__43063\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__43132\,
            I => \N__43063\
        );

    \I__7702\ : Span4Mux_v
    port map (
            O => \N__43129\,
            I => \N__43055\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__43126\,
            I => \N__43055\
        );

    \I__7700\ : InMux
    port map (
            O => \N__43125\,
            I => \N__43050\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__43122\,
            I => \N__43047\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__43119\,
            I => \N__43044\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__43114\,
            I => \N__43035\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__43109\,
            I => \N__43035\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__43106\,
            I => \N__43035\
        );

    \I__7694\ : Span4Mux_h
    port map (
            O => \N__43103\,
            I => \N__43035\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__43100\,
            I => \N__43029\
        );

    \I__7692\ : Span4Mux_h
    port map (
            O => \N__43097\,
            I => \N__43024\
        );

    \I__7691\ : Span4Mux_h
    port map (
            O => \N__43094\,
            I => \N__43024\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__43091\,
            I => \N__43021\
        );

    \I__7689\ : Span4Mux_v
    port map (
            O => \N__43088\,
            I => \N__43018\
        );

    \I__7688\ : InMux
    port map (
            O => \N__43087\,
            I => \N__43009\
        );

    \I__7687\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43009\
        );

    \I__7686\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43009\
        );

    \I__7685\ : InMux
    port map (
            O => \N__43084\,
            I => \N__43009\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__43081\,
            I => \N__43006\
        );

    \I__7683\ : Span4Mux_v
    port map (
            O => \N__43068\,
            I => \N__43001\
        );

    \I__7682\ : Span4Mux_v
    port map (
            O => \N__43063\,
            I => \N__43001\
        );

    \I__7681\ : InMux
    port map (
            O => \N__43062\,
            I => \N__42998\
        );

    \I__7680\ : InMux
    port map (
            O => \N__43061\,
            I => \N__42993\
        );

    \I__7679\ : InMux
    port map (
            O => \N__43060\,
            I => \N__42993\
        );

    \I__7678\ : Sp12to4
    port map (
            O => \N__43055\,
            I => \N__42990\
        );

    \I__7677\ : InMux
    port map (
            O => \N__43054\,
            I => \N__42987\
        );

    \I__7676\ : InMux
    port map (
            O => \N__43053\,
            I => \N__42984\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__43050\,
            I => \N__42979\
        );

    \I__7674\ : Span4Mux_h
    port map (
            O => \N__43047\,
            I => \N__42979\
        );

    \I__7673\ : Span4Mux_h
    port map (
            O => \N__43044\,
            I => \N__42974\
        );

    \I__7672\ : Span4Mux_h
    port map (
            O => \N__43035\,
            I => \N__42974\
        );

    \I__7671\ : InMux
    port map (
            O => \N__43034\,
            I => \N__42967\
        );

    \I__7670\ : InMux
    port map (
            O => \N__43033\,
            I => \N__42967\
        );

    \I__7669\ : InMux
    port map (
            O => \N__43032\,
            I => \N__42967\
        );

    \I__7668\ : Span4Mux_h
    port map (
            O => \N__43029\,
            I => \N__42960\
        );

    \I__7667\ : Span4Mux_v
    port map (
            O => \N__43024\,
            I => \N__42960\
        );

    \I__7666\ : Span4Mux_h
    port map (
            O => \N__43021\,
            I => \N__42960\
        );

    \I__7665\ : Span4Mux_v
    port map (
            O => \N__43018\,
            I => \N__42953\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__43009\,
            I => \N__42953\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__43006\,
            I => \N__42953\
        );

    \I__7662\ : Sp12to4
    port map (
            O => \N__43001\,
            I => \N__42948\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__42998\,
            I => \N__42948\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__42993\,
            I => \N__42943\
        );

    \I__7659\ : Span12Mux_h
    port map (
            O => \N__42990\,
            I => \N__42943\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__42987\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__42984\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7656\ : Odrv4
    port map (
            O => \N__42979\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7655\ : Odrv4
    port map (
            O => \N__42974\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__42967\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__42960\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7652\ : Odrv4
    port map (
            O => \N__42953\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7651\ : Odrv12
    port map (
            O => \N__42948\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7650\ : Odrv12
    port map (
            O => \N__42943\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7649\ : InMux
    port map (
            O => \N__42924\,
            I => \N__42920\
        );

    \I__7648\ : InMux
    port map (
            O => \N__42923\,
            I => \N__42917\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__42920\,
            I => \N__42914\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__42917\,
            I => data_out_frame_9_4
        );

    \I__7645\ : Odrv12
    port map (
            O => \N__42914\,
            I => data_out_frame_9_4
        );

    \I__7644\ : InMux
    port map (
            O => \N__42909\,
            I => \N__42906\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__42906\,
            I => \N__42902\
        );

    \I__7642\ : InMux
    port map (
            O => \N__42905\,
            I => \N__42899\
        );

    \I__7641\ : Span4Mux_v
    port map (
            O => \N__42902\,
            I => \N__42896\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__42899\,
            I => data_out_frame_8_4
        );

    \I__7639\ : Odrv4
    port map (
            O => \N__42896\,
            I => data_out_frame_8_4
        );

    \I__7638\ : InMux
    port map (
            O => \N__42891\,
            I => \N__42888\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__42888\,
            I => \N__42885\
        );

    \I__7636\ : Odrv4
    port map (
            O => \N__42885\,
            I => \c0.n24782\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__42882\,
            I => \N__42878\
        );

    \I__7634\ : CascadeMux
    port map (
            O => \N__42881\,
            I => \N__42875\
        );

    \I__7633\ : InMux
    port map (
            O => \N__42878\,
            I => \N__42872\
        );

    \I__7632\ : InMux
    port map (
            O => \N__42875\,
            I => \N__42869\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__42872\,
            I => \N__42866\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__42869\,
            I => \N__42863\
        );

    \I__7629\ : Span4Mux_v
    port map (
            O => \N__42866\,
            I => \N__42860\
        );

    \I__7628\ : Span4Mux_v
    port map (
            O => \N__42863\,
            I => \N__42857\
        );

    \I__7627\ : Span4Mux_h
    port map (
            O => \N__42860\,
            I => \N__42852\
        );

    \I__7626\ : Span4Mux_v
    port map (
            O => \N__42857\,
            I => \N__42849\
        );

    \I__7625\ : InMux
    port map (
            O => \N__42856\,
            I => \N__42846\
        );

    \I__7624\ : InMux
    port map (
            O => \N__42855\,
            I => \N__42842\
        );

    \I__7623\ : Sp12to4
    port map (
            O => \N__42852\,
            I => \N__42839\
        );

    \I__7622\ : Span4Mux_h
    port map (
            O => \N__42849\,
            I => \N__42834\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__42846\,
            I => \N__42834\
        );

    \I__7620\ : InMux
    port map (
            O => \N__42845\,
            I => \N__42831\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__42842\,
            I => encoder0_position_8
        );

    \I__7618\ : Odrv12
    port map (
            O => \N__42839\,
            I => encoder0_position_8
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__42834\,
            I => encoder0_position_8
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__42831\,
            I => encoder0_position_8
        );

    \I__7615\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42819\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__42819\,
            I => \N__42815\
        );

    \I__7613\ : InMux
    port map (
            O => \N__42818\,
            I => \N__42812\
        );

    \I__7612\ : Span4Mux_h
    port map (
            O => \N__42815\,
            I => \N__42809\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__42812\,
            I => \N__42806\
        );

    \I__7610\ : Span4Mux_v
    port map (
            O => \N__42809\,
            I => \N__42803\
        );

    \I__7609\ : Span4Mux_h
    port map (
            O => \N__42806\,
            I => \N__42800\
        );

    \I__7608\ : Span4Mux_v
    port map (
            O => \N__42803\,
            I => \N__42797\
        );

    \I__7607\ : Span4Mux_v
    port map (
            O => \N__42800\,
            I => \N__42794\
        );

    \I__7606\ : Odrv4
    port map (
            O => \N__42797\,
            I => \c0.n22423\
        );

    \I__7605\ : Odrv4
    port map (
            O => \N__42794\,
            I => \c0.n22423\
        );

    \I__7604\ : CascadeMux
    port map (
            O => \N__42789\,
            I => \N__42784\
        );

    \I__7603\ : CascadeMux
    port map (
            O => \N__42788\,
            I => \N__42781\
        );

    \I__7602\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42778\
        );

    \I__7601\ : InMux
    port map (
            O => \N__42784\,
            I => \N__42775\
        );

    \I__7600\ : InMux
    port map (
            O => \N__42781\,
            I => \N__42772\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__42778\,
            I => \N__42767\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__42775\,
            I => \N__42764\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__42772\,
            I => \N__42761\
        );

    \I__7596\ : InMux
    port map (
            O => \N__42771\,
            I => \N__42758\
        );

    \I__7595\ : InMux
    port map (
            O => \N__42770\,
            I => \N__42755\
        );

    \I__7594\ : Span4Mux_v
    port map (
            O => \N__42767\,
            I => \N__42752\
        );

    \I__7593\ : Span4Mux_v
    port map (
            O => \N__42764\,
            I => \N__42749\
        );

    \I__7592\ : Span4Mux_h
    port map (
            O => \N__42761\,
            I => \N__42746\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__42758\,
            I => \N__42743\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__42755\,
            I => \N__42738\
        );

    \I__7589\ : Span4Mux_v
    port map (
            O => \N__42752\,
            I => \N__42738\
        );

    \I__7588\ : Span4Mux_v
    port map (
            O => \N__42749\,
            I => \N__42733\
        );

    \I__7587\ : Span4Mux_h
    port map (
            O => \N__42746\,
            I => \N__42733\
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__42743\,
            I => encoder0_position_6
        );

    \I__7585\ : Odrv4
    port map (
            O => \N__42738\,
            I => encoder0_position_6
        );

    \I__7584\ : Odrv4
    port map (
            O => \N__42733\,
            I => encoder0_position_6
        );

    \I__7583\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42723\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__42723\,
            I => \c0.n6_adj_4293\
        );

    \I__7581\ : CascadeMux
    port map (
            O => \N__42720\,
            I => \N__42717\
        );

    \I__7580\ : InMux
    port map (
            O => \N__42717\,
            I => \N__42713\
        );

    \I__7579\ : CascadeMux
    port map (
            O => \N__42716\,
            I => \N__42710\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__42713\,
            I => \N__42707\
        );

    \I__7577\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42704\
        );

    \I__7576\ : Span4Mux_h
    port map (
            O => \N__42707\,
            I => \N__42698\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__42704\,
            I => \N__42695\
        );

    \I__7574\ : InMux
    port map (
            O => \N__42703\,
            I => \N__42692\
        );

    \I__7573\ : InMux
    port map (
            O => \N__42702\,
            I => \N__42689\
        );

    \I__7572\ : InMux
    port map (
            O => \N__42701\,
            I => \N__42685\
        );

    \I__7571\ : Span4Mux_h
    port map (
            O => \N__42698\,
            I => \N__42680\
        );

    \I__7570\ : Span4Mux_v
    port map (
            O => \N__42695\,
            I => \N__42680\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__42692\,
            I => \N__42675\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__42689\,
            I => \N__42675\
        );

    \I__7567\ : InMux
    port map (
            O => \N__42688\,
            I => \N__42672\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__42685\,
            I => encoder0_position_23
        );

    \I__7565\ : Odrv4
    port map (
            O => \N__42680\,
            I => encoder0_position_23
        );

    \I__7564\ : Odrv4
    port map (
            O => \N__42675\,
            I => encoder0_position_23
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__42672\,
            I => encoder0_position_23
        );

    \I__7562\ : InMux
    port map (
            O => \N__42663\,
            I => \N__42660\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__42660\,
            I => \N__42652\
        );

    \I__7560\ : InMux
    port map (
            O => \N__42659\,
            I => \N__42649\
        );

    \I__7559\ : InMux
    port map (
            O => \N__42658\,
            I => \N__42646\
        );

    \I__7558\ : InMux
    port map (
            O => \N__42657\,
            I => \N__42643\
        );

    \I__7557\ : InMux
    port map (
            O => \N__42656\,
            I => \N__42640\
        );

    \I__7556\ : InMux
    port map (
            O => \N__42655\,
            I => \N__42637\
        );

    \I__7555\ : Sp12to4
    port map (
            O => \N__42652\,
            I => \N__42632\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__42649\,
            I => \N__42632\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__42646\,
            I => \N__42629\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__42643\,
            I => encoder0_position_9
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__42640\,
            I => encoder0_position_9
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__42637\,
            I => encoder0_position_9
        );

    \I__7549\ : Odrv12
    port map (
            O => \N__42632\,
            I => encoder0_position_9
        );

    \I__7548\ : Odrv12
    port map (
            O => \N__42629\,
            I => encoder0_position_9
        );

    \I__7547\ : CascadeMux
    port map (
            O => \N__42618\,
            I => \N__42615\
        );

    \I__7546\ : InMux
    port map (
            O => \N__42615\,
            I => \N__42612\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__42612\,
            I => \N__42608\
        );

    \I__7544\ : CascadeMux
    port map (
            O => \N__42611\,
            I => \N__42605\
        );

    \I__7543\ : Span4Mux_v
    port map (
            O => \N__42608\,
            I => \N__42602\
        );

    \I__7542\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42598\
        );

    \I__7541\ : Span4Mux_h
    port map (
            O => \N__42602\,
            I => \N__42594\
        );

    \I__7540\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42591\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__42598\,
            I => \N__42588\
        );

    \I__7538\ : InMux
    port map (
            O => \N__42597\,
            I => \N__42585\
        );

    \I__7537\ : Span4Mux_h
    port map (
            O => \N__42594\,
            I => \N__42580\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__42591\,
            I => \N__42580\
        );

    \I__7535\ : Span12Mux_v
    port map (
            O => \N__42588\,
            I => \N__42577\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__42585\,
            I => control_mode_7
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__42580\,
            I => control_mode_7
        );

    \I__7532\ : Odrv12
    port map (
            O => \N__42577\,
            I => control_mode_7
        );

    \I__7531\ : CascadeMux
    port map (
            O => \N__42570\,
            I => \c0.n22385_cascade_\
        );

    \I__7530\ : CascadeMux
    port map (
            O => \N__42567\,
            I => \N__42564\
        );

    \I__7529\ : InMux
    port map (
            O => \N__42564\,
            I => \N__42561\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__42561\,
            I => \N__42556\
        );

    \I__7527\ : InMux
    port map (
            O => \N__42560\,
            I => \N__42553\
        );

    \I__7526\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42549\
        );

    \I__7525\ : Span4Mux_h
    port map (
            O => \N__42556\,
            I => \N__42544\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__42553\,
            I => \N__42544\
        );

    \I__7523\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42541\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__42549\,
            I => \N__42538\
        );

    \I__7521\ : Span4Mux_v
    port map (
            O => \N__42544\,
            I => \N__42532\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__42541\,
            I => \N__42529\
        );

    \I__7519\ : Span4Mux_h
    port map (
            O => \N__42538\,
            I => \N__42526\
        );

    \I__7518\ : InMux
    port map (
            O => \N__42537\,
            I => \N__42523\
        );

    \I__7517\ : InMux
    port map (
            O => \N__42536\,
            I => \N__42520\
        );

    \I__7516\ : InMux
    port map (
            O => \N__42535\,
            I => \N__42517\
        );

    \I__7515\ : Span4Mux_v
    port map (
            O => \N__42532\,
            I => \N__42514\
        );

    \I__7514\ : Span4Mux_h
    port map (
            O => \N__42529\,
            I => \N__42509\
        );

    \I__7513\ : Span4Mux_v
    port map (
            O => \N__42526\,
            I => \N__42509\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__42523\,
            I => encoder0_position_24
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__42520\,
            I => encoder0_position_24
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__42517\,
            I => encoder0_position_24
        );

    \I__7509\ : Odrv4
    port map (
            O => \N__42514\,
            I => encoder0_position_24
        );

    \I__7508\ : Odrv4
    port map (
            O => \N__42509\,
            I => encoder0_position_24
        );

    \I__7507\ : InMux
    port map (
            O => \N__42498\,
            I => \N__42494\
        );

    \I__7506\ : InMux
    port map (
            O => \N__42497\,
            I => \N__42491\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__42494\,
            I => \N__42488\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__42491\,
            I => \N__42485\
        );

    \I__7503\ : Span4Mux_h
    port map (
            O => \N__42488\,
            I => \N__42482\
        );

    \I__7502\ : Span4Mux_v
    port map (
            O => \N__42485\,
            I => \N__42479\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__42482\,
            I => \N__42474\
        );

    \I__7500\ : Span4Mux_h
    port map (
            O => \N__42479\,
            I => \N__42474\
        );

    \I__7499\ : Odrv4
    port map (
            O => \N__42474\,
            I => \c0.n20325\
        );

    \I__7498\ : InMux
    port map (
            O => \N__42471\,
            I => \N__42467\
        );

    \I__7497\ : CascadeMux
    port map (
            O => \N__42470\,
            I => \N__42463\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__42467\,
            I => \N__42459\
        );

    \I__7495\ : InMux
    port map (
            O => \N__42466\,
            I => \N__42454\
        );

    \I__7494\ : InMux
    port map (
            O => \N__42463\,
            I => \N__42454\
        );

    \I__7493\ : InMux
    port map (
            O => \N__42462\,
            I => \N__42451\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__42459\,
            I => \N__42448\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__42454\,
            I => \N__42445\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__42451\,
            I => data_in_2_5
        );

    \I__7489\ : Odrv4
    port map (
            O => \N__42448\,
            I => data_in_2_5
        );

    \I__7488\ : Odrv4
    port map (
            O => \N__42445\,
            I => data_in_2_5
        );

    \I__7487\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42431\
        );

    \I__7486\ : InMux
    port map (
            O => \N__42437\,
            I => \N__42431\
        );

    \I__7485\ : InMux
    port map (
            O => \N__42436\,
            I => \N__42428\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__42431\,
            I => \N__42424\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__42428\,
            I => \N__42421\
        );

    \I__7482\ : InMux
    port map (
            O => \N__42427\,
            I => \N__42418\
        );

    \I__7481\ : Span4Mux_h
    port map (
            O => \N__42424\,
            I => \N__42415\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__42421\,
            I => data_in_1_5
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__42418\,
            I => data_in_1_5
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__42415\,
            I => data_in_1_5
        );

    \I__7477\ : CascadeMux
    port map (
            O => \N__42408\,
            I => \N__42405\
        );

    \I__7476\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42402\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__42402\,
            I => \N__42397\
        );

    \I__7474\ : InMux
    port map (
            O => \N__42401\,
            I => \N__42394\
        );

    \I__7473\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42391\
        );

    \I__7472\ : Span4Mux_v
    port map (
            O => \N__42397\,
            I => \N__42382\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__42394\,
            I => \N__42382\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__42391\,
            I => \N__42382\
        );

    \I__7469\ : InMux
    port map (
            O => \N__42390\,
            I => \N__42377\
        );

    \I__7468\ : InMux
    port map (
            O => \N__42389\,
            I => \N__42374\
        );

    \I__7467\ : Span4Mux_h
    port map (
            O => \N__42382\,
            I => \N__42371\
        );

    \I__7466\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42366\
        );

    \I__7465\ : InMux
    port map (
            O => \N__42380\,
            I => \N__42366\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__42377\,
            I => \N__42363\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__42374\,
            I => encoder0_position_19
        );

    \I__7462\ : Odrv4
    port map (
            O => \N__42371\,
            I => encoder0_position_19
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__42366\,
            I => encoder0_position_19
        );

    \I__7460\ : Odrv12
    port map (
            O => \N__42363\,
            I => encoder0_position_19
        );

    \I__7459\ : CascadeMux
    port map (
            O => \N__42354\,
            I => \c0.n22199_cascade_\
        );

    \I__7458\ : InMux
    port map (
            O => \N__42351\,
            I => \N__42348\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__42348\,
            I => \N__42345\
        );

    \I__7456\ : Span4Mux_h
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__7455\ : Span4Mux_v
    port map (
            O => \N__42342\,
            I => \N__42338\
        );

    \I__7454\ : InMux
    port map (
            O => \N__42341\,
            I => \N__42335\
        );

    \I__7453\ : Odrv4
    port map (
            O => \N__42338\,
            I => \c0.n22834\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__42335\,
            I => \c0.n22834\
        );

    \I__7451\ : InMux
    port map (
            O => \N__42330\,
            I => \N__42325\
        );

    \I__7450\ : CascadeMux
    port map (
            O => \N__42329\,
            I => \N__42322\
        );

    \I__7449\ : InMux
    port map (
            O => \N__42328\,
            I => \N__42319\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__42325\,
            I => \N__42316\
        );

    \I__7447\ : InMux
    port map (
            O => \N__42322\,
            I => \N__42313\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__42319\,
            I => \N__42308\
        );

    \I__7445\ : Span4Mux_h
    port map (
            O => \N__42316\,
            I => \N__42308\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__42313\,
            I => \N__42304\
        );

    \I__7443\ : Span4Mux_v
    port map (
            O => \N__42308\,
            I => \N__42301\
        );

    \I__7442\ : InMux
    port map (
            O => \N__42307\,
            I => \N__42298\
        );

    \I__7441\ : Span4Mux_v
    port map (
            O => \N__42304\,
            I => \N__42292\
        );

    \I__7440\ : Span4Mux_v
    port map (
            O => \N__42301\,
            I => \N__42292\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__42298\,
            I => \N__42289\
        );

    \I__7438\ : InMux
    port map (
            O => \N__42297\,
            I => \N__42285\
        );

    \I__7437\ : Span4Mux_h
    port map (
            O => \N__42292\,
            I => \N__42282\
        );

    \I__7436\ : Sp12to4
    port map (
            O => \N__42289\,
            I => \N__42279\
        );

    \I__7435\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42276\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__42285\,
            I => encoder0_position_13
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__42282\,
            I => encoder0_position_13
        );

    \I__7432\ : Odrv12
    port map (
            O => \N__42279\,
            I => encoder0_position_13
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__42276\,
            I => encoder0_position_13
        );

    \I__7430\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42264\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__42264\,
            I => \N__42258\
        );

    \I__7428\ : InMux
    port map (
            O => \N__42263\,
            I => \N__42254\
        );

    \I__7427\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42251\
        );

    \I__7426\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42248\
        );

    \I__7425\ : Span4Mux_h
    port map (
            O => \N__42258\,
            I => \N__42244\
        );

    \I__7424\ : InMux
    port map (
            O => \N__42257\,
            I => \N__42241\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__42254\,
            I => \N__42238\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__42251\,
            I => \N__42235\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__42248\,
            I => \N__42232\
        );

    \I__7420\ : InMux
    port map (
            O => \N__42247\,
            I => \N__42229\
        );

    \I__7419\ : Span4Mux_v
    port map (
            O => \N__42244\,
            I => \N__42226\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__42241\,
            I => \N__42223\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__42238\,
            I => \N__42216\
        );

    \I__7416\ : Span4Mux_v
    port map (
            O => \N__42235\,
            I => \N__42216\
        );

    \I__7415\ : Span4Mux_v
    port map (
            O => \N__42232\,
            I => \N__42216\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__42229\,
            I => encoder0_position_22
        );

    \I__7413\ : Odrv4
    port map (
            O => \N__42226\,
            I => encoder0_position_22
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__42223\,
            I => encoder0_position_22
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__42216\,
            I => encoder0_position_22
        );

    \I__7410\ : InMux
    port map (
            O => \N__42207\,
            I => \N__42204\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__42204\,
            I => \c0.n6_adj_4366\
        );

    \I__7408\ : InMux
    port map (
            O => \N__42201\,
            I => \N__42195\
        );

    \I__7407\ : InMux
    port map (
            O => \N__42200\,
            I => \N__42195\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__42195\,
            I => \N__42190\
        );

    \I__7405\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42187\
        );

    \I__7404\ : InMux
    port map (
            O => \N__42193\,
            I => \N__42184\
        );

    \I__7403\ : Sp12to4
    port map (
            O => \N__42190\,
            I => \N__42181\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__42187\,
            I => data_in_2_0
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__42184\,
            I => data_in_2_0
        );

    \I__7400\ : Odrv12
    port map (
            O => \N__42181\,
            I => data_in_2_0
        );

    \I__7399\ : CascadeMux
    port map (
            O => \N__42174\,
            I => \N__42171\
        );

    \I__7398\ : InMux
    port map (
            O => \N__42171\,
            I => \N__42167\
        );

    \I__7397\ : InMux
    port map (
            O => \N__42170\,
            I => \N__42164\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__42167\,
            I => \N__42161\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__42164\,
            I => \N__42158\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__42161\,
            I => \N__42155\
        );

    \I__7393\ : Odrv12
    port map (
            O => \N__42158\,
            I => \c0.n22635\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__42155\,
            I => \c0.n22635\
        );

    \I__7391\ : CascadeMux
    port map (
            O => \N__42150\,
            I => \c0.n22256_cascade_\
        );

    \I__7390\ : InMux
    port map (
            O => \N__42147\,
            I => \N__42144\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__42144\,
            I => \N__42140\
        );

    \I__7388\ : InMux
    port map (
            O => \N__42143\,
            I => \N__42137\
        );

    \I__7387\ : Span4Mux_v
    port map (
            O => \N__42140\,
            I => \N__42134\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__42137\,
            I => \N__42131\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__42134\,
            I => \N__42128\
        );

    \I__7384\ : Odrv12
    port map (
            O => \N__42131\,
            I => \c0.n22772\
        );

    \I__7383\ : Odrv4
    port map (
            O => \N__42128\,
            I => \c0.n22772\
        );

    \I__7382\ : InMux
    port map (
            O => \N__42123\,
            I => \N__42118\
        );

    \I__7381\ : CascadeMux
    port map (
            O => \N__42122\,
            I => \N__42115\
        );

    \I__7380\ : InMux
    port map (
            O => \N__42121\,
            I => \N__42111\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__42118\,
            I => \N__42108\
        );

    \I__7378\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42105\
        );

    \I__7377\ : InMux
    port map (
            O => \N__42114\,
            I => \N__42102\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__42111\,
            I => data_in_1_3
        );

    \I__7375\ : Odrv4
    port map (
            O => \N__42108\,
            I => data_in_1_3
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__42105\,
            I => data_in_1_3
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__42102\,
            I => data_in_1_3
        );

    \I__7372\ : InMux
    port map (
            O => \N__42093\,
            I => \N__42088\
        );

    \I__7371\ : InMux
    port map (
            O => \N__42092\,
            I => \N__42083\
        );

    \I__7370\ : InMux
    port map (
            O => \N__42091\,
            I => \N__42083\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__42088\,
            I => data_in_3_4
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__42083\,
            I => data_in_3_4
        );

    \I__7367\ : InMux
    port map (
            O => \N__42078\,
            I => \N__42075\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__42075\,
            I => \N__42072\
        );

    \I__7365\ : Span4Mux_v
    port map (
            O => \N__42072\,
            I => \N__42069\
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__42069\,
            I => n2334
        );

    \I__7363\ : CascadeMux
    port map (
            O => \N__42066\,
            I => \N__42060\
        );

    \I__7362\ : InMux
    port map (
            O => \N__42065\,
            I => \N__42057\
        );

    \I__7361\ : InMux
    port map (
            O => \N__42064\,
            I => \N__42054\
        );

    \I__7360\ : InMux
    port map (
            O => \N__42063\,
            I => \N__42049\
        );

    \I__7359\ : InMux
    port map (
            O => \N__42060\,
            I => \N__42049\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__42057\,
            I => data_in_1_0
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__42054\,
            I => data_in_1_0
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__42049\,
            I => data_in_1_0
        );

    \I__7355\ : InMux
    port map (
            O => \N__42042\,
            I => \N__42039\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__42036\
        );

    \I__7353\ : Span4Mux_v
    port map (
            O => \N__42036\,
            I => \N__42033\
        );

    \I__7352\ : Span4Mux_v
    port map (
            O => \N__42033\,
            I => \N__42030\
        );

    \I__7351\ : Odrv4
    port map (
            O => \N__42030\,
            I => n2349
        );

    \I__7350\ : InMux
    port map (
            O => \N__42027\,
            I => \N__42023\
        );

    \I__7349\ : InMux
    port map (
            O => \N__42026\,
            I => \N__42019\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__42023\,
            I => \N__42014\
        );

    \I__7347\ : InMux
    port map (
            O => \N__42022\,
            I => \N__42011\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__42019\,
            I => \N__42008\
        );

    \I__7345\ : InMux
    port map (
            O => \N__42018\,
            I => \N__42004\
        );

    \I__7344\ : InMux
    port map (
            O => \N__42017\,
            I => \N__42001\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__42014\,
            I => \N__41996\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__42011\,
            I => \N__41996\
        );

    \I__7341\ : Span4Mux_v
    port map (
            O => \N__42008\,
            I => \N__41993\
        );

    \I__7340\ : InMux
    port map (
            O => \N__42007\,
            I => \N__41990\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__42004\,
            I => \N__41987\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__42001\,
            I => \N__41984\
        );

    \I__7337\ : Span4Mux_v
    port map (
            O => \N__41996\,
            I => \N__41981\
        );

    \I__7336\ : Sp12to4
    port map (
            O => \N__41993\,
            I => \N__41978\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__41990\,
            I => \N__41975\
        );

    \I__7334\ : Span4Mux_h
    port map (
            O => \N__41987\,
            I => \N__41972\
        );

    \I__7333\ : Span4Mux_v
    port map (
            O => \N__41984\,
            I => \N__41967\
        );

    \I__7332\ : Span4Mux_v
    port map (
            O => \N__41981\,
            I => \N__41967\
        );

    \I__7331\ : Span12Mux_h
    port map (
            O => \N__41978\,
            I => \N__41964\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__41975\,
            I => \N__41959\
        );

    \I__7329\ : Span4Mux_v
    port map (
            O => \N__41972\,
            I => \N__41959\
        );

    \I__7328\ : Odrv4
    port map (
            O => \N__41967\,
            I => \c0.rx.r_SM_Main_2_N_3680_2\
        );

    \I__7327\ : Odrv12
    port map (
            O => \N__41964\,
            I => \c0.rx.r_SM_Main_2_N_3680_2\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__41959\,
            I => \c0.rx.r_SM_Main_2_N_3680_2\
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__41952\,
            I => \N__41949\
        );

    \I__7324\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41946\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__41946\,
            I => \N__41940\
        );

    \I__7322\ : InMux
    port map (
            O => \N__41945\,
            I => \N__41935\
        );

    \I__7321\ : InMux
    port map (
            O => \N__41944\,
            I => \N__41935\
        );

    \I__7320\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41932\
        );

    \I__7319\ : Odrv4
    port map (
            O => \N__41940\,
            I => \c0.n24028\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__41935\,
            I => \c0.n24028\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__41932\,
            I => \c0.n24028\
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__41925\,
            I => \c0.n14_adj_4478_cascade_\
        );

    \I__7315\ : InMux
    port map (
            O => \N__41922\,
            I => \N__41916\
        );

    \I__7314\ : InMux
    port map (
            O => \N__41921\,
            I => \N__41916\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__41916\,
            I => \c0.n22193\
        );

    \I__7312\ : InMux
    port map (
            O => \N__41913\,
            I => \N__41908\
        );

    \I__7311\ : InMux
    port map (
            O => \N__41912\,
            I => \N__41904\
        );

    \I__7310\ : InMux
    port map (
            O => \N__41911\,
            I => \N__41901\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__41908\,
            I => \N__41898\
        );

    \I__7308\ : InMux
    port map (
            O => \N__41907\,
            I => \N__41895\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__41904\,
            I => \N__41890\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__41901\,
            I => \N__41890\
        );

    \I__7305\ : Span12Mux_v
    port map (
            O => \N__41898\,
            I => \N__41885\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__41895\,
            I => \N__41885\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__41890\,
            I => \N__41882\
        );

    \I__7302\ : Odrv12
    port map (
            O => \N__41885\,
            I => \c0.n13422\
        );

    \I__7301\ : Odrv4
    port map (
            O => \N__41882\,
            I => \c0.n13422\
        );

    \I__7300\ : CascadeMux
    port map (
            O => \N__41877\,
            I => \N__41874\
        );

    \I__7299\ : InMux
    port map (
            O => \N__41874\,
            I => \N__41871\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__41871\,
            I => \N__41868\
        );

    \I__7297\ : Odrv4
    port map (
            O => \N__41868\,
            I => \c0.n22722\
        );

    \I__7296\ : InMux
    port map (
            O => \N__41865\,
            I => \N__41862\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__41862\,
            I => \N__41858\
        );

    \I__7294\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41855\
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__41858\,
            I => \data_out_frame_29__2__N_1748\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__41855\,
            I => \data_out_frame_29__2__N_1748\
        );

    \I__7291\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41847\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41844\
        );

    \I__7289\ : Span12Mux_v
    port map (
            O => \N__41844\,
            I => \N__41841\
        );

    \I__7288\ : Odrv12
    port map (
            O => \N__41841\,
            I => \c0.n19_adj_4720\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__41838\,
            I => \N__41834\
        );

    \I__7286\ : InMux
    port map (
            O => \N__41837\,
            I => \N__41831\
        );

    \I__7285\ : InMux
    port map (
            O => \N__41834\,
            I => \N__41828\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__41831\,
            I => \N__41825\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__41828\,
            I => \N__41822\
        );

    \I__7282\ : Span4Mux_h
    port map (
            O => \N__41825\,
            I => \N__41815\
        );

    \I__7281\ : Span4Mux_v
    port map (
            O => \N__41822\,
            I => \N__41815\
        );

    \I__7280\ : InMux
    port map (
            O => \N__41821\,
            I => \N__41810\
        );

    \I__7279\ : InMux
    port map (
            O => \N__41820\,
            I => \N__41810\
        );

    \I__7278\ : Odrv4
    port map (
            O => \N__41815\,
            I => data_in_2_1
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__41810\,
            I => data_in_2_1
        );

    \I__7276\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41802\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__41802\,
            I => \N__41798\
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__41801\,
            I => \N__41795\
        );

    \I__7273\ : Span4Mux_h
    port map (
            O => \N__41798\,
            I => \N__41792\
        );

    \I__7272\ : InMux
    port map (
            O => \N__41795\,
            I => \N__41789\
        );

    \I__7271\ : Span4Mux_v
    port map (
            O => \N__41792\,
            I => \N__41786\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__41789\,
            I => data_out_frame_29_3
        );

    \I__7269\ : Odrv4
    port map (
            O => \N__41786\,
            I => data_out_frame_29_3
        );

    \I__7268\ : CascadeMux
    port map (
            O => \N__41781\,
            I => \N__41776\
        );

    \I__7267\ : CascadeMux
    port map (
            O => \N__41780\,
            I => \N__41773\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__41779\,
            I => \N__41770\
        );

    \I__7265\ : InMux
    port map (
            O => \N__41776\,
            I => \N__41767\
        );

    \I__7264\ : InMux
    port map (
            O => \N__41773\,
            I => \N__41764\
        );

    \I__7263\ : InMux
    port map (
            O => \N__41770\,
            I => \N__41761\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__41767\,
            I => \N__41757\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__41764\,
            I => \N__41754\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__41761\,
            I => \N__41749\
        );

    \I__7259\ : InMux
    port map (
            O => \N__41760\,
            I => \N__41746\
        );

    \I__7258\ : Span12Mux_v
    port map (
            O => \N__41757\,
            I => \N__41743\
        );

    \I__7257\ : Span12Mux_h
    port map (
            O => \N__41754\,
            I => \N__41740\
        );

    \I__7256\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41737\
        );

    \I__7255\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41734\
        );

    \I__7254\ : Span4Mux_v
    port map (
            O => \N__41749\,
            I => \N__41731\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__41746\,
            I => encoder1_position_12
        );

    \I__7252\ : Odrv12
    port map (
            O => \N__41743\,
            I => encoder1_position_12
        );

    \I__7251\ : Odrv12
    port map (
            O => \N__41740\,
            I => encoder1_position_12
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__41737\,
            I => encoder1_position_12
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__41734\,
            I => encoder1_position_12
        );

    \I__7248\ : Odrv4
    port map (
            O => \N__41731\,
            I => encoder1_position_12
        );

    \I__7247\ : InMux
    port map (
            O => \N__41718\,
            I => \N__41715\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__41715\,
            I => \N__41711\
        );

    \I__7245\ : InMux
    port map (
            O => \N__41714\,
            I => \N__41708\
        );

    \I__7244\ : Span4Mux_v
    port map (
            O => \N__41711\,
            I => \N__41705\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__41708\,
            I => data_out_frame_12_4
        );

    \I__7242\ : Odrv4
    port map (
            O => \N__41705\,
            I => data_out_frame_12_4
        );

    \I__7241\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41695\
        );

    \I__7240\ : InMux
    port map (
            O => \N__41699\,
            I => \N__41692\
        );

    \I__7239\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41689\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__41695\,
            I => data_in_0_3
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__41692\,
            I => data_in_0_3
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__41689\,
            I => data_in_0_3
        );

    \I__7235\ : InMux
    port map (
            O => \N__41682\,
            I => \N__41679\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__41679\,
            I => \N__41676\
        );

    \I__7233\ : Span4Mux_h
    port map (
            O => \N__41676\,
            I => \N__41673\
        );

    \I__7232\ : Odrv4
    port map (
            O => \N__41673\,
            I => \c0.n15\
        );

    \I__7231\ : CascadeMux
    port map (
            O => \N__41670\,
            I => \c0.n21311_cascade_\
        );

    \I__7230\ : InMux
    port map (
            O => \N__41667\,
            I => \N__41664\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__41664\,
            I => \N__41661\
        );

    \I__7228\ : Span4Mux_v
    port map (
            O => \N__41661\,
            I => \N__41658\
        );

    \I__7227\ : Span4Mux_h
    port map (
            O => \N__41658\,
            I => \N__41654\
        );

    \I__7226\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41651\
        );

    \I__7225\ : Odrv4
    port map (
            O => \N__41654\,
            I => \c0.n21244\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__41651\,
            I => \c0.n21244\
        );

    \I__7223\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41643\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__41643\,
            I => \N__41640\
        );

    \I__7221\ : Span4Mux_h
    port map (
            O => \N__41640\,
            I => \N__41636\
        );

    \I__7220\ : InMux
    port map (
            O => \N__41639\,
            I => \N__41633\
        );

    \I__7219\ : Span4Mux_h
    port map (
            O => \N__41636\,
            I => \N__41630\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__41633\,
            I => \c0.n21496\
        );

    \I__7217\ : Odrv4
    port map (
            O => \N__41630\,
            I => \c0.n21496\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__41625\,
            I => \c0.n21273_cascade_\
        );

    \I__7215\ : InMux
    port map (
            O => \N__41622\,
            I => \N__41619\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__41619\,
            I => \N__41616\
        );

    \I__7213\ : Span4Mux_h
    port map (
            O => \N__41616\,
            I => \N__41613\
        );

    \I__7212\ : Odrv4
    port map (
            O => \N__41613\,
            I => \c0.data_out_frame_29_6\
        );

    \I__7211\ : InMux
    port map (
            O => \N__41610\,
            I => \N__41607\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__41607\,
            I => \N__41604\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__41604\,
            I => \c0.data_out_frame_28_6\
        );

    \I__7208\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41598\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__41598\,
            I => \N__41595\
        );

    \I__7206\ : Span12Mux_h
    port map (
            O => \N__41595\,
            I => \N__41592\
        );

    \I__7205\ : Odrv12
    port map (
            O => \N__41592\,
            I => \c0.n26_adj_4702\
        );

    \I__7204\ : InMux
    port map (
            O => \N__41589\,
            I => \N__41585\
        );

    \I__7203\ : InMux
    port map (
            O => \N__41588\,
            I => \N__41582\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__41585\,
            I => \N__41577\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__41582\,
            I => \N__41577\
        );

    \I__7200\ : Span4Mux_h
    port map (
            O => \N__41577\,
            I => \N__41574\
        );

    \I__7199\ : Odrv4
    port map (
            O => \N__41574\,
            I => \c0.n22617\
        );

    \I__7198\ : InMux
    port map (
            O => \N__41571\,
            I => \N__41568\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__41568\,
            I => \N__41565\
        );

    \I__7196\ : Span4Mux_v
    port map (
            O => \N__41565\,
            I => \N__41559\
        );

    \I__7195\ : InMux
    port map (
            O => \N__41564\,
            I => \N__41556\
        );

    \I__7194\ : InMux
    port map (
            O => \N__41563\,
            I => \N__41551\
        );

    \I__7193\ : InMux
    port map (
            O => \N__41562\,
            I => \N__41551\
        );

    \I__7192\ : Span4Mux_h
    port map (
            O => \N__41559\,
            I => \N__41546\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__41556\,
            I => \N__41546\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__41551\,
            I => \c0.n20341\
        );

    \I__7189\ : Odrv4
    port map (
            O => \N__41546\,
            I => \c0.n20341\
        );

    \I__7188\ : CascadeMux
    port map (
            O => \N__41541\,
            I => \c0.n18_adj_4684_cascade_\
        );

    \I__7187\ : InMux
    port map (
            O => \N__41538\,
            I => \N__41532\
        );

    \I__7186\ : InMux
    port map (
            O => \N__41537\,
            I => \N__41529\
        );

    \I__7185\ : InMux
    port map (
            O => \N__41536\,
            I => \N__41524\
        );

    \I__7184\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41524\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__41532\,
            I => \c0.n13268\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__41529\,
            I => \c0.n13268\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__41524\,
            I => \c0.n13268\
        );

    \I__7180\ : InMux
    port map (
            O => \N__41517\,
            I => \N__41514\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__41514\,
            I => \N__41511\
        );

    \I__7178\ : Span4Mux_v
    port map (
            O => \N__41511\,
            I => \N__41508\
        );

    \I__7177\ : Odrv4
    port map (
            O => \N__41508\,
            I => \c0.n15_adj_4686\
        );

    \I__7176\ : CascadeMux
    port map (
            O => \N__41505\,
            I => \c0.n20_adj_4685_cascade_\
        );

    \I__7175\ : InMux
    port map (
            O => \N__41502\,
            I => \N__41499\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__41499\,
            I => \N__41496\
        );

    \I__7173\ : Span4Mux_h
    port map (
            O => \N__41496\,
            I => \N__41492\
        );

    \I__7172\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41488\
        );

    \I__7171\ : Span4Mux_h
    port map (
            O => \N__41492\,
            I => \N__41485\
        );

    \I__7170\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41482\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__41488\,
            I => \N__41479\
        );

    \I__7168\ : Odrv4
    port map (
            O => \N__41485\,
            I => \c0.n21475\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__41482\,
            I => \c0.n21475\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__41479\,
            I => \c0.n21475\
        );

    \I__7165\ : InMux
    port map (
            O => \N__41472\,
            I => \N__41469\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__41469\,
            I => \N__41466\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__41466\,
            I => \N__41463\
        );

    \I__7162\ : Span4Mux_h
    port map (
            O => \N__41463\,
            I => \N__41460\
        );

    \I__7161\ : Sp12to4
    port map (
            O => \N__41460\,
            I => \N__41457\
        );

    \I__7160\ : Odrv12
    port map (
            O => \N__41457\,
            I => \c0.data_out_frame_28_7\
        );

    \I__7159\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41451\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__41451\,
            I => \c0.n22461\
        );

    \I__7157\ : InMux
    port map (
            O => \N__41448\,
            I => \N__41444\
        );

    \I__7156\ : InMux
    port map (
            O => \N__41447\,
            I => \N__41441\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__41444\,
            I => \c0.n21358\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__41441\,
            I => \c0.n21358\
        );

    \I__7153\ : CascadeMux
    port map (
            O => \N__41436\,
            I => \c0.n22461_cascade_\
        );

    \I__7152\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41426\
        );

    \I__7151\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41423\
        );

    \I__7150\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41420\
        );

    \I__7149\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41417\
        );

    \I__7148\ : InMux
    port map (
            O => \N__41429\,
            I => \N__41414\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__41426\,
            I => \N__41409\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__41423\,
            I => \N__41400\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__41420\,
            I => \N__41400\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__41417\,
            I => \N__41400\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__41414\,
            I => \N__41400\
        );

    \I__7142\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41397\
        );

    \I__7141\ : InMux
    port map (
            O => \N__41412\,
            I => \N__41394\
        );

    \I__7140\ : Span4Mux_v
    port map (
            O => \N__41409\,
            I => \N__41391\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__41400\,
            I => \N__41386\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__41397\,
            I => \N__41386\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__41394\,
            I => \N__41383\
        );

    \I__7136\ : Span4Mux_v
    port map (
            O => \N__41391\,
            I => \N__41378\
        );

    \I__7135\ : Span4Mux_v
    port map (
            O => \N__41386\,
            I => \N__41378\
        );

    \I__7134\ : Span4Mux_h
    port map (
            O => \N__41383\,
            I => \N__41375\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__41378\,
            I => \c0.n21406\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__41375\,
            I => \c0.n21406\
        );

    \I__7131\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41367\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__41367\,
            I => \N__41361\
        );

    \I__7129\ : InMux
    port map (
            O => \N__41366\,
            I => \N__41358\
        );

    \I__7128\ : InMux
    port map (
            O => \N__41365\,
            I => \N__41355\
        );

    \I__7127\ : InMux
    port map (
            O => \N__41364\,
            I => \N__41352\
        );

    \I__7126\ : Span4Mux_v
    port map (
            O => \N__41361\,
            I => \N__41347\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__41358\,
            I => \N__41347\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__41355\,
            I => \N__41342\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__41352\,
            I => \N__41342\
        );

    \I__7122\ : Span4Mux_h
    port map (
            O => \N__41347\,
            I => \N__41339\
        );

    \I__7121\ : Odrv12
    port map (
            O => \N__41342\,
            I => \c0.n21441\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__41339\,
            I => \c0.n21441\
        );

    \I__7119\ : CascadeMux
    port map (
            O => \N__41334\,
            I => \N__41331\
        );

    \I__7118\ : InMux
    port map (
            O => \N__41331\,
            I => \N__41328\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__41328\,
            I => \N__41322\
        );

    \I__7116\ : CascadeMux
    port map (
            O => \N__41327\,
            I => \N__41319\
        );

    \I__7115\ : InMux
    port map (
            O => \N__41326\,
            I => \N__41314\
        );

    \I__7114\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41311\
        );

    \I__7113\ : Span4Mux_h
    port map (
            O => \N__41322\,
            I => \N__41308\
        );

    \I__7112\ : InMux
    port map (
            O => \N__41319\,
            I => \N__41305\
        );

    \I__7111\ : InMux
    port map (
            O => \N__41318\,
            I => \N__41302\
        );

    \I__7110\ : InMux
    port map (
            O => \N__41317\,
            I => \N__41299\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__41314\,
            I => \N__41296\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__41311\,
            I => encoder0_position_25
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__41308\,
            I => encoder0_position_25
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__41305\,
            I => encoder0_position_25
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__41302\,
            I => encoder0_position_25
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__41299\,
            I => encoder0_position_25
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__41296\,
            I => encoder0_position_25
        );

    \I__7102\ : InMux
    port map (
            O => \N__41283\,
            I => \N__41280\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__41280\,
            I => \N__41277\
        );

    \I__7100\ : Span4Mux_v
    port map (
            O => \N__41277\,
            I => \N__41273\
        );

    \I__7099\ : InMux
    port map (
            O => \N__41276\,
            I => \N__41270\
        );

    \I__7098\ : Span4Mux_h
    port map (
            O => \N__41273\,
            I => \N__41267\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__41270\,
            I => data_out_frame_6_1
        );

    \I__7096\ : Odrv4
    port map (
            O => \N__41267\,
            I => data_out_frame_6_1
        );

    \I__7095\ : InMux
    port map (
            O => \N__41262\,
            I => \N__41258\
        );

    \I__7094\ : CascadeMux
    port map (
            O => \N__41261\,
            I => \N__41255\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__41258\,
            I => \N__41252\
        );

    \I__7092\ : InMux
    port map (
            O => \N__41255\,
            I => \N__41249\
        );

    \I__7091\ : Span4Mux_h
    port map (
            O => \N__41252\,
            I => \N__41246\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__41249\,
            I => data_out_frame_29_2
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__41246\,
            I => data_out_frame_29_2
        );

    \I__7088\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41238\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__41238\,
            I => \c0.n12_adj_4312\
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__41235\,
            I => \c0.n24113_cascade_\
        );

    \I__7085\ : InMux
    port map (
            O => \N__41232\,
            I => \N__41226\
        );

    \I__7084\ : InMux
    port map (
            O => \N__41231\,
            I => \N__41223\
        );

    \I__7083\ : InMux
    port map (
            O => \N__41230\,
            I => \N__41220\
        );

    \I__7082\ : InMux
    port map (
            O => \N__41229\,
            I => \N__41217\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__41226\,
            I => \N__41214\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__41223\,
            I => \N__41211\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__41220\,
            I => \N__41208\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__41217\,
            I => \N__41205\
        );

    \I__7077\ : Span4Mux_h
    port map (
            O => \N__41214\,
            I => \N__41202\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__41211\,
            I => \N__41197\
        );

    \I__7075\ : Span4Mux_v
    port map (
            O => \N__41208\,
            I => \N__41197\
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__41205\,
            I => \c0.n10529\
        );

    \I__7073\ : Odrv4
    port map (
            O => \N__41202\,
            I => \c0.n10529\
        );

    \I__7072\ : Odrv4
    port map (
            O => \N__41197\,
            I => \c0.n10529\
        );

    \I__7071\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41186\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__41189\,
            I => \N__41182\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__41186\,
            I => \N__41176\
        );

    \I__7068\ : InMux
    port map (
            O => \N__41185\,
            I => \N__41173\
        );

    \I__7067\ : InMux
    port map (
            O => \N__41182\,
            I => \N__41169\
        );

    \I__7066\ : InMux
    port map (
            O => \N__41181\,
            I => \N__41164\
        );

    \I__7065\ : InMux
    port map (
            O => \N__41180\,
            I => \N__41164\
        );

    \I__7064\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41161\
        );

    \I__7063\ : Span4Mux_v
    port map (
            O => \N__41176\,
            I => \N__41156\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__41173\,
            I => \N__41156\
        );

    \I__7061\ : CascadeMux
    port map (
            O => \N__41172\,
            I => \N__41153\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__41169\,
            I => \N__41148\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__41164\,
            I => \N__41148\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__41161\,
            I => \N__41143\
        );

    \I__7057\ : Span4Mux_v
    port map (
            O => \N__41156\,
            I => \N__41143\
        );

    \I__7056\ : InMux
    port map (
            O => \N__41153\,
            I => \N__41140\
        );

    \I__7055\ : Span4Mux_v
    port map (
            O => \N__41148\,
            I => \N__41136\
        );

    \I__7054\ : Span4Mux_h
    port map (
            O => \N__41143\,
            I => \N__41131\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__41140\,
            I => \N__41131\
        );

    \I__7052\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41128\
        );

    \I__7051\ : Span4Mux_h
    port map (
            O => \N__41136\,
            I => \N__41125\
        );

    \I__7050\ : Span4Mux_h
    port map (
            O => \N__41131\,
            I => \N__41122\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__41128\,
            I => encoder1_position_5
        );

    \I__7048\ : Odrv4
    port map (
            O => \N__41125\,
            I => encoder1_position_5
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__41122\,
            I => encoder1_position_5
        );

    \I__7046\ : CascadeMux
    port map (
            O => \N__41115\,
            I => \N__41112\
        );

    \I__7045\ : InMux
    port map (
            O => \N__41112\,
            I => \N__41109\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__41109\,
            I => \N__41099\
        );

    \I__7043\ : InMux
    port map (
            O => \N__41108\,
            I => \N__41094\
        );

    \I__7042\ : InMux
    port map (
            O => \N__41107\,
            I => \N__41094\
        );

    \I__7041\ : InMux
    port map (
            O => \N__41106\,
            I => \N__41089\
        );

    \I__7040\ : InMux
    port map (
            O => \N__41105\,
            I => \N__41089\
        );

    \I__7039\ : InMux
    port map (
            O => \N__41104\,
            I => \N__41086\
        );

    \I__7038\ : InMux
    port map (
            O => \N__41103\,
            I => \N__41081\
        );

    \I__7037\ : InMux
    port map (
            O => \N__41102\,
            I => \N__41081\
        );

    \I__7036\ : Span4Mux_h
    port map (
            O => \N__41099\,
            I => \N__41074\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__41094\,
            I => \N__41074\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__41089\,
            I => \N__41074\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__41086\,
            I => \c0.n21364\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__41081\,
            I => \c0.n21364\
        );

    \I__7031\ : Odrv4
    port map (
            O => \N__41074\,
            I => \c0.n21364\
        );

    \I__7030\ : InMux
    port map (
            O => \N__41067\,
            I => \N__41063\
        );

    \I__7029\ : InMux
    port map (
            O => \N__41066\,
            I => \N__41060\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__41063\,
            I => \c0.n24113\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__41060\,
            I => \c0.n24113\
        );

    \I__7026\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41050\
        );

    \I__7025\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41047\
        );

    \I__7024\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41042\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__41050\,
            I => \N__41039\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__41047\,
            I => \N__41035\
        );

    \I__7021\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41030\
        );

    \I__7020\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41027\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__41042\,
            I => \N__41014\
        );

    \I__7018\ : Span4Mux_v
    port map (
            O => \N__41039\,
            I => \N__41011\
        );

    \I__7017\ : InMux
    port map (
            O => \N__41038\,
            I => \N__41005\
        );

    \I__7016\ : Span4Mux_v
    port map (
            O => \N__41035\,
            I => \N__41002\
        );

    \I__7015\ : InMux
    port map (
            O => \N__41034\,
            I => \N__40997\
        );

    \I__7014\ : CascadeMux
    port map (
            O => \N__41033\,
            I => \N__40991\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__41030\,
            I => \N__40986\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__41027\,
            I => \N__40986\
        );

    \I__7011\ : InMux
    port map (
            O => \N__41026\,
            I => \N__40983\
        );

    \I__7010\ : InMux
    port map (
            O => \N__41025\,
            I => \N__40980\
        );

    \I__7009\ : InMux
    port map (
            O => \N__41024\,
            I => \N__40973\
        );

    \I__7008\ : InMux
    port map (
            O => \N__41023\,
            I => \N__40973\
        );

    \I__7007\ : InMux
    port map (
            O => \N__41022\,
            I => \N__40973\
        );

    \I__7006\ : InMux
    port map (
            O => \N__41021\,
            I => \N__40966\
        );

    \I__7005\ : InMux
    port map (
            O => \N__41020\,
            I => \N__40966\
        );

    \I__7004\ : InMux
    port map (
            O => \N__41019\,
            I => \N__40966\
        );

    \I__7003\ : InMux
    port map (
            O => \N__41018\,
            I => \N__40961\
        );

    \I__7002\ : InMux
    port map (
            O => \N__41017\,
            I => \N__40961\
        );

    \I__7001\ : Span4Mux_v
    port map (
            O => \N__41014\,
            I => \N__40958\
        );

    \I__7000\ : Span4Mux_v
    port map (
            O => \N__41011\,
            I => \N__40955\
        );

    \I__6999\ : InMux
    port map (
            O => \N__41010\,
            I => \N__40950\
        );

    \I__6998\ : InMux
    port map (
            O => \N__41009\,
            I => \N__40950\
        );

    \I__6997\ : InMux
    port map (
            O => \N__41008\,
            I => \N__40946\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__41005\,
            I => \N__40941\
        );

    \I__6995\ : Span4Mux_v
    port map (
            O => \N__41002\,
            I => \N__40941\
        );

    \I__6994\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40936\
        );

    \I__6993\ : InMux
    port map (
            O => \N__41000\,
            I => \N__40936\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__40997\,
            I => \N__40933\
        );

    \I__6991\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40930\
        );

    \I__6990\ : InMux
    port map (
            O => \N__40995\,
            I => \N__40926\
        );

    \I__6989\ : InMux
    port map (
            O => \N__40994\,
            I => \N__40923\
        );

    \I__6988\ : InMux
    port map (
            O => \N__40991\,
            I => \N__40920\
        );

    \I__6987\ : Span4Mux_v
    port map (
            O => \N__40986\,
            I => \N__40913\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__40983\,
            I => \N__40913\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__40980\,
            I => \N__40913\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__40973\,
            I => \N__40904\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__40966\,
            I => \N__40904\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__40961\,
            I => \N__40904\
        );

    \I__6981\ : Span4Mux_v
    port map (
            O => \N__40958\,
            I => \N__40904\
        );

    \I__6980\ : Span4Mux_v
    port map (
            O => \N__40955\,
            I => \N__40901\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__40950\,
            I => \N__40898\
        );

    \I__6978\ : InMux
    port map (
            O => \N__40949\,
            I => \N__40895\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__40946\,
            I => \N__40890\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__40941\,
            I => \N__40890\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__40936\,
            I => \N__40883\
        );

    \I__6974\ : Span4Mux_h
    port map (
            O => \N__40933\,
            I => \N__40883\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__40930\,
            I => \N__40883\
        );

    \I__6972\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40880\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__40926\,
            I => \N__40867\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__40923\,
            I => \N__40867\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__40920\,
            I => \N__40867\
        );

    \I__6968\ : Span4Mux_v
    port map (
            O => \N__40913\,
            I => \N__40867\
        );

    \I__6967\ : Span4Mux_v
    port map (
            O => \N__40904\,
            I => \N__40867\
        );

    \I__6966\ : Span4Mux_h
    port map (
            O => \N__40901\,
            I => \N__40867\
        );

    \I__6965\ : Odrv12
    port map (
            O => \N__40898\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__40895\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__40890\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6962\ : Odrv4
    port map (
            O => \N__40883\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__40880\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6960\ : Odrv4
    port map (
            O => \N__40867\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__6959\ : InMux
    port map (
            O => \N__40854\,
            I => \N__40851\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__40851\,
            I => \N__40848\
        );

    \I__6957\ : Span4Mux_h
    port map (
            O => \N__40848\,
            I => \N__40845\
        );

    \I__6956\ : Span4Mux_v
    port map (
            O => \N__40845\,
            I => \N__40842\
        );

    \I__6955\ : Span4Mux_v
    port map (
            O => \N__40842\,
            I => \N__40839\
        );

    \I__6954\ : Odrv4
    port map (
            O => \N__40839\,
            I => \c0.n5_adj_4217\
        );

    \I__6953\ : CascadeMux
    port map (
            O => \N__40836\,
            I => \N__40832\
        );

    \I__6952\ : InMux
    port map (
            O => \N__40835\,
            I => \N__40829\
        );

    \I__6951\ : InMux
    port map (
            O => \N__40832\,
            I => \N__40826\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__40829\,
            I => \N__40823\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__40826\,
            I => \N__40812\
        );

    \I__6948\ : Span4Mux_v
    port map (
            O => \N__40823\,
            I => \N__40801\
        );

    \I__6947\ : InMux
    port map (
            O => \N__40822\,
            I => \N__40796\
        );

    \I__6946\ : InMux
    port map (
            O => \N__40821\,
            I => \N__40796\
        );

    \I__6945\ : InMux
    port map (
            O => \N__40820\,
            I => \N__40793\
        );

    \I__6944\ : InMux
    port map (
            O => \N__40819\,
            I => \N__40790\
        );

    \I__6943\ : InMux
    port map (
            O => \N__40818\,
            I => \N__40787\
        );

    \I__6942\ : InMux
    port map (
            O => \N__40817\,
            I => \N__40782\
        );

    \I__6941\ : InMux
    port map (
            O => \N__40816\,
            I => \N__40782\
        );

    \I__6940\ : CascadeMux
    port map (
            O => \N__40815\,
            I => \N__40764\
        );

    \I__6939\ : Span4Mux_v
    port map (
            O => \N__40812\,
            I => \N__40761\
        );

    \I__6938\ : InMux
    port map (
            O => \N__40811\,
            I => \N__40758\
        );

    \I__6937\ : InMux
    port map (
            O => \N__40810\,
            I => \N__40755\
        );

    \I__6936\ : InMux
    port map (
            O => \N__40809\,
            I => \N__40746\
        );

    \I__6935\ : InMux
    port map (
            O => \N__40808\,
            I => \N__40746\
        );

    \I__6934\ : InMux
    port map (
            O => \N__40807\,
            I => \N__40746\
        );

    \I__6933\ : InMux
    port map (
            O => \N__40806\,
            I => \N__40746\
        );

    \I__6932\ : InMux
    port map (
            O => \N__40805\,
            I => \N__40741\
        );

    \I__6931\ : InMux
    port map (
            O => \N__40804\,
            I => \N__40741\
        );

    \I__6930\ : Span4Mux_v
    port map (
            O => \N__40801\,
            I => \N__40736\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__40796\,
            I => \N__40736\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__40793\,
            I => \N__40727\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__40790\,
            I => \N__40727\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__40787\,
            I => \N__40727\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__40782\,
            I => \N__40727\
        );

    \I__6924\ : InMux
    port map (
            O => \N__40781\,
            I => \N__40720\
        );

    \I__6923\ : InMux
    port map (
            O => \N__40780\,
            I => \N__40720\
        );

    \I__6922\ : InMux
    port map (
            O => \N__40779\,
            I => \N__40720\
        );

    \I__6921\ : InMux
    port map (
            O => \N__40778\,
            I => \N__40715\
        );

    \I__6920\ : InMux
    port map (
            O => \N__40777\,
            I => \N__40715\
        );

    \I__6919\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40706\
        );

    \I__6918\ : InMux
    port map (
            O => \N__40775\,
            I => \N__40706\
        );

    \I__6917\ : InMux
    port map (
            O => \N__40774\,
            I => \N__40706\
        );

    \I__6916\ : InMux
    port map (
            O => \N__40773\,
            I => \N__40706\
        );

    \I__6915\ : InMux
    port map (
            O => \N__40772\,
            I => \N__40703\
        );

    \I__6914\ : InMux
    port map (
            O => \N__40771\,
            I => \N__40694\
        );

    \I__6913\ : InMux
    port map (
            O => \N__40770\,
            I => \N__40694\
        );

    \I__6912\ : InMux
    port map (
            O => \N__40769\,
            I => \N__40694\
        );

    \I__6911\ : InMux
    port map (
            O => \N__40768\,
            I => \N__40694\
        );

    \I__6910\ : InMux
    port map (
            O => \N__40767\,
            I => \N__40689\
        );

    \I__6909\ : InMux
    port map (
            O => \N__40764\,
            I => \N__40689\
        );

    \I__6908\ : Span4Mux_h
    port map (
            O => \N__40761\,
            I => \N__40686\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__40758\,
            I => \N__40681\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__40755\,
            I => \N__40672\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__40746\,
            I => \N__40672\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__40741\,
            I => \N__40672\
        );

    \I__6903\ : Span4Mux_h
    port map (
            O => \N__40736\,
            I => \N__40672\
        );

    \I__6902\ : Span4Mux_v
    port map (
            O => \N__40727\,
            I => \N__40667\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__40720\,
            I => \N__40667\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__40715\,
            I => \N__40654\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__40706\,
            I => \N__40654\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__40703\,
            I => \N__40654\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__40694\,
            I => \N__40654\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__40689\,
            I => \N__40654\
        );

    \I__6895\ : Span4Mux_v
    port map (
            O => \N__40686\,
            I => \N__40654\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__40685\,
            I => \N__40651\
        );

    \I__6893\ : InMux
    port map (
            O => \N__40684\,
            I => \N__40645\
        );

    \I__6892\ : Span4Mux_v
    port map (
            O => \N__40681\,
            I => \N__40642\
        );

    \I__6891\ : Span4Mux_h
    port map (
            O => \N__40672\,
            I => \N__40639\
        );

    \I__6890\ : Span4Mux_v
    port map (
            O => \N__40667\,
            I => \N__40634\
        );

    \I__6889\ : Span4Mux_v
    port map (
            O => \N__40654\,
            I => \N__40634\
        );

    \I__6888\ : InMux
    port map (
            O => \N__40651\,
            I => \N__40627\
        );

    \I__6887\ : InMux
    port map (
            O => \N__40650\,
            I => \N__40627\
        );

    \I__6886\ : InMux
    port map (
            O => \N__40649\,
            I => \N__40627\
        );

    \I__6885\ : InMux
    port map (
            O => \N__40648\,
            I => \N__40624\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__40645\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6883\ : Odrv4
    port map (
            O => \N__40642\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__40639\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__40634\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__40627\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__40624\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6878\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40608\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__40608\,
            I => \N__40605\
        );

    \I__6876\ : Span4Mux_h
    port map (
            O => \N__40605\,
            I => \N__40602\
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__40602\,
            I => \c0.n24901\
        );

    \I__6874\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40596\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__40596\,
            I => \N__40593\
        );

    \I__6872\ : Odrv12
    port map (
            O => \N__40593\,
            I => \c0.n25062\
        );

    \I__6871\ : InMux
    port map (
            O => \N__40590\,
            I => \N__40587\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__40587\,
            I => \N__40584\
        );

    \I__6869\ : Span4Mux_h
    port map (
            O => \N__40584\,
            I => \N__40581\
        );

    \I__6868\ : Span4Mux_v
    port map (
            O => \N__40581\,
            I => \N__40578\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__40578\,
            I => n2260
        );

    \I__6866\ : CascadeMux
    port map (
            O => \N__40575\,
            I => \N__40570\
        );

    \I__6865\ : InMux
    port map (
            O => \N__40574\,
            I => \N__40559\
        );

    \I__6864\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40555\
        );

    \I__6863\ : InMux
    port map (
            O => \N__40570\,
            I => \N__40552\
        );

    \I__6862\ : InMux
    port map (
            O => \N__40569\,
            I => \N__40549\
        );

    \I__6861\ : InMux
    port map (
            O => \N__40568\,
            I => \N__40546\
        );

    \I__6860\ : InMux
    port map (
            O => \N__40567\,
            I => \N__40537\
        );

    \I__6859\ : CascadeMux
    port map (
            O => \N__40566\,
            I => \N__40532\
        );

    \I__6858\ : InMux
    port map (
            O => \N__40565\,
            I => \N__40529\
        );

    \I__6857\ : InMux
    port map (
            O => \N__40564\,
            I => \N__40519\
        );

    \I__6856\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40519\
        );

    \I__6855\ : InMux
    port map (
            O => \N__40562\,
            I => \N__40519\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__40559\,
            I => \N__40516\
        );

    \I__6853\ : InMux
    port map (
            O => \N__40558\,
            I => \N__40513\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__40555\,
            I => \N__40504\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__40552\,
            I => \N__40504\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__40549\,
            I => \N__40504\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__40546\,
            I => \N__40504\
        );

    \I__6848\ : InMux
    port map (
            O => \N__40545\,
            I => \N__40499\
        );

    \I__6847\ : InMux
    port map (
            O => \N__40544\,
            I => \N__40499\
        );

    \I__6846\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40494\
        );

    \I__6845\ : InMux
    port map (
            O => \N__40542\,
            I => \N__40494\
        );

    \I__6844\ : InMux
    port map (
            O => \N__40541\,
            I => \N__40489\
        );

    \I__6843\ : InMux
    port map (
            O => \N__40540\,
            I => \N__40489\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__40537\,
            I => \N__40486\
        );

    \I__6841\ : InMux
    port map (
            O => \N__40536\,
            I => \N__40480\
        );

    \I__6840\ : InMux
    port map (
            O => \N__40535\,
            I => \N__40480\
        );

    \I__6839\ : InMux
    port map (
            O => \N__40532\,
            I => \N__40476\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__40529\,
            I => \N__40473\
        );

    \I__6837\ : InMux
    port map (
            O => \N__40528\,
            I => \N__40468\
        );

    \I__6836\ : InMux
    port map (
            O => \N__40527\,
            I => \N__40468\
        );

    \I__6835\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40464\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__40519\,
            I => \N__40457\
        );

    \I__6833\ : Span4Mux_v
    port map (
            O => \N__40516\,
            I => \N__40457\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__40513\,
            I => \N__40457\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__40504\,
            I => \N__40452\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__40499\,
            I => \N__40452\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__40494\,
            I => \N__40447\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__40489\,
            I => \N__40447\
        );

    \I__6827\ : Span4Mux_h
    port map (
            O => \N__40486\,
            I => \N__40444\
        );

    \I__6826\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40441\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__40480\,
            I => \N__40437\
        );

    \I__6824\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40434\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__40476\,
            I => \N__40431\
        );

    \I__6822\ : Span4Mux_v
    port map (
            O => \N__40473\,
            I => \N__40426\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__40468\,
            I => \N__40426\
        );

    \I__6820\ : InMux
    port map (
            O => \N__40467\,
            I => \N__40423\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__40464\,
            I => \N__40420\
        );

    \I__6818\ : Span4Mux_v
    port map (
            O => \N__40457\,
            I => \N__40417\
        );

    \I__6817\ : Span4Mux_h
    port map (
            O => \N__40452\,
            I => \N__40414\
        );

    \I__6816\ : Span4Mux_h
    port map (
            O => \N__40447\,
            I => \N__40402\
        );

    \I__6815\ : Span4Mux_h
    port map (
            O => \N__40444\,
            I => \N__40402\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__40441\,
            I => \N__40402\
        );

    \I__6813\ : InMux
    port map (
            O => \N__40440\,
            I => \N__40399\
        );

    \I__6812\ : Span4Mux_v
    port map (
            O => \N__40437\,
            I => \N__40396\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__40434\,
            I => \N__40391\
        );

    \I__6810\ : Span4Mux_v
    port map (
            O => \N__40431\,
            I => \N__40391\
        );

    \I__6809\ : Span4Mux_h
    port map (
            O => \N__40426\,
            I => \N__40380\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__40423\,
            I => \N__40380\
        );

    \I__6807\ : Span4Mux_h
    port map (
            O => \N__40420\,
            I => \N__40380\
        );

    \I__6806\ : Span4Mux_h
    port map (
            O => \N__40417\,
            I => \N__40380\
        );

    \I__6805\ : Span4Mux_v
    port map (
            O => \N__40414\,
            I => \N__40380\
        );

    \I__6804\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40377\
        );

    \I__6803\ : InMux
    port map (
            O => \N__40412\,
            I => \N__40374\
        );

    \I__6802\ : InMux
    port map (
            O => \N__40411\,
            I => \N__40371\
        );

    \I__6801\ : InMux
    port map (
            O => \N__40410\,
            I => \N__40368\
        );

    \I__6800\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40365\
        );

    \I__6799\ : Span4Mux_v
    port map (
            O => \N__40402\,
            I => \N__40362\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__40399\,
            I => \N__40355\
        );

    \I__6797\ : Span4Mux_v
    port map (
            O => \N__40396\,
            I => \N__40355\
        );

    \I__6796\ : Span4Mux_h
    port map (
            O => \N__40391\,
            I => \N__40355\
        );

    \I__6795\ : Span4Mux_v
    port map (
            O => \N__40380\,
            I => \N__40352\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__40377\,
            I => count_enable_adj_4769
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__40374\,
            I => count_enable_adj_4769
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__40371\,
            I => count_enable_adj_4769
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__40368\,
            I => count_enable_adj_4769
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__40365\,
            I => count_enable_adj_4769
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__40362\,
            I => count_enable_adj_4769
        );

    \I__6788\ : Odrv4
    port map (
            O => \N__40355\,
            I => count_enable_adj_4769
        );

    \I__6787\ : Odrv4
    port map (
            O => \N__40352\,
            I => count_enable_adj_4769
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__40335\,
            I => \N__40332\
        );

    \I__6785\ : InMux
    port map (
            O => \N__40332\,
            I => \N__40328\
        );

    \I__6784\ : InMux
    port map (
            O => \N__40331\,
            I => \N__40325\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__40328\,
            I => \N__40321\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__40325\,
            I => \N__40318\
        );

    \I__6781\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40315\
        );

    \I__6780\ : Sp12to4
    port map (
            O => \N__40321\,
            I => \N__40311\
        );

    \I__6779\ : Span4Mux_v
    port map (
            O => \N__40318\,
            I => \N__40308\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__40315\,
            I => \N__40305\
        );

    \I__6777\ : InMux
    port map (
            O => \N__40314\,
            I => \N__40302\
        );

    \I__6776\ : Span12Mux_h
    port map (
            O => \N__40311\,
            I => \N__40299\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__40308\,
            I => \N__40296\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__40305\,
            I => \N__40293\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__40302\,
            I => encoder1_position_31
        );

    \I__6772\ : Odrv12
    port map (
            O => \N__40299\,
            I => encoder1_position_31
        );

    \I__6771\ : Odrv4
    port map (
            O => \N__40296\,
            I => encoder1_position_31
        );

    \I__6770\ : Odrv4
    port map (
            O => \N__40293\,
            I => encoder1_position_31
        );

    \I__6769\ : InMux
    port map (
            O => \N__40284\,
            I => \N__40281\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__40281\,
            I => n2338
        );

    \I__6767\ : CascadeMux
    port map (
            O => \N__40278\,
            I => \N__40275\
        );

    \I__6766\ : InMux
    port map (
            O => \N__40275\,
            I => \N__40271\
        );

    \I__6765\ : InMux
    port map (
            O => \N__40274\,
            I => \N__40268\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__40271\,
            I => \N__40261\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__40268\,
            I => \N__40258\
        );

    \I__6762\ : InMux
    port map (
            O => \N__40267\,
            I => \N__40255\
        );

    \I__6761\ : InMux
    port map (
            O => \N__40266\,
            I => \N__40252\
        );

    \I__6760\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40249\
        );

    \I__6759\ : InMux
    port map (
            O => \N__40264\,
            I => \N__40246\
        );

    \I__6758\ : Span4Mux_h
    port map (
            O => \N__40261\,
            I => \N__40241\
        );

    \I__6757\ : Span4Mux_h
    port map (
            O => \N__40258\,
            I => \N__40241\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__40255\,
            I => \N__40236\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__40252\,
            I => \N__40236\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__40249\,
            I => encoder1_position_21
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__40246\,
            I => encoder1_position_21
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__40241\,
            I => encoder1_position_21
        );

    \I__6751\ : Odrv12
    port map (
            O => \N__40236\,
            I => encoder1_position_21
        );

    \I__6750\ : CascadeMux
    port map (
            O => \N__40227\,
            I => \N__40224\
        );

    \I__6749\ : InMux
    port map (
            O => \N__40224\,
            I => \N__40221\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__40221\,
            I => \N__40218\
        );

    \I__6747\ : Span4Mux_v
    port map (
            O => \N__40218\,
            I => \N__40215\
        );

    \I__6746\ : Sp12to4
    port map (
            O => \N__40215\,
            I => \N__40210\
        );

    \I__6745\ : InMux
    port map (
            O => \N__40214\,
            I => \N__40207\
        );

    \I__6744\ : InMux
    port map (
            O => \N__40213\,
            I => \N__40201\
        );

    \I__6743\ : Span12Mux_h
    port map (
            O => \N__40210\,
            I => \N__40196\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__40207\,
            I => \N__40196\
        );

    \I__6741\ : InMux
    port map (
            O => \N__40206\,
            I => \N__40193\
        );

    \I__6740\ : InMux
    port map (
            O => \N__40205\,
            I => \N__40188\
        );

    \I__6739\ : InMux
    port map (
            O => \N__40204\,
            I => \N__40188\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__40201\,
            I => encoder0_position_17
        );

    \I__6737\ : Odrv12
    port map (
            O => \N__40196\,
            I => encoder0_position_17
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__40193\,
            I => encoder0_position_17
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__40188\,
            I => encoder0_position_17
        );

    \I__6734\ : CascadeMux
    port map (
            O => \N__40179\,
            I => \N__40175\
        );

    \I__6733\ : InMux
    port map (
            O => \N__40178\,
            I => \N__40171\
        );

    \I__6732\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40168\
        );

    \I__6731\ : CascadeMux
    port map (
            O => \N__40174\,
            I => \N__40165\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__40171\,
            I => \N__40162\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__40168\,
            I => \N__40159\
        );

    \I__6728\ : InMux
    port map (
            O => \N__40165\,
            I => \N__40156\
        );

    \I__6727\ : Span4Mux_h
    port map (
            O => \N__40162\,
            I => \N__40153\
        );

    \I__6726\ : Span4Mux_v
    port map (
            O => \N__40159\,
            I => \N__40148\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__40156\,
            I => \N__40148\
        );

    \I__6724\ : Span4Mux_h
    port map (
            O => \N__40153\,
            I => \N__40145\
        );

    \I__6723\ : Span4Mux_v
    port map (
            O => \N__40148\,
            I => \N__40138\
        );

    \I__6722\ : Span4Mux_h
    port map (
            O => \N__40145\,
            I => \N__40138\
        );

    \I__6721\ : InMux
    port map (
            O => \N__40144\,
            I => \N__40133\
        );

    \I__6720\ : InMux
    port map (
            O => \N__40143\,
            I => \N__40133\
        );

    \I__6719\ : Odrv4
    port map (
            O => \N__40138\,
            I => encoder1_position_8
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__40133\,
            I => encoder1_position_8
        );

    \I__6717\ : InMux
    port map (
            O => \N__40128\,
            I => \N__40124\
        );

    \I__6716\ : InMux
    port map (
            O => \N__40127\,
            I => \N__40121\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__40124\,
            I => \N__40118\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__40121\,
            I => \N__40115\
        );

    \I__6713\ : Span4Mux_h
    port map (
            O => \N__40118\,
            I => \N__40112\
        );

    \I__6712\ : Span4Mux_h
    port map (
            O => \N__40115\,
            I => \N__40109\
        );

    \I__6711\ : Span4Mux_h
    port map (
            O => \N__40112\,
            I => \N__40106\
        );

    \I__6710\ : Span4Mux_v
    port map (
            O => \N__40109\,
            I => \N__40103\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__40106\,
            I => \c0.n22593\
        );

    \I__6708\ : Odrv4
    port map (
            O => \N__40103\,
            I => \c0.n22593\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__40098\,
            I => \N__40095\
        );

    \I__6706\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40091\
        );

    \I__6705\ : CascadeMux
    port map (
            O => \N__40094\,
            I => \N__40088\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__40091\,
            I => \N__40085\
        );

    \I__6703\ : InMux
    port map (
            O => \N__40088\,
            I => \N__40081\
        );

    \I__6702\ : Span4Mux_v
    port map (
            O => \N__40085\,
            I => \N__40076\
        );

    \I__6701\ : InMux
    port map (
            O => \N__40084\,
            I => \N__40073\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__40081\,
            I => \N__40070\
        );

    \I__6699\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40065\
        );

    \I__6698\ : InMux
    port map (
            O => \N__40079\,
            I => \N__40065\
        );

    \I__6697\ : Span4Mux_h
    port map (
            O => \N__40076\,
            I => \N__40059\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__40073\,
            I => \N__40059\
        );

    \I__6695\ : Span4Mux_h
    port map (
            O => \N__40070\,
            I => \N__40054\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__40065\,
            I => \N__40054\
        );

    \I__6693\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40051\
        );

    \I__6692\ : Span4Mux_v
    port map (
            O => \N__40059\,
            I => \N__40048\
        );

    \I__6691\ : Span4Mux_h
    port map (
            O => \N__40054\,
            I => \N__40045\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__40051\,
            I => encoder1_position_9
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__40048\,
            I => encoder1_position_9
        );

    \I__6688\ : Odrv4
    port map (
            O => \N__40045\,
            I => encoder1_position_9
        );

    \I__6687\ : InMux
    port map (
            O => \N__40038\,
            I => \N__40035\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__40035\,
            I => \c0.n6_adj_4276\
        );

    \I__6685\ : CascadeMux
    port map (
            O => \N__40032\,
            I => \N__40029\
        );

    \I__6684\ : InMux
    port map (
            O => \N__40029\,
            I => \N__40026\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__40026\,
            I => \N__40023\
        );

    \I__6682\ : Span4Mux_v
    port map (
            O => \N__40023\,
            I => \N__40018\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__40022\,
            I => \N__40015\
        );

    \I__6680\ : InMux
    port map (
            O => \N__40021\,
            I => \N__40012\
        );

    \I__6679\ : Span4Mux_h
    port map (
            O => \N__40018\,
            I => \N__40009\
        );

    \I__6678\ : InMux
    port map (
            O => \N__40015\,
            I => \N__40006\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__40012\,
            I => \N__40003\
        );

    \I__6676\ : Span4Mux_h
    port map (
            O => \N__40009\,
            I => \N__40000\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__40006\,
            I => \N__39995\
        );

    \I__6674\ : Span4Mux_v
    port map (
            O => \N__40003\,
            I => \N__39995\
        );

    \I__6673\ : Odrv4
    port map (
            O => \N__40000\,
            I => \c0.n22372\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__39995\,
            I => \c0.n22372\
        );

    \I__6671\ : CascadeMux
    port map (
            O => \N__39990\,
            I => \N__39986\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__39989\,
            I => \N__39983\
        );

    \I__6669\ : InMux
    port map (
            O => \N__39986\,
            I => \N__39979\
        );

    \I__6668\ : InMux
    port map (
            O => \N__39983\,
            I => \N__39976\
        );

    \I__6667\ : InMux
    port map (
            O => \N__39982\,
            I => \N__39973\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__39979\,
            I => \N__39969\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__39976\,
            I => \N__39966\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__39973\,
            I => \N__39963\
        );

    \I__6663\ : CascadeMux
    port map (
            O => \N__39972\,
            I => \N__39959\
        );

    \I__6662\ : Span4Mux_h
    port map (
            O => \N__39969\,
            I => \N__39956\
        );

    \I__6661\ : Span4Mux_h
    port map (
            O => \N__39966\,
            I => \N__39953\
        );

    \I__6660\ : Span4Mux_h
    port map (
            O => \N__39963\,
            I => \N__39950\
        );

    \I__6659\ : InMux
    port map (
            O => \N__39962\,
            I => \N__39947\
        );

    \I__6658\ : InMux
    port map (
            O => \N__39959\,
            I => \N__39944\
        );

    \I__6657\ : Span4Mux_v
    port map (
            O => \N__39956\,
            I => \N__39939\
        );

    \I__6656\ : Span4Mux_v
    port map (
            O => \N__39953\,
            I => \N__39939\
        );

    \I__6655\ : Span4Mux_v
    port map (
            O => \N__39950\,
            I => \N__39936\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__39947\,
            I => encoder1_position_28
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__39944\,
            I => encoder1_position_28
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__39939\,
            I => encoder1_position_28
        );

    \I__6651\ : Odrv4
    port map (
            O => \N__39936\,
            I => encoder1_position_28
        );

    \I__6650\ : InMux
    port map (
            O => \N__39927\,
            I => \N__39924\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__39924\,
            I => \N__39921\
        );

    \I__6648\ : Span4Mux_v
    port map (
            O => \N__39921\,
            I => \N__39918\
        );

    \I__6647\ : Odrv4
    port map (
            O => \N__39918\,
            I => \c0.n31_adj_4325\
        );

    \I__6646\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39911\
        );

    \I__6645\ : InMux
    port map (
            O => \N__39914\,
            I => \N__39908\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__39911\,
            I => \N__39905\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__39908\,
            I => \N__39902\
        );

    \I__6642\ : Span4Mux_h
    port map (
            O => \N__39905\,
            I => \N__39899\
        );

    \I__6641\ : Span4Mux_h
    port map (
            O => \N__39902\,
            I => \N__39896\
        );

    \I__6640\ : Odrv4
    port map (
            O => \N__39899\,
            I => \c0.n22775\
        );

    \I__6639\ : Odrv4
    port map (
            O => \N__39896\,
            I => \c0.n22775\
        );

    \I__6638\ : InMux
    port map (
            O => \N__39891\,
            I => \N__39888\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__39888\,
            I => n2348
        );

    \I__6636\ : InMux
    port map (
            O => \N__39885\,
            I => \N__39882\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__39882\,
            I => n2336
        );

    \I__6634\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39876\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__39876\,
            I => \N__39872\
        );

    \I__6632\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39869\
        );

    \I__6631\ : Span4Mux_h
    port map (
            O => \N__39872\,
            I => \N__39864\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__39869\,
            I => \N__39864\
        );

    \I__6629\ : Odrv4
    port map (
            O => \N__39864\,
            I => \c0.n22608\
        );

    \I__6628\ : CascadeMux
    port map (
            O => \N__39861\,
            I => \N__39858\
        );

    \I__6627\ : InMux
    port map (
            O => \N__39858\,
            I => \N__39855\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__39855\,
            I => \N__39852\
        );

    \I__6625\ : Span4Mux_h
    port map (
            O => \N__39852\,
            I => \N__39849\
        );

    \I__6624\ : Span4Mux_v
    port map (
            O => \N__39849\,
            I => \N__39845\
        );

    \I__6623\ : InMux
    port map (
            O => \N__39848\,
            I => \N__39842\
        );

    \I__6622\ : Span4Mux_v
    port map (
            O => \N__39845\,
            I => \N__39837\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__39842\,
            I => \N__39832\
        );

    \I__6620\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39829\
        );

    \I__6619\ : InMux
    port map (
            O => \N__39840\,
            I => \N__39826\
        );

    \I__6618\ : Span4Mux_v
    port map (
            O => \N__39837\,
            I => \N__39823\
        );

    \I__6617\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39820\
        );

    \I__6616\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39817\
        );

    \I__6615\ : Span4Mux_v
    port map (
            O => \N__39832\,
            I => \N__39814\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__39829\,
            I => \N__39811\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__39826\,
            I => encoder0_position_2
        );

    \I__6612\ : Odrv4
    port map (
            O => \N__39823\,
            I => encoder0_position_2
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__39820\,
            I => encoder0_position_2
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__39817\,
            I => encoder0_position_2
        );

    \I__6609\ : Odrv4
    port map (
            O => \N__39814\,
            I => encoder0_position_2
        );

    \I__6608\ : Odrv4
    port map (
            O => \N__39811\,
            I => encoder0_position_2
        );

    \I__6607\ : InMux
    port map (
            O => \N__39798\,
            I => \N__39794\
        );

    \I__6606\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39791\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__39794\,
            I => \N__39788\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__39791\,
            I => \N__39785\
        );

    \I__6603\ : Odrv4
    port map (
            O => \N__39788\,
            I => \c0.n22785\
        );

    \I__6602\ : Odrv12
    port map (
            O => \N__39785\,
            I => \c0.n22785\
        );

    \I__6601\ : InMux
    port map (
            O => \N__39780\,
            I => \N__39776\
        );

    \I__6600\ : InMux
    port map (
            O => \N__39779\,
            I => \N__39773\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__39776\,
            I => \N__39770\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__39773\,
            I => \N__39767\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__39770\,
            I => \c0.n13630\
        );

    \I__6596\ : Odrv4
    port map (
            O => \N__39767\,
            I => \c0.n13630\
        );

    \I__6595\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39759\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__39759\,
            I => n2340
        );

    \I__6593\ : InMux
    port map (
            O => \N__39756\,
            I => \N__39751\
        );

    \I__6592\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39746\
        );

    \I__6591\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39746\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__39751\,
            I => \N__39741\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__39746\,
            I => \N__39738\
        );

    \I__6588\ : InMux
    port map (
            O => \N__39745\,
            I => \N__39735\
        );

    \I__6587\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39732\
        );

    \I__6586\ : Span4Mux_h
    port map (
            O => \N__39741\,
            I => \N__39729\
        );

    \I__6585\ : Span4Mux_h
    port map (
            O => \N__39738\,
            I => \N__39726\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__39735\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__39732\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__39729\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__6581\ : Odrv4
    port map (
            O => \N__39726\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__6580\ : SRMux
    port map (
            O => \N__39717\,
            I => \N__39714\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__39714\,
            I => \N__39711\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__39711\,
            I => \N__39708\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__39708\,
            I => \c0.n21639\
        );

    \I__6576\ : CascadeMux
    port map (
            O => \N__39705\,
            I => \N__39701\
        );

    \I__6575\ : InMux
    port map (
            O => \N__39704\,
            I => \N__39698\
        );

    \I__6574\ : InMux
    port map (
            O => \N__39701\,
            I => \N__39695\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__39698\,
            I => \N__39691\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__39695\,
            I => \N__39688\
        );

    \I__6571\ : InMux
    port map (
            O => \N__39694\,
            I => \N__39685\
        );

    \I__6570\ : Span4Mux_v
    port map (
            O => \N__39691\,
            I => \N__39682\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__39688\,
            I => \N__39679\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__39685\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__6567\ : Odrv4
    port map (
            O => \N__39682\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__6566\ : Odrv4
    port map (
            O => \N__39679\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__6565\ : SRMux
    port map (
            O => \N__39672\,
            I => \N__39669\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__39669\,
            I => \N__39666\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__39666\,
            I => \N__39663\
        );

    \I__6562\ : Span4Mux_v
    port map (
            O => \N__39663\,
            I => \N__39660\
        );

    \I__6561\ : Odrv4
    port map (
            O => \N__39660\,
            I => \c0.n8_adj_4555\
        );

    \I__6560\ : SRMux
    port map (
            O => \N__39657\,
            I => \N__39654\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__39654\,
            I => \N__39651\
        );

    \I__6558\ : Span4Mux_h
    port map (
            O => \N__39651\,
            I => \N__39648\
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__39648\,
            I => \c0.n21641\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__39645\,
            I => \N__39642\
        );

    \I__6555\ : InMux
    port map (
            O => \N__39642\,
            I => \N__39639\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__39639\,
            I => \N__39636\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__39636\,
            I => \N__39633\
        );

    \I__6552\ : Span4Mux_h
    port map (
            O => \N__39633\,
            I => \N__39630\
        );

    \I__6551\ : Span4Mux_v
    port map (
            O => \N__39630\,
            I => \N__39627\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__39627\,
            I => \N__39620\
        );

    \I__6549\ : InMux
    port map (
            O => \N__39626\,
            I => \N__39617\
        );

    \I__6548\ : InMux
    port map (
            O => \N__39625\,
            I => \N__39614\
        );

    \I__6547\ : InMux
    port map (
            O => \N__39624\,
            I => \N__39609\
        );

    \I__6546\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39606\
        );

    \I__6545\ : Span4Mux_h
    port map (
            O => \N__39620\,
            I => \N__39599\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__39617\,
            I => \N__39599\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__39614\,
            I => \N__39599\
        );

    \I__6542\ : InMux
    port map (
            O => \N__39613\,
            I => \N__39596\
        );

    \I__6541\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39592\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__39609\,
            I => \N__39589\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__39606\,
            I => \N__39586\
        );

    \I__6538\ : Span4Mux_v
    port map (
            O => \N__39599\,
            I => \N__39581\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__39596\,
            I => \N__39581\
        );

    \I__6536\ : InMux
    port map (
            O => \N__39595\,
            I => \N__39578\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__39592\,
            I => encoder0_position_30
        );

    \I__6534\ : Odrv12
    port map (
            O => \N__39589\,
            I => encoder0_position_30
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__39586\,
            I => encoder0_position_30
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__39581\,
            I => encoder0_position_30
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__39578\,
            I => encoder0_position_30
        );

    \I__6530\ : InMux
    port map (
            O => \N__39567\,
            I => \N__39564\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__39564\,
            I => \N__39561\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__39561\,
            I => n2342
        );

    \I__6527\ : InMux
    port map (
            O => \N__39558\,
            I => \N__39555\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__39555\,
            I => \N__39550\
        );

    \I__6525\ : InMux
    port map (
            O => \N__39554\,
            I => \N__39546\
        );

    \I__6524\ : InMux
    port map (
            O => \N__39553\,
            I => \N__39543\
        );

    \I__6523\ : Sp12to4
    port map (
            O => \N__39550\,
            I => \N__39539\
        );

    \I__6522\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39536\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__39546\,
            I => \N__39533\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__39543\,
            I => \N__39530\
        );

    \I__6519\ : InMux
    port map (
            O => \N__39542\,
            I => \N__39526\
        );

    \I__6518\ : Span12Mux_v
    port map (
            O => \N__39539\,
            I => \N__39521\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__39536\,
            I => \N__39521\
        );

    \I__6516\ : Span4Mux_v
    port map (
            O => \N__39533\,
            I => \N__39516\
        );

    \I__6515\ : Span4Mux_h
    port map (
            O => \N__39530\,
            I => \N__39516\
        );

    \I__6514\ : InMux
    port map (
            O => \N__39529\,
            I => \N__39513\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__39526\,
            I => encoder0_position_15
        );

    \I__6512\ : Odrv12
    port map (
            O => \N__39521\,
            I => encoder0_position_15
        );

    \I__6511\ : Odrv4
    port map (
            O => \N__39516\,
            I => encoder0_position_15
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__39513\,
            I => encoder0_position_15
        );

    \I__6509\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39501\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__39501\,
            I => n2352
        );

    \I__6507\ : CascadeMux
    port map (
            O => \N__39498\,
            I => \c0.n30_adj_4730_cascade_\
        );

    \I__6506\ : InMux
    port map (
            O => \N__39495\,
            I => \N__39492\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__39492\,
            I => \N__39489\
        );

    \I__6504\ : Span4Mux_h
    port map (
            O => \N__39489\,
            I => \N__39485\
        );

    \I__6503\ : InMux
    port map (
            O => \N__39488\,
            I => \N__39482\
        );

    \I__6502\ : Span4Mux_v
    port map (
            O => \N__39485\,
            I => \N__39479\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__39482\,
            I => \N__39476\
        );

    \I__6500\ : Span4Mux_v
    port map (
            O => \N__39479\,
            I => \N__39473\
        );

    \I__6499\ : Span12Mux_v
    port map (
            O => \N__39476\,
            I => \N__39470\
        );

    \I__6498\ : Odrv4
    port map (
            O => \N__39473\,
            I => \c0.n17539\
        );

    \I__6497\ : Odrv12
    port map (
            O => \N__39470\,
            I => \c0.n17539\
        );

    \I__6496\ : InMux
    port map (
            O => \N__39465\,
            I => \N__39462\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__39462\,
            I => \N__39459\
        );

    \I__6494\ : Span4Mux_v
    port map (
            O => \N__39459\,
            I => \N__39455\
        );

    \I__6493\ : CascadeMux
    port map (
            O => \N__39458\,
            I => \N__39452\
        );

    \I__6492\ : Span4Mux_h
    port map (
            O => \N__39455\,
            I => \N__39448\
        );

    \I__6491\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39445\
        );

    \I__6490\ : InMux
    port map (
            O => \N__39451\,
            I => \N__39442\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__39448\,
            I => \N__39434\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__39445\,
            I => \N__39434\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__39442\,
            I => \N__39434\
        );

    \I__6486\ : InMux
    port map (
            O => \N__39441\,
            I => \N__39431\
        );

    \I__6485\ : Span4Mux_v
    port map (
            O => \N__39434\,
            I => \N__39428\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__39431\,
            I => \c0.n17846\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__39428\,
            I => \c0.n17846\
        );

    \I__6482\ : InMux
    port map (
            O => \N__39423\,
            I => \N__39418\
        );

    \I__6481\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39413\
        );

    \I__6480\ : InMux
    port map (
            O => \N__39421\,
            I => \N__39413\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__39418\,
            I => \N__39407\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__39413\,
            I => \N__39407\
        );

    \I__6477\ : InMux
    port map (
            O => \N__39412\,
            I => \N__39404\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__39407\,
            I => \c0.n4_adj_4654\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__39404\,
            I => \c0.n4_adj_4654\
        );

    \I__6474\ : CascadeMux
    port map (
            O => \N__39399\,
            I => \N__39396\
        );

    \I__6473\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39393\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__39393\,
            I => \N__39389\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__39392\,
            I => \N__39386\
        );

    \I__6470\ : Span4Mux_h
    port map (
            O => \N__39389\,
            I => \N__39383\
        );

    \I__6469\ : InMux
    port map (
            O => \N__39386\,
            I => \N__39380\
        );

    \I__6468\ : Odrv4
    port map (
            O => \N__39383\,
            I => \c0.n17533\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__39380\,
            I => \c0.n17533\
        );

    \I__6466\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39372\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39367\
        );

    \I__6464\ : InMux
    port map (
            O => \N__39371\,
            I => \N__39364\
        );

    \I__6463\ : InMux
    port map (
            O => \N__39370\,
            I => \N__39361\
        );

    \I__6462\ : Span4Mux_h
    port map (
            O => \N__39367\,
            I => \N__39358\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__39364\,
            I => \N__39353\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__39361\,
            I => \N__39353\
        );

    \I__6459\ : Odrv4
    port map (
            O => \N__39358\,
            I => \c0.n22907\
        );

    \I__6458\ : Odrv12
    port map (
            O => \N__39353\,
            I => \c0.n22907\
        );

    \I__6457\ : InMux
    port map (
            O => \N__39348\,
            I => \N__39345\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__39345\,
            I => \N__39342\
        );

    \I__6455\ : Odrv4
    port map (
            O => \N__39342\,
            I => \c0.n24422\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__39339\,
            I => \c0.n24596_cascade_\
        );

    \I__6453\ : InMux
    port map (
            O => \N__39336\,
            I => \N__39330\
        );

    \I__6452\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39327\
        );

    \I__6451\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39322\
        );

    \I__6450\ : InMux
    port map (
            O => \N__39333\,
            I => \N__39322\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__39330\,
            I => \c0.n2004\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__39327\,
            I => \c0.n2004\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__39322\,
            I => \c0.n2004\
        );

    \I__6446\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39311\
        );

    \I__6445\ : InMux
    port map (
            O => \N__39314\,
            I => \N__39308\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__39311\,
            I => \N__39305\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__39308\,
            I => \N__39302\
        );

    \I__6442\ : Span12Mux_s10_h
    port map (
            O => \N__39305\,
            I => \N__39297\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__39302\,
            I => \N__39294\
        );

    \I__6440\ : InMux
    port map (
            O => \N__39301\,
            I => \N__39289\
        );

    \I__6439\ : InMux
    port map (
            O => \N__39300\,
            I => \N__39289\
        );

    \I__6438\ : Odrv12
    port map (
            O => \N__39297\,
            I => \c0.rx.r_SM_Main_2_N_3686_0\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__39294\,
            I => \c0.rx.r_SM_Main_2_N_3686_0\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__39289\,
            I => \c0.rx.r_SM_Main_2_N_3686_0\
        );

    \I__6435\ : CascadeMux
    port map (
            O => \N__39282\,
            I => \c0.rx.n6_cascade_\
        );

    \I__6434\ : CEMux
    port map (
            O => \N__39279\,
            I => \N__39276\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__39276\,
            I => \N__39272\
        );

    \I__6432\ : InMux
    port map (
            O => \N__39275\,
            I => \N__39269\
        );

    \I__6431\ : Span12Mux_h
    port map (
            O => \N__39272\,
            I => \N__39266\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__39269\,
            I => \N__39263\
        );

    \I__6429\ : Odrv12
    port map (
            O => \N__39266\,
            I => n14439
        );

    \I__6428\ : Odrv12
    port map (
            O => \N__39263\,
            I => n14439
        );

    \I__6427\ : InMux
    port map (
            O => \N__39258\,
            I => \N__39254\
        );

    \I__6426\ : InMux
    port map (
            O => \N__39257\,
            I => \N__39251\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__39254\,
            I => \N__39247\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__39251\,
            I => \N__39244\
        );

    \I__6423\ : InMux
    port map (
            O => \N__39250\,
            I => \N__39241\
        );

    \I__6422\ : Span4Mux_v
    port map (
            O => \N__39247\,
            I => \N__39237\
        );

    \I__6421\ : Span4Mux_h
    port map (
            O => \N__39244\,
            I => \N__39234\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__39241\,
            I => \N__39231\
        );

    \I__6419\ : InMux
    port map (
            O => \N__39240\,
            I => \N__39228\
        );

    \I__6418\ : Odrv4
    port map (
            O => \N__39237\,
            I => \c0.n7570\
        );

    \I__6417\ : Odrv4
    port map (
            O => \N__39234\,
            I => \c0.n7570\
        );

    \I__6416\ : Odrv12
    port map (
            O => \N__39231\,
            I => \c0.n7570\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__39228\,
            I => \c0.n7570\
        );

    \I__6414\ : InMux
    port map (
            O => \N__39219\,
            I => \N__39216\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__39216\,
            I => \N__39213\
        );

    \I__6412\ : Odrv4
    port map (
            O => \N__39213\,
            I => \c0.n24386\
        );

    \I__6411\ : CascadeMux
    port map (
            O => \N__39210\,
            I => \c0.n24302_cascade_\
        );

    \I__6410\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39203\
        );

    \I__6409\ : InMux
    port map (
            O => \N__39206\,
            I => \N__39199\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__39203\,
            I => \N__39196\
        );

    \I__6407\ : InMux
    port map (
            O => \N__39202\,
            I => \N__39193\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__39199\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__39196\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__39193\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__6403\ : SRMux
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__6401\ : Span4Mux_h
    port map (
            O => \N__39180\,
            I => \N__39177\
        );

    \I__6400\ : Span4Mux_h
    port map (
            O => \N__39177\,
            I => \N__39174\
        );

    \I__6399\ : Odrv4
    port map (
            O => \N__39174\,
            I => \c0.n8_adj_4556\
        );

    \I__6398\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39165\
        );

    \I__6397\ : InMux
    port map (
            O => \N__39170\,
            I => \N__39162\
        );

    \I__6396\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39157\
        );

    \I__6395\ : InMux
    port map (
            O => \N__39168\,
            I => \N__39157\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__39165\,
            I => \N__39154\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__39162\,
            I => \N__39151\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__39157\,
            I => data_in_3_5
        );

    \I__6391\ : Odrv4
    port map (
            O => \N__39154\,
            I => data_in_3_5
        );

    \I__6390\ : Odrv12
    port map (
            O => \N__39151\,
            I => data_in_3_5
        );

    \I__6389\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39140\
        );

    \I__6388\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39137\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__39140\,
            I => \N__39134\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__39137\,
            I => \N__39129\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__39134\,
            I => \N__39129\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__39129\,
            I => \N__39126\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__39126\,
            I => \c0.n13063\
        );

    \I__6382\ : CascadeMux
    port map (
            O => \N__39123\,
            I => \c0.n13063_cascade_\
        );

    \I__6381\ : InMux
    port map (
            O => \N__39120\,
            I => \N__39117\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__39117\,
            I => \c0.n6_adj_4263\
        );

    \I__6379\ : InMux
    port map (
            O => \N__39114\,
            I => \N__39103\
        );

    \I__6378\ : InMux
    port map (
            O => \N__39113\,
            I => \N__39103\
        );

    \I__6377\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39098\
        );

    \I__6376\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39098\
        );

    \I__6375\ : InMux
    port map (
            O => \N__39110\,
            I => \N__39094\
        );

    \I__6374\ : InMux
    port map (
            O => \N__39109\,
            I => \N__39091\
        );

    \I__6373\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39085\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__39103\,
            I => \N__39080\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__39098\,
            I => \N__39080\
        );

    \I__6370\ : InMux
    port map (
            O => \N__39097\,
            I => \N__39077\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__39094\,
            I => \N__39072\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__39091\,
            I => \N__39072\
        );

    \I__6367\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39068\
        );

    \I__6366\ : InMux
    port map (
            O => \N__39089\,
            I => \N__39063\
        );

    \I__6365\ : InMux
    port map (
            O => \N__39088\,
            I => \N__39063\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__39085\,
            I => \N__39056\
        );

    \I__6363\ : Span4Mux_v
    port map (
            O => \N__39080\,
            I => \N__39056\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__39077\,
            I => \N__39056\
        );

    \I__6361\ : Span4Mux_h
    port map (
            O => \N__39072\,
            I => \N__39053\
        );

    \I__6360\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39050\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__39068\,
            I => \c0.n9706\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__39063\,
            I => \c0.n9706\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__39056\,
            I => \c0.n9706\
        );

    \I__6356\ : Odrv4
    port map (
            O => \N__39053\,
            I => \c0.n9706\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__39050\,
            I => \c0.n9706\
        );

    \I__6354\ : InMux
    port map (
            O => \N__39039\,
            I => \N__39035\
        );

    \I__6353\ : InMux
    port map (
            O => \N__39038\,
            I => \N__39032\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__39035\,
            I => \N__39029\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__39032\,
            I => \N__39026\
        );

    \I__6350\ : Span4Mux_v
    port map (
            O => \N__39029\,
            I => \N__39021\
        );

    \I__6349\ : Span4Mux_v
    port map (
            O => \N__39026\,
            I => \N__39021\
        );

    \I__6348\ : Span4Mux_h
    port map (
            O => \N__39021\,
            I => \N__39017\
        );

    \I__6347\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39014\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__39017\,
            I => \c0.n3325\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__39014\,
            I => \c0.n3325\
        );

    \I__6344\ : InMux
    port map (
            O => \N__39009\,
            I => \N__39004\
        );

    \I__6343\ : InMux
    port map (
            O => \N__39008\,
            I => \N__39001\
        );

    \I__6342\ : InMux
    port map (
            O => \N__39007\,
            I => \N__38998\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__39004\,
            I => \N__38995\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__39001\,
            I => data_in_2_7
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__38998\,
            I => data_in_2_7
        );

    \I__6338\ : Odrv12
    port map (
            O => \N__38995\,
            I => data_in_2_7
        );

    \I__6337\ : InMux
    port map (
            O => \N__38988\,
            I => \N__38982\
        );

    \I__6336\ : InMux
    port map (
            O => \N__38987\,
            I => \N__38982\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__38982\,
            I => \N__38978\
        );

    \I__6334\ : InMux
    port map (
            O => \N__38981\,
            I => \N__38975\
        );

    \I__6333\ : Sp12to4
    port map (
            O => \N__38978\,
            I => \N__38972\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__38975\,
            I => data_in_1_7
        );

    \I__6331\ : Odrv12
    port map (
            O => \N__38972\,
            I => data_in_1_7
        );

    \I__6330\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38961\
        );

    \I__6329\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38961\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__38961\,
            I => \N__38958\
        );

    \I__6327\ : Odrv4
    port map (
            O => \N__38958\,
            I => \c0.n17682\
        );

    \I__6326\ : InMux
    port map (
            O => \N__38955\,
            I => \N__38948\
        );

    \I__6325\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38935\
        );

    \I__6324\ : InMux
    port map (
            O => \N__38953\,
            I => \N__38935\
        );

    \I__6323\ : InMux
    port map (
            O => \N__38952\,
            I => \N__38935\
        );

    \I__6322\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38935\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__38948\,
            I => \N__38930\
        );

    \I__6320\ : InMux
    port map (
            O => \N__38947\,
            I => \N__38921\
        );

    \I__6319\ : InMux
    port map (
            O => \N__38946\,
            I => \N__38921\
        );

    \I__6318\ : InMux
    port map (
            O => \N__38945\,
            I => \N__38921\
        );

    \I__6317\ : InMux
    port map (
            O => \N__38944\,
            I => \N__38921\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__38935\,
            I => \N__38918\
        );

    \I__6315\ : InMux
    port map (
            O => \N__38934\,
            I => \N__38915\
        );

    \I__6314\ : InMux
    port map (
            O => \N__38933\,
            I => \N__38910\
        );

    \I__6313\ : Span4Mux_v
    port map (
            O => \N__38930\,
            I => \N__38905\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__38921\,
            I => \N__38905\
        );

    \I__6311\ : Span4Mux_h
    port map (
            O => \N__38918\,
            I => \N__38900\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__38915\,
            I => \N__38900\
        );

    \I__6309\ : InMux
    port map (
            O => \N__38914\,
            I => \N__38895\
        );

    \I__6308\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38895\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__38910\,
            I => \c0.n1\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__38905\,
            I => \c0.n1\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__38900\,
            I => \c0.n1\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__38895\,
            I => \c0.n1\
        );

    \I__6303\ : InMux
    port map (
            O => \N__38886\,
            I => \N__38883\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__38883\,
            I => \c0.n24745\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__38880\,
            I => \N__38876\
        );

    \I__6300\ : InMux
    port map (
            O => \N__38879\,
            I => \N__38872\
        );

    \I__6299\ : InMux
    port map (
            O => \N__38876\,
            I => \N__38869\
        );

    \I__6298\ : InMux
    port map (
            O => \N__38875\,
            I => \N__38865\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__38872\,
            I => \N__38860\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__38869\,
            I => \N__38860\
        );

    \I__6295\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38857\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__38865\,
            I => \N__38852\
        );

    \I__6293\ : Span4Mux_v
    port map (
            O => \N__38860\,
            I => \N__38852\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__38857\,
            I => data_in_2_6
        );

    \I__6291\ : Odrv4
    port map (
            O => \N__38852\,
            I => data_in_2_6
        );

    \I__6290\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38842\
        );

    \I__6289\ : InMux
    port map (
            O => \N__38846\,
            I => \N__38839\
        );

    \I__6288\ : InMux
    port map (
            O => \N__38845\,
            I => \N__38836\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__38842\,
            I => data_in_0_5
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__38839\,
            I => data_in_0_5
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__38836\,
            I => data_in_0_5
        );

    \I__6284\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38826\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__38826\,
            I => \c0.n17_adj_4232\
        );

    \I__6282\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38820\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__38820\,
            I => \N__38817\
        );

    \I__6280\ : Span4Mux_v
    port map (
            O => \N__38817\,
            I => \N__38814\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__38814\,
            I => n2261
        );

    \I__6278\ : CascadeMux
    port map (
            O => \N__38811\,
            I => \N__38805\
        );

    \I__6277\ : InMux
    port map (
            O => \N__38810\,
            I => \N__38802\
        );

    \I__6276\ : InMux
    port map (
            O => \N__38809\,
            I => \N__38799\
        );

    \I__6275\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38796\
        );

    \I__6274\ : InMux
    port map (
            O => \N__38805\,
            I => \N__38793\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__38802\,
            I => \N__38788\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38788\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__38796\,
            I => \N__38782\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__38793\,
            I => \N__38782\
        );

    \I__6269\ : Span12Mux_h
    port map (
            O => \N__38788\,
            I => \N__38779\
        );

    \I__6268\ : InMux
    port map (
            O => \N__38787\,
            I => \N__38776\
        );

    \I__6267\ : Span4Mux_h
    port map (
            O => \N__38782\,
            I => \N__38773\
        );

    \I__6266\ : Span12Mux_v
    port map (
            O => \N__38779\,
            I => \N__38770\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__38776\,
            I => encoder1_position_30
        );

    \I__6264\ : Odrv4
    port map (
            O => \N__38773\,
            I => encoder1_position_30
        );

    \I__6263\ : Odrv12
    port map (
            O => \N__38770\,
            I => encoder1_position_30
        );

    \I__6262\ : InMux
    port map (
            O => \N__38763\,
            I => \N__38758\
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__38762\,
            I => \N__38755\
        );

    \I__6260\ : InMux
    port map (
            O => \N__38761\,
            I => \N__38751\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__38758\,
            I => \N__38748\
        );

    \I__6258\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38743\
        );

    \I__6257\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38743\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__38751\,
            I => data_in_3_7
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__38748\,
            I => data_in_3_7
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__38743\,
            I => data_in_3_7
        );

    \I__6253\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38731\
        );

    \I__6252\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38728\
        );

    \I__6251\ : InMux
    port map (
            O => \N__38734\,
            I => \N__38725\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__38731\,
            I => \N__38722\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__38728\,
            I => \N__38719\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__38725\,
            I => \N__38713\
        );

    \I__6247\ : Span4Mux_h
    port map (
            O => \N__38722\,
            I => \N__38713\
        );

    \I__6246\ : Span4Mux_h
    port map (
            O => \N__38719\,
            I => \N__38710\
        );

    \I__6245\ : InMux
    port map (
            O => \N__38718\,
            I => \N__38707\
        );

    \I__6244\ : Span4Mux_v
    port map (
            O => \N__38713\,
            I => \N__38704\
        );

    \I__6243\ : Odrv4
    port map (
            O => \N__38710\,
            I => data_in_2_2
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__38707\,
            I => data_in_2_2
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__38704\,
            I => data_in_2_2
        );

    \I__6240\ : CascadeMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__6239\ : InMux
    port map (
            O => \N__38694\,
            I => \N__38688\
        );

    \I__6238\ : InMux
    port map (
            O => \N__38693\,
            I => \N__38688\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__38688\,
            I => data_out_frame_8_1
        );

    \I__6236\ : CascadeMux
    port map (
            O => \N__38685\,
            I => \N__38682\
        );

    \I__6235\ : InMux
    port map (
            O => \N__38682\,
            I => \N__38679\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__6233\ : Span4Mux_h
    port map (
            O => \N__38676\,
            I => \N__38670\
        );

    \I__6232\ : InMux
    port map (
            O => \N__38675\,
            I => \N__38667\
        );

    \I__6231\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38664\
        );

    \I__6230\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38661\
        );

    \I__6229\ : Span4Mux_v
    port map (
            O => \N__38670\,
            I => \N__38658\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__38667\,
            I => encoder1_position_29
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__38664\,
            I => encoder1_position_29
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__38661\,
            I => encoder1_position_29
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__38658\,
            I => encoder1_position_29
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__38649\,
            I => \N__38645\
        );

    \I__6223\ : InMux
    port map (
            O => \N__38648\,
            I => \N__38642\
        );

    \I__6222\ : InMux
    port map (
            O => \N__38645\,
            I => \N__38639\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__38642\,
            I => \N__38636\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__38639\,
            I => data_out_frame_10_5
        );

    \I__6219\ : Odrv12
    port map (
            O => \N__38636\,
            I => data_out_frame_10_5
        );

    \I__6218\ : InMux
    port map (
            O => \N__38631\,
            I => \N__38627\
        );

    \I__6217\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38624\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__38627\,
            I => \N__38619\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__38624\,
            I => \N__38619\
        );

    \I__6214\ : Odrv12
    port map (
            O => \N__38619\,
            I => \c0.n13046\
        );

    \I__6213\ : InMux
    port map (
            O => \N__38616\,
            I => \N__38613\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__38613\,
            I => \N__38609\
        );

    \I__6211\ : InMux
    port map (
            O => \N__38612\,
            I => \N__38606\
        );

    \I__6210\ : Span4Mux_v
    port map (
            O => \N__38609\,
            I => \N__38601\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__38606\,
            I => \N__38601\
        );

    \I__6208\ : Odrv4
    port map (
            O => \N__38601\,
            I => \c0.n12898\
        );

    \I__6207\ : CascadeMux
    port map (
            O => \N__38598\,
            I => \c0.n20_adj_4308_cascade_\
        );

    \I__6206\ : InMux
    port map (
            O => \N__38595\,
            I => \N__38592\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__38592\,
            I => \c0.n19_adj_4307\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__38589\,
            I => \c0.n16_adj_4231_cascade_\
        );

    \I__6203\ : CascadeMux
    port map (
            O => \N__38586\,
            I => \N__38582\
        );

    \I__6202\ : InMux
    port map (
            O => \N__38585\,
            I => \N__38579\
        );

    \I__6201\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38576\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__38579\,
            I => \N__38571\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__38576\,
            I => \N__38571\
        );

    \I__6198\ : Odrv12
    port map (
            O => \N__38571\,
            I => \c0.n12986\
        );

    \I__6197\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38565\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__38565\,
            I => \c0.n17_adj_4234\
        );

    \I__6195\ : InMux
    port map (
            O => \N__38562\,
            I => \N__38559\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__38559\,
            I => \N__38556\
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__38556\,
            I => n2268
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__38553\,
            I => \N__38548\
        );

    \I__6191\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38543\
        );

    \I__6190\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38543\
        );

    \I__6189\ : InMux
    port map (
            O => \N__38548\,
            I => \N__38539\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__38543\,
            I => \N__38536\
        );

    \I__6187\ : InMux
    port map (
            O => \N__38542\,
            I => \N__38532\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__38539\,
            I => \N__38529\
        );

    \I__6185\ : Span4Mux_h
    port map (
            O => \N__38536\,
            I => \N__38526\
        );

    \I__6184\ : InMux
    port map (
            O => \N__38535\,
            I => \N__38523\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__38532\,
            I => \N__38520\
        );

    \I__6182\ : Span4Mux_v
    port map (
            O => \N__38529\,
            I => \N__38515\
        );

    \I__6181\ : Span4Mux_v
    port map (
            O => \N__38526\,
            I => \N__38515\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__38523\,
            I => encoder1_position_23
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__38520\,
            I => encoder1_position_23
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__38515\,
            I => encoder1_position_23
        );

    \I__6177\ : InMux
    port map (
            O => \N__38508\,
            I => \N__38505\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__38505\,
            I => \N__38502\
        );

    \I__6175\ : Span4Mux_v
    port map (
            O => \N__38502\,
            I => \N__38499\
        );

    \I__6174\ : Span4Mux_v
    port map (
            O => \N__38499\,
            I => \N__38496\
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__38496\,
            I => n2344
        );

    \I__6172\ : InMux
    port map (
            O => \N__38493\,
            I => \N__38490\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__38490\,
            I => \N__38487\
        );

    \I__6170\ : Odrv12
    port map (
            O => \N__38487\,
            I => \c0.n10_adj_4240\
        );

    \I__6169\ : CEMux
    port map (
            O => \N__38484\,
            I => \N__38479\
        );

    \I__6168\ : CEMux
    port map (
            O => \N__38483\,
            I => \N__38475\
        );

    \I__6167\ : InMux
    port map (
            O => \N__38482\,
            I => \N__38472\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__38479\,
            I => \N__38468\
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__38478\,
            I => \N__38464\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__38475\,
            I => \N__38460\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__38472\,
            I => \N__38457\
        );

    \I__6162\ : InMux
    port map (
            O => \N__38471\,
            I => \N__38454\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__38468\,
            I => \N__38451\
        );

    \I__6160\ : InMux
    port map (
            O => \N__38467\,
            I => \N__38446\
        );

    \I__6159\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38446\
        );

    \I__6158\ : InMux
    port map (
            O => \N__38463\,
            I => \N__38443\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__38460\,
            I => \N__38438\
        );

    \I__6156\ : Span4Mux_v
    port map (
            O => \N__38457\,
            I => \N__38438\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__38454\,
            I => \N__38435\
        );

    \I__6154\ : Span4Mux_h
    port map (
            O => \N__38451\,
            I => \N__38430\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__38446\,
            I => \N__38430\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__38443\,
            I => \N__38427\
        );

    \I__6151\ : Span4Mux_h
    port map (
            O => \N__38438\,
            I => \N__38420\
        );

    \I__6150\ : Span4Mux_v
    port map (
            O => \N__38435\,
            I => \N__38420\
        );

    \I__6149\ : Span4Mux_v
    port map (
            O => \N__38430\,
            I => \N__38420\
        );

    \I__6148\ : Odrv4
    port map (
            O => \N__38427\,
            I => n14374
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__38420\,
            I => n14374
        );

    \I__6146\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38412\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__38412\,
            I => \N__38409\
        );

    \I__6144\ : Span4Mux_h
    port map (
            O => \N__38409\,
            I => \N__38406\
        );

    \I__6143\ : Span4Mux_h
    port map (
            O => \N__38406\,
            I => \N__38403\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__38403\,
            I => \c0.tx.n24889\
        );

    \I__6141\ : InMux
    port map (
            O => \N__38400\,
            I => \N__38397\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__38397\,
            I => \N__38394\
        );

    \I__6139\ : Span4Mux_v
    port map (
            O => \N__38394\,
            I => \N__38390\
        );

    \I__6138\ : InMux
    port map (
            O => \N__38393\,
            I => \N__38387\
        );

    \I__6137\ : Sp12to4
    port map (
            O => \N__38390\,
            I => \N__38384\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__38387\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__6135\ : Odrv12
    port map (
            O => \N__38384\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__6134\ : InMux
    port map (
            O => \N__38379\,
            I => \N__38376\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__38376\,
            I => \N__38373\
        );

    \I__6132\ : Span4Mux_h
    port map (
            O => \N__38373\,
            I => \N__38370\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__38370\,
            I => n2265
        );

    \I__6130\ : CascadeMux
    port map (
            O => \N__38367\,
            I => \N__38362\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__38366\,
            I => \N__38359\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__38365\,
            I => \N__38356\
        );

    \I__6127\ : InMux
    port map (
            O => \N__38362\,
            I => \N__38353\
        );

    \I__6126\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38350\
        );

    \I__6125\ : InMux
    port map (
            O => \N__38356\,
            I => \N__38347\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__38353\,
            I => \N__38344\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__38350\,
            I => \N__38338\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__38347\,
            I => \N__38338\
        );

    \I__6121\ : Span4Mux_h
    port map (
            O => \N__38344\,
            I => \N__38335\
        );

    \I__6120\ : InMux
    port map (
            O => \N__38343\,
            I => \N__38332\
        );

    \I__6119\ : Span4Mux_v
    port map (
            O => \N__38338\,
            I => \N__38329\
        );

    \I__6118\ : Span4Mux_v
    port map (
            O => \N__38335\,
            I => \N__38326\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__38332\,
            I => encoder1_position_26
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__38329\,
            I => encoder1_position_26
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__38326\,
            I => encoder1_position_26
        );

    \I__6114\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38315\
        );

    \I__6113\ : InMux
    port map (
            O => \N__38318\,
            I => \N__38312\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__38315\,
            I => data_out_frame_10_1
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__38312\,
            I => data_out_frame_10_1
        );

    \I__6110\ : CascadeMux
    port map (
            O => \N__38307\,
            I => \N__38303\
        );

    \I__6109\ : InMux
    port map (
            O => \N__38306\,
            I => \N__38300\
        );

    \I__6108\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38297\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__38300\,
            I => data_out_frame_11_1
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__38297\,
            I => data_out_frame_11_1
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__38292\,
            I => \c0.n25116_cascade_\
        );

    \I__6104\ : InMux
    port map (
            O => \N__38289\,
            I => \N__38285\
        );

    \I__6103\ : InMux
    port map (
            O => \N__38288\,
            I => \N__38282\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__38285\,
            I => \N__38279\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__38282\,
            I => data_out_frame_9_1
        );

    \I__6100\ : Odrv4
    port map (
            O => \N__38279\,
            I => data_out_frame_9_1
        );

    \I__6099\ : InMux
    port map (
            O => \N__38274\,
            I => \N__38271\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__38271\,
            I => \N__38268\
        );

    \I__6097\ : Odrv12
    port map (
            O => \N__38268\,
            I => \c0.n25119\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__38265\,
            I => \N__38259\
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__38264\,
            I => \N__38255\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__38263\,
            I => \N__38251\
        );

    \I__6093\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38248\
        );

    \I__6092\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38245\
        );

    \I__6091\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38242\
        );

    \I__6090\ : InMux
    port map (
            O => \N__38255\,
            I => \N__38239\
        );

    \I__6089\ : InMux
    port map (
            O => \N__38254\,
            I => \N__38234\
        );

    \I__6088\ : InMux
    port map (
            O => \N__38251\,
            I => \N__38234\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38229\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__38245\,
            I => \N__38229\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__38242\,
            I => \N__38223\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__38239\,
            I => \N__38220\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__38234\,
            I => \N__38217\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__38229\,
            I => \N__38214\
        );

    \I__6081\ : InMux
    port map (
            O => \N__38228\,
            I => \N__38209\
        );

    \I__6080\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38209\
        );

    \I__6079\ : InMux
    port map (
            O => \N__38226\,
            I => \N__38206\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__38223\,
            I => \N__38203\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__38220\,
            I => \c0.n22291\
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__38217\,
            I => \c0.n22291\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__38214\,
            I => \c0.n22291\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__38209\,
            I => \c0.n22291\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__38206\,
            I => \c0.n22291\
        );

    \I__6072\ : Odrv4
    port map (
            O => \N__38203\,
            I => \c0.n22291\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__38190\,
            I => \N__38186\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__38189\,
            I => \N__38181\
        );

    \I__6069\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38169\
        );

    \I__6068\ : InMux
    port map (
            O => \N__38185\,
            I => \N__38169\
        );

    \I__6067\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38166\
        );

    \I__6066\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38155\
        );

    \I__6065\ : InMux
    port map (
            O => \N__38180\,
            I => \N__38155\
        );

    \I__6064\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38155\
        );

    \I__6063\ : InMux
    port map (
            O => \N__38178\,
            I => \N__38155\
        );

    \I__6062\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38150\
        );

    \I__6061\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38150\
        );

    \I__6060\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38147\
        );

    \I__6059\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38144\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__38169\,
            I => \N__38139\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__38166\,
            I => \N__38139\
        );

    \I__6056\ : InMux
    port map (
            O => \N__38165\,
            I => \N__38134\
        );

    \I__6055\ : InMux
    port map (
            O => \N__38164\,
            I => \N__38134\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__38155\,
            I => \N__38129\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__38150\,
            I => \N__38129\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__38147\,
            I => \N__38126\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__38144\,
            I => \N__38123\
        );

    \I__6050\ : Span4Mux_v
    port map (
            O => \N__38139\,
            I => \N__38115\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__38134\,
            I => \N__38115\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__38129\,
            I => \N__38115\
        );

    \I__6047\ : Span4Mux_v
    port map (
            O => \N__38126\,
            I => \N__38112\
        );

    \I__6046\ : Span12Mux_s11_h
    port map (
            O => \N__38123\,
            I => \N__38109\
        );

    \I__6045\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38106\
        );

    \I__6044\ : Span4Mux_v
    port map (
            O => \N__38115\,
            I => \N__38101\
        );

    \I__6043\ : Span4Mux_v
    port map (
            O => \N__38112\,
            I => \N__38101\
        );

    \I__6042\ : Odrv12
    port map (
            O => \N__38109\,
            I => \c0.n20333\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__38106\,
            I => \c0.n20333\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__38101\,
            I => \c0.n20333\
        );

    \I__6039\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38084\
        );

    \I__6038\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38084\
        );

    \I__6037\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38077\
        );

    \I__6036\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38077\
        );

    \I__6035\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38072\
        );

    \I__6034\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38072\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__38084\,
            I => \N__38069\
        );

    \I__6032\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38066\
        );

    \I__6031\ : InMux
    port map (
            O => \N__38082\,
            I => \N__38063\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__38077\,
            I => \N__38060\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__38072\,
            I => \N__38052\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__38069\,
            I => \N__38052\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__38066\,
            I => \N__38052\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__38063\,
            I => \N__38049\
        );

    \I__6025\ : Span4Mux_h
    port map (
            O => \N__38060\,
            I => \N__38046\
        );

    \I__6024\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38043\
        );

    \I__6023\ : Span4Mux_v
    port map (
            O => \N__38052\,
            I => \N__38038\
        );

    \I__6022\ : Span4Mux_v
    port map (
            O => \N__38049\,
            I => \N__38038\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__38046\,
            I => \c0.data_out_frame_29__7__N_1148\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__38043\,
            I => \c0.data_out_frame_29__7__N_1148\
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__38038\,
            I => \c0.data_out_frame_29__7__N_1148\
        );

    \I__6018\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38026\
        );

    \I__6017\ : InMux
    port map (
            O => \N__38030\,
            I => \N__38022\
        );

    \I__6016\ : InMux
    port map (
            O => \N__38029\,
            I => \N__38018\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__38015\
        );

    \I__6014\ : InMux
    port map (
            O => \N__38025\,
            I => \N__38012\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__38022\,
            I => \N__38007\
        );

    \I__6012\ : InMux
    port map (
            O => \N__38021\,
            I => \N__38003\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__38018\,
            I => \N__38000\
        );

    \I__6010\ : Span4Mux_v
    port map (
            O => \N__38015\,
            I => \N__37995\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__38012\,
            I => \N__37995\
        );

    \I__6008\ : InMux
    port map (
            O => \N__38011\,
            I => \N__37990\
        );

    \I__6007\ : InMux
    port map (
            O => \N__38010\,
            I => \N__37990\
        );

    \I__6006\ : Span4Mux_h
    port map (
            O => \N__38007\,
            I => \N__37987\
        );

    \I__6005\ : InMux
    port map (
            O => \N__38006\,
            I => \N__37984\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__38003\,
            I => \N__37979\
        );

    \I__6003\ : Span4Mux_h
    port map (
            O => \N__38000\,
            I => \N__37979\
        );

    \I__6002\ : Span4Mux_h
    port map (
            O => \N__37995\,
            I => \N__37976\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__37990\,
            I => \N__37973\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__37987\,
            I => \c0.n21464\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__37984\,
            I => \c0.n21464\
        );

    \I__5998\ : Odrv4
    port map (
            O => \N__37979\,
            I => \c0.n21464\
        );

    \I__5997\ : Odrv4
    port map (
            O => \N__37976\,
            I => \c0.n21464\
        );

    \I__5996\ : Odrv12
    port map (
            O => \N__37973\,
            I => \c0.n21464\
        );

    \I__5995\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37959\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__37959\,
            I => \N__37956\
        );

    \I__5993\ : Span4Mux_v
    port map (
            O => \N__37956\,
            I => \N__37953\
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__37953\,
            I => n2267
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__37950\,
            I => \N__37947\
        );

    \I__5990\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37943\
        );

    \I__5989\ : CascadeMux
    port map (
            O => \N__37946\,
            I => \N__37940\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__37943\,
            I => \N__37935\
        );

    \I__5987\ : InMux
    port map (
            O => \N__37940\,
            I => \N__37932\
        );

    \I__5986\ : InMux
    port map (
            O => \N__37939\,
            I => \N__37927\
        );

    \I__5985\ : InMux
    port map (
            O => \N__37938\,
            I => \N__37927\
        );

    \I__5984\ : Span4Mux_h
    port map (
            O => \N__37935\,
            I => \N__37923\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__37932\,
            I => \N__37920\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__37927\,
            I => \N__37917\
        );

    \I__5981\ : InMux
    port map (
            O => \N__37926\,
            I => \N__37914\
        );

    \I__5980\ : Span4Mux_h
    port map (
            O => \N__37923\,
            I => \N__37911\
        );

    \I__5979\ : Span4Mux_h
    port map (
            O => \N__37920\,
            I => \N__37906\
        );

    \I__5978\ : Span4Mux_h
    port map (
            O => \N__37917\,
            I => \N__37906\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__37914\,
            I => encoder1_position_24
        );

    \I__5976\ : Odrv4
    port map (
            O => \N__37911\,
            I => encoder1_position_24
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__37906\,
            I => encoder1_position_24
        );

    \I__5974\ : InMux
    port map (
            O => \N__37899\,
            I => \N__37896\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__37896\,
            I => \N__37893\
        );

    \I__5972\ : Span4Mux_h
    port map (
            O => \N__37893\,
            I => \N__37890\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__37890\,
            I => \N__37887\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__37887\,
            I => \c0.n10_adj_4367\
        );

    \I__5969\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37881\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__37881\,
            I => \c0.n10_adj_4239\
        );

    \I__5967\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37875\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__37875\,
            I => \c0.n13049\
        );

    \I__5965\ : InMux
    port map (
            O => \N__37872\,
            I => \N__37869\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__37869\,
            I => \N__37866\
        );

    \I__5963\ : Span4Mux_v
    port map (
            O => \N__37866\,
            I => \N__37862\
        );

    \I__5962\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37857\
        );

    \I__5961\ : Span4Mux_h
    port map (
            O => \N__37862\,
            I => \N__37854\
        );

    \I__5960\ : InMux
    port map (
            O => \N__37861\,
            I => \N__37851\
        );

    \I__5959\ : InMux
    port map (
            O => \N__37860\,
            I => \N__37848\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__37857\,
            I => data_in_2_4
        );

    \I__5957\ : Odrv4
    port map (
            O => \N__37854\,
            I => data_in_2_4
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__37851\,
            I => data_in_2_4
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__37848\,
            I => data_in_2_4
        );

    \I__5954\ : CascadeMux
    port map (
            O => \N__37839\,
            I => \c0.n13049_cascade_\
        );

    \I__5953\ : CascadeMux
    port map (
            O => \N__37836\,
            I => \c0.n18_adj_4236_cascade_\
        );

    \I__5952\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37830\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__37830\,
            I => \c0.n20_adj_4237\
        );

    \I__5950\ : CascadeMux
    port map (
            O => \N__37827\,
            I => \N__37823\
        );

    \I__5949\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37819\
        );

    \I__5948\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37816\
        );

    \I__5947\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37813\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__37819\,
            I => \N__37809\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__37816\,
            I => \N__37804\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__37813\,
            I => \N__37804\
        );

    \I__5943\ : InMux
    port map (
            O => \N__37812\,
            I => \N__37801\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__37809\,
            I => \N__37796\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__37804\,
            I => \N__37796\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__37801\,
            I => data_in_1_4
        );

    \I__5939\ : Odrv4
    port map (
            O => \N__37796\,
            I => data_in_1_4
        );

    \I__5938\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37788\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__37788\,
            I => \c0.n14_adj_4241\
        );

    \I__5936\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37782\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__37782\,
            I => \c0.n22489\
        );

    \I__5934\ : InMux
    port map (
            O => \N__37779\,
            I => \N__37775\
        );

    \I__5933\ : InMux
    port map (
            O => \N__37778\,
            I => \N__37772\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__37775\,
            I => \N__37769\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__37772\,
            I => \N__37766\
        );

    \I__5930\ : Odrv4
    port map (
            O => \N__37769\,
            I => \c0.n21393\
        );

    \I__5929\ : Odrv4
    port map (
            O => \N__37766\,
            I => \c0.n21393\
        );

    \I__5928\ : CascadeMux
    port map (
            O => \N__37761\,
            I => \N__37758\
        );

    \I__5927\ : InMux
    port map (
            O => \N__37758\,
            I => \N__37755\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__37755\,
            I => \c0.n22797\
        );

    \I__5925\ : InMux
    port map (
            O => \N__37752\,
            I => \N__37749\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__37749\,
            I => \N__37746\
        );

    \I__5923\ : Odrv12
    port map (
            O => \N__37746\,
            I => \c0.n26_adj_4697\
        );

    \I__5922\ : InMux
    port map (
            O => \N__37743\,
            I => \N__37739\
        );

    \I__5921\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37736\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__37739\,
            I => \N__37733\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__37736\,
            I => \N__37730\
        );

    \I__5918\ : Odrv12
    port map (
            O => \N__37733\,
            I => \c0.n22475\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__37730\,
            I => \c0.n22475\
        );

    \I__5916\ : InMux
    port map (
            O => \N__37725\,
            I => \N__37722\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__37722\,
            I => \N__37718\
        );

    \I__5914\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37715\
        );

    \I__5913\ : Odrv12
    port map (
            O => \N__37718\,
            I => \c0.data_out_frame_29__7__N_1143\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__37715\,
            I => \c0.data_out_frame_29__7__N_1143\
        );

    \I__5911\ : InMux
    port map (
            O => \N__37710\,
            I => \N__37707\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__37707\,
            I => \N__37704\
        );

    \I__5909\ : Span4Mux_h
    port map (
            O => \N__37704\,
            I => \N__37701\
        );

    \I__5908\ : Odrv4
    port map (
            O => \N__37701\,
            I => \c0.n10_adj_4214\
        );

    \I__5907\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37695\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__37695\,
            I => \N__37692\
        );

    \I__5905\ : Span4Mux_h
    port map (
            O => \N__37692\,
            I => \N__37689\
        );

    \I__5904\ : Span4Mux_h
    port map (
            O => \N__37689\,
            I => \N__37686\
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__37686\,
            I => \c0.data_out_frame_28_1\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__37683\,
            I => \N__37680\
        );

    \I__5901\ : InMux
    port map (
            O => \N__37680\,
            I => \N__37677\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__37677\,
            I => \N__37674\
        );

    \I__5899\ : Odrv12
    port map (
            O => \N__37674\,
            I => \c0.n24033\
        );

    \I__5898\ : InMux
    port map (
            O => \N__37671\,
            I => \N__37668\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__37668\,
            I => \c0.n27_adj_4696\
        );

    \I__5896\ : InMux
    port map (
            O => \N__37665\,
            I => \N__37661\
        );

    \I__5895\ : InMux
    port map (
            O => \N__37664\,
            I => \N__37658\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__37661\,
            I => data_in_0_0
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__37658\,
            I => data_in_0_0
        );

    \I__5892\ : CascadeMux
    port map (
            O => \N__37653\,
            I => \N__37649\
        );

    \I__5891\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37644\
        );

    \I__5890\ : InMux
    port map (
            O => \N__37649\,
            I => \N__37644\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__37644\,
            I => data_in_0_4
        );

    \I__5888\ : CascadeMux
    port map (
            O => \N__37641\,
            I => \c0.n15_adj_4242_cascade_\
        );

    \I__5887\ : InMux
    port map (
            O => \N__37638\,
            I => \N__37634\
        );

    \I__5886\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37631\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__37634\,
            I => \c0.n20766\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__37631\,
            I => \c0.n20766\
        );

    \I__5883\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37623\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__37623\,
            I => \N__37620\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__37620\,
            I => n2335
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__37617\,
            I => \N__37614\
        );

    \I__5879\ : InMux
    port map (
            O => \N__37614\,
            I => \N__37611\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__37611\,
            I => \c0.n10427\
        );

    \I__5877\ : CascadeMux
    port map (
            O => \N__37608\,
            I => \c0.n21360_cascade_\
        );

    \I__5876\ : InMux
    port map (
            O => \N__37605\,
            I => \N__37602\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__37602\,
            I => \N__37598\
        );

    \I__5874\ : InMux
    port map (
            O => \N__37601\,
            I => \N__37594\
        );

    \I__5873\ : Span4Mux_h
    port map (
            O => \N__37598\,
            I => \N__37591\
        );

    \I__5872\ : InMux
    port map (
            O => \N__37597\,
            I => \N__37588\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__37594\,
            I => \c0.n10504\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__37591\,
            I => \c0.n10504\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__37588\,
            I => \c0.n10504\
        );

    \I__5868\ : InMux
    port map (
            O => \N__37581\,
            I => \N__37578\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__37578\,
            I => \N__37574\
        );

    \I__5866\ : InMux
    port map (
            O => \N__37577\,
            I => \N__37571\
        );

    \I__5865\ : Span4Mux_h
    port map (
            O => \N__37574\,
            I => \N__37568\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__37571\,
            I => \N__37565\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__37568\,
            I => \c0.n22366\
        );

    \I__5862\ : Odrv12
    port map (
            O => \N__37565\,
            I => \c0.n22366\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__37560\,
            I => \c0.n10504_cascade_\
        );

    \I__5860\ : InMux
    port map (
            O => \N__37557\,
            I => \N__37551\
        );

    \I__5859\ : InMux
    port map (
            O => \N__37556\,
            I => \N__37551\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__37551\,
            I => \N__37548\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__37548\,
            I => \c0.n22327\
        );

    \I__5856\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37542\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__37542\,
            I => \N__37539\
        );

    \I__5854\ : Span4Mux_v
    port map (
            O => \N__37539\,
            I => \N__37536\
        );

    \I__5853\ : Span4Mux_h
    port map (
            O => \N__37536\,
            I => \N__37532\
        );

    \I__5852\ : InMux
    port map (
            O => \N__37535\,
            I => \N__37529\
        );

    \I__5851\ : Sp12to4
    port map (
            O => \N__37532\,
            I => \N__37524\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__37529\,
            I => \N__37524\
        );

    \I__5849\ : Odrv12
    port map (
            O => \N__37524\,
            I => n21484
        );

    \I__5848\ : InMux
    port map (
            O => \N__37521\,
            I => \N__37518\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__37518\,
            I => \N__37515\
        );

    \I__5846\ : Span4Mux_h
    port map (
            O => \N__37515\,
            I => \N__37512\
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__37512\,
            I => \c0.n28_adj_4698\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__37509\,
            I => \c0.n25_adj_4695_cascade_\
        );

    \I__5843\ : CascadeMux
    port map (
            O => \N__37506\,
            I => \N__37503\
        );

    \I__5842\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37500\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__37500\,
            I => \N__37497\
        );

    \I__5840\ : Span12Mux_v
    port map (
            O => \N__37497\,
            I => \N__37494\
        );

    \I__5839\ : Odrv12
    port map (
            O => \N__37494\,
            I => \c0.data_out_frame_29_1\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__37491\,
            I => \N__37480\
        );

    \I__5837\ : CascadeMux
    port map (
            O => \N__37490\,
            I => \N__37475\
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__37489\,
            I => \N__37471\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__37488\,
            I => \N__37467\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__37487\,
            I => \N__37463\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__37486\,
            I => \N__37459\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__37485\,
            I => \N__37455\
        );

    \I__5831\ : CascadeMux
    port map (
            O => \N__37484\,
            I => \N__37451\
        );

    \I__5830\ : InMux
    port map (
            O => \N__37483\,
            I => \N__37441\
        );

    \I__5829\ : InMux
    port map (
            O => \N__37480\,
            I => \N__37436\
        );

    \I__5828\ : InMux
    port map (
            O => \N__37479\,
            I => \N__37436\
        );

    \I__5827\ : InMux
    port map (
            O => \N__37478\,
            I => \N__37423\
        );

    \I__5826\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37423\
        );

    \I__5825\ : InMux
    port map (
            O => \N__37474\,
            I => \N__37423\
        );

    \I__5824\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37423\
        );

    \I__5823\ : InMux
    port map (
            O => \N__37470\,
            I => \N__37423\
        );

    \I__5822\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37423\
        );

    \I__5821\ : InMux
    port map (
            O => \N__37466\,
            I => \N__37406\
        );

    \I__5820\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37406\
        );

    \I__5819\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37406\
        );

    \I__5818\ : InMux
    port map (
            O => \N__37459\,
            I => \N__37406\
        );

    \I__5817\ : InMux
    port map (
            O => \N__37458\,
            I => \N__37406\
        );

    \I__5816\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37406\
        );

    \I__5815\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37406\
        );

    \I__5814\ : InMux
    port map (
            O => \N__37451\,
            I => \N__37406\
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__37450\,
            I => \N__37403\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__37449\,
            I => \N__37400\
        );

    \I__5811\ : CascadeMux
    port map (
            O => \N__37448\,
            I => \N__37397\
        );

    \I__5810\ : CascadeMux
    port map (
            O => \N__37447\,
            I => \N__37394\
        );

    \I__5809\ : CascadeMux
    port map (
            O => \N__37446\,
            I => \N__37391\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__37445\,
            I => \N__37388\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__37444\,
            I => \N__37385\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__37441\,
            I => \N__37371\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__37436\,
            I => \N__37371\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__37423\,
            I => \N__37371\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__37406\,
            I => \N__37371\
        );

    \I__5802\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37362\
        );

    \I__5801\ : InMux
    port map (
            O => \N__37400\,
            I => \N__37362\
        );

    \I__5800\ : InMux
    port map (
            O => \N__37397\,
            I => \N__37362\
        );

    \I__5799\ : InMux
    port map (
            O => \N__37394\,
            I => \N__37362\
        );

    \I__5798\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37353\
        );

    \I__5797\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37353\
        );

    \I__5796\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37353\
        );

    \I__5795\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37353\
        );

    \I__5794\ : CascadeMux
    port map (
            O => \N__37383\,
            I => \N__37350\
        );

    \I__5793\ : CascadeMux
    port map (
            O => \N__37382\,
            I => \N__37346\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__37381\,
            I => \N__37342\
        );

    \I__5791\ : CascadeMux
    port map (
            O => \N__37380\,
            I => \N__37338\
        );

    \I__5790\ : Span4Mux_v
    port map (
            O => \N__37371\,
            I => \N__37334\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__37362\,
            I => \N__37331\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__37353\,
            I => \N__37328\
        );

    \I__5787\ : InMux
    port map (
            O => \N__37350\,
            I => \N__37311\
        );

    \I__5786\ : InMux
    port map (
            O => \N__37349\,
            I => \N__37311\
        );

    \I__5785\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37311\
        );

    \I__5784\ : InMux
    port map (
            O => \N__37345\,
            I => \N__37311\
        );

    \I__5783\ : InMux
    port map (
            O => \N__37342\,
            I => \N__37311\
        );

    \I__5782\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37311\
        );

    \I__5781\ : InMux
    port map (
            O => \N__37338\,
            I => \N__37311\
        );

    \I__5780\ : InMux
    port map (
            O => \N__37337\,
            I => \N__37311\
        );

    \I__5779\ : Span4Mux_h
    port map (
            O => \N__37334\,
            I => \N__37304\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__37331\,
            I => \N__37304\
        );

    \I__5777\ : Span4Mux_h
    port map (
            O => \N__37328\,
            I => \N__37304\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__37311\,
            I => \N__37301\
        );

    \I__5775\ : Span4Mux_h
    port map (
            O => \N__37304\,
            I => \N__37298\
        );

    \I__5774\ : Odrv12
    port map (
            O => \N__37301\,
            I => \quad_counter0.n2313\
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__37298\,
            I => \quad_counter0.n2313\
        );

    \I__5772\ : InMux
    port map (
            O => \N__37293\,
            I => \bfn_14_13_0_\
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__37290\,
            I => \n2326_cascade_\
        );

    \I__5770\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37284\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__37284\,
            I => \N__37280\
        );

    \I__5768\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37277\
        );

    \I__5767\ : Span12Mux_s10_h
    port map (
            O => \N__37280\,
            I => \N__37272\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__37277\,
            I => \N__37272\
        );

    \I__5765\ : Span12Mux_h
    port map (
            O => \N__37272\,
            I => \N__37269\
        );

    \I__5764\ : Odrv12
    port map (
            O => \N__37269\,
            I => \c0.n22218\
        );

    \I__5763\ : CascadeMux
    port map (
            O => \N__37266\,
            I => \N__37262\
        );

    \I__5762\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37259\
        );

    \I__5761\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37255\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__37259\,
            I => \N__37252\
        );

    \I__5759\ : InMux
    port map (
            O => \N__37258\,
            I => \N__37249\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__37255\,
            I => \N__37246\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__37252\,
            I => \N__37243\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__37249\,
            I => \N__37240\
        );

    \I__5755\ : Span4Mux_v
    port map (
            O => \N__37246\,
            I => \N__37235\
        );

    \I__5754\ : Span4Mux_h
    port map (
            O => \N__37243\,
            I => \N__37235\
        );

    \I__5753\ : Span4Mux_v
    port map (
            O => \N__37240\,
            I => \N__37232\
        );

    \I__5752\ : Odrv4
    port map (
            O => \N__37235\,
            I => \c0.n21323\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__37232\,
            I => \c0.n21323\
        );

    \I__5750\ : InMux
    port map (
            O => \N__37227\,
            I => \N__37224\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__37224\,
            I => \N__37221\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__37221\,
            I => \c0.n22671\
        );

    \I__5747\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37215\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__37215\,
            I => \N__37212\
        );

    \I__5745\ : Odrv12
    port map (
            O => \N__37212\,
            I => \c0.n20_adj_4694\
        );

    \I__5744\ : InMux
    port map (
            O => \N__37209\,
            I => \N__37205\
        );

    \I__5743\ : InMux
    port map (
            O => \N__37208\,
            I => \N__37202\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__37205\,
            I => \N__37198\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__37202\,
            I => \N__37195\
        );

    \I__5740\ : InMux
    port map (
            O => \N__37201\,
            I => \N__37192\
        );

    \I__5739\ : Span4Mux_h
    port map (
            O => \N__37198\,
            I => \N__37189\
        );

    \I__5738\ : Span4Mux_h
    port map (
            O => \N__37195\,
            I => \N__37183\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__37192\,
            I => \N__37183\
        );

    \I__5736\ : Span4Mux_v
    port map (
            O => \N__37189\,
            I => \N__37180\
        );

    \I__5735\ : InMux
    port map (
            O => \N__37188\,
            I => \N__37177\
        );

    \I__5734\ : Odrv4
    port map (
            O => \N__37183\,
            I => \c0.n20348\
        );

    \I__5733\ : Odrv4
    port map (
            O => \N__37180\,
            I => \c0.n20348\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__37177\,
            I => \c0.n20348\
        );

    \I__5731\ : CascadeMux
    port map (
            O => \N__37170\,
            I => \N__37165\
        );

    \I__5730\ : InMux
    port map (
            O => \N__37169\,
            I => \N__37161\
        );

    \I__5729\ : InMux
    port map (
            O => \N__37168\,
            I => \N__37158\
        );

    \I__5728\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37153\
        );

    \I__5727\ : InMux
    port map (
            O => \N__37164\,
            I => \N__37153\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__37161\,
            I => \c0.n21330\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__37158\,
            I => \c0.n21330\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__37153\,
            I => \c0.n21330\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__37146\,
            I => \c0.n21355_cascade_\
        );

    \I__5722\ : InMux
    port map (
            O => \N__37143\,
            I => \N__37140\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__37140\,
            I => \N__37134\
        );

    \I__5720\ : InMux
    port map (
            O => \N__37139\,
            I => \N__37131\
        );

    \I__5719\ : CascadeMux
    port map (
            O => \N__37138\,
            I => \N__37128\
        );

    \I__5718\ : InMux
    port map (
            O => \N__37137\,
            I => \N__37125\
        );

    \I__5717\ : Span4Mux_v
    port map (
            O => \N__37134\,
            I => \N__37120\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__37131\,
            I => \N__37120\
        );

    \I__5715\ : InMux
    port map (
            O => \N__37128\,
            I => \N__37117\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__37125\,
            I => \N__37112\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__37120\,
            I => \N__37107\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__37117\,
            I => \N__37107\
        );

    \I__5711\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37104\
        );

    \I__5710\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37101\
        );

    \I__5709\ : Odrv4
    port map (
            O => \N__37112\,
            I => \c0.n12464\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__37107\,
            I => \c0.n12464\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__37104\,
            I => \c0.n12464\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__37101\,
            I => \c0.n12464\
        );

    \I__5705\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37088\
        );

    \I__5704\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37085\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__37088\,
            I => \c0.n20404\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__37085\,
            I => \c0.n20404\
        );

    \I__5701\ : InMux
    port map (
            O => \N__37080\,
            I => \quad_counter0.n19785\
        );

    \I__5700\ : InMux
    port map (
            O => \N__37077\,
            I => \bfn_14_12_0_\
        );

    \I__5699\ : InMux
    port map (
            O => \N__37074\,
            I => \N__37071\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__37071\,
            I => n2333
        );

    \I__5697\ : InMux
    port map (
            O => \N__37068\,
            I => \quad_counter0.n19787\
        );

    \I__5696\ : InMux
    port map (
            O => \N__37065\,
            I => \N__37062\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__37062\,
            I => n2332
        );

    \I__5694\ : InMux
    port map (
            O => \N__37059\,
            I => \quad_counter0.n19788\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__37056\,
            I => \N__37053\
        );

    \I__5692\ : InMux
    port map (
            O => \N__37053\,
            I => \N__37049\
        );

    \I__5691\ : InMux
    port map (
            O => \N__37052\,
            I => \N__37046\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__37049\,
            I => \N__37042\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__37046\,
            I => \N__37039\
        );

    \I__5688\ : CascadeMux
    port map (
            O => \N__37045\,
            I => \N__37036\
        );

    \I__5687\ : Span12Mux_v
    port map (
            O => \N__37042\,
            I => \N__37030\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__37039\,
            I => \N__37027\
        );

    \I__5685\ : InMux
    port map (
            O => \N__37036\,
            I => \N__37022\
        );

    \I__5684\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37022\
        );

    \I__5683\ : InMux
    port map (
            O => \N__37034\,
            I => \N__37017\
        );

    \I__5682\ : InMux
    port map (
            O => \N__37033\,
            I => \N__37017\
        );

    \I__5681\ : Odrv12
    port map (
            O => \N__37030\,
            I => encoder0_position_26
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__37027\,
            I => encoder0_position_26
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__37022\,
            I => encoder0_position_26
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__37017\,
            I => encoder0_position_26
        );

    \I__5677\ : InMux
    port map (
            O => \N__37008\,
            I => \N__37005\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__37005\,
            I => \N__37002\
        );

    \I__5675\ : Span4Mux_v
    port map (
            O => \N__37002\,
            I => \N__36999\
        );

    \I__5674\ : Odrv4
    port map (
            O => \N__36999\,
            I => n2331
        );

    \I__5673\ : InMux
    port map (
            O => \N__36996\,
            I => \quad_counter0.n19789\
        );

    \I__5672\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36990\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__36990\,
            I => n2330
        );

    \I__5670\ : InMux
    port map (
            O => \N__36987\,
            I => \quad_counter0.n19790\
        );

    \I__5669\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36981\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__36981\,
            I => \N__36978\
        );

    \I__5667\ : Span4Mux_v
    port map (
            O => \N__36978\,
            I => \N__36971\
        );

    \I__5666\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36968\
        );

    \I__5665\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36965\
        );

    \I__5664\ : CascadeMux
    port map (
            O => \N__36975\,
            I => \N__36961\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__36974\,
            I => \N__36958\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__36971\,
            I => \N__36952\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__36968\,
            I => \N__36952\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__36965\,
            I => \N__36948\
        );

    \I__5659\ : InMux
    port map (
            O => \N__36964\,
            I => \N__36945\
        );

    \I__5658\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36940\
        );

    \I__5657\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36940\
        );

    \I__5656\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36937\
        );

    \I__5655\ : Span4Mux_v
    port map (
            O => \N__36952\,
            I => \N__36934\
        );

    \I__5654\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36931\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__36948\,
            I => \N__36928\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__36945\,
            I => \N__36923\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__36940\,
            I => \N__36923\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__36937\,
            I => encoder0_position_28
        );

    \I__5649\ : Odrv4
    port map (
            O => \N__36934\,
            I => encoder0_position_28
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__36931\,
            I => encoder0_position_28
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__36928\,
            I => encoder0_position_28
        );

    \I__5646\ : Odrv4
    port map (
            O => \N__36923\,
            I => encoder0_position_28
        );

    \I__5645\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36909\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__36909\,
            I => \N__36906\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__36906\,
            I => \N__36903\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__36903\,
            I => n2329
        );

    \I__5641\ : InMux
    port map (
            O => \N__36900\,
            I => \quad_counter0.n19791\
        );

    \I__5640\ : InMux
    port map (
            O => \N__36897\,
            I => \N__36894\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__36894\,
            I => \N__36890\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__36893\,
            I => \N__36887\
        );

    \I__5637\ : Span4Mux_v
    port map (
            O => \N__36890\,
            I => \N__36884\
        );

    \I__5636\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36881\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__36884\,
            I => \N__36878\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__36881\,
            I => \N__36875\
        );

    \I__5633\ : Span4Mux_v
    port map (
            O => \N__36878\,
            I => \N__36867\
        );

    \I__5632\ : Span4Mux_h
    port map (
            O => \N__36875\,
            I => \N__36864\
        );

    \I__5631\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36857\
        );

    \I__5630\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36857\
        );

    \I__5629\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36857\
        );

    \I__5628\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36852\
        );

    \I__5627\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36852\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__36867\,
            I => encoder0_position_29
        );

    \I__5625\ : Odrv4
    port map (
            O => \N__36864\,
            I => encoder0_position_29
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__36857\,
            I => encoder0_position_29
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__36852\,
            I => encoder0_position_29
        );

    \I__5622\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36840\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__36840\,
            I => \N__36837\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__36837\,
            I => \N__36834\
        );

    \I__5619\ : Span4Mux_h
    port map (
            O => \N__36834\,
            I => \N__36831\
        );

    \I__5618\ : Odrv4
    port map (
            O => \N__36831\,
            I => n2328
        );

    \I__5617\ : InMux
    port map (
            O => \N__36828\,
            I => \quad_counter0.n19792\
        );

    \I__5616\ : InMux
    port map (
            O => \N__36825\,
            I => \N__36822\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__36822\,
            I => \N__36819\
        );

    \I__5614\ : Odrv12
    port map (
            O => \N__36819\,
            I => n2327
        );

    \I__5613\ : InMux
    port map (
            O => \N__36816\,
            I => \quad_counter0.n19793\
        );

    \I__5612\ : InMux
    port map (
            O => \N__36813\,
            I => \quad_counter0.n19776\
        );

    \I__5611\ : InMux
    port map (
            O => \N__36810\,
            I => \quad_counter0.n19777\
        );

    \I__5610\ : InMux
    port map (
            O => \N__36807\,
            I => \bfn_14_11_0_\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__36804\,
            I => \N__36798\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__36803\,
            I => \N__36795\
        );

    \I__5607\ : InMux
    port map (
            O => \N__36802\,
            I => \N__36792\
        );

    \I__5606\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36789\
        );

    \I__5605\ : InMux
    port map (
            O => \N__36798\,
            I => \N__36785\
        );

    \I__5604\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36781\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__36792\,
            I => \N__36776\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__36789\,
            I => \N__36776\
        );

    \I__5601\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36773\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__36785\,
            I => \N__36770\
        );

    \I__5599\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36767\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__36781\,
            I => \N__36760\
        );

    \I__5597\ : Span4Mux_v
    port map (
            O => \N__36776\,
            I => \N__36760\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__36773\,
            I => \N__36760\
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__36770\,
            I => encoder0_position_16
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__36767\,
            I => encoder0_position_16
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__36760\,
            I => encoder0_position_16
        );

    \I__5592\ : InMux
    port map (
            O => \N__36753\,
            I => \N__36750\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36747\
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__36747\,
            I => n2341
        );

    \I__5589\ : InMux
    port map (
            O => \N__36744\,
            I => \quad_counter0.n19779\
        );

    \I__5588\ : InMux
    port map (
            O => \N__36741\,
            I => \quad_counter0.n19780\
        );

    \I__5587\ : InMux
    port map (
            O => \N__36738\,
            I => \quad_counter0.n19781\
        );

    \I__5586\ : InMux
    port map (
            O => \N__36735\,
            I => \quad_counter0.n19782\
        );

    \I__5585\ : InMux
    port map (
            O => \N__36732\,
            I => \quad_counter0.n19783\
        );

    \I__5584\ : InMux
    port map (
            O => \N__36729\,
            I => \quad_counter0.n19784\
        );

    \I__5583\ : InMux
    port map (
            O => \N__36726\,
            I => \quad_counter0.n19768\
        );

    \I__5582\ : InMux
    port map (
            O => \N__36723\,
            I => \N__36720\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__36720\,
            I => \N__36717\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__36717\,
            I => n2351
        );

    \I__5579\ : InMux
    port map (
            O => \N__36714\,
            I => \quad_counter0.n19769\
        );

    \I__5578\ : CascadeMux
    port map (
            O => \N__36711\,
            I => \N__36708\
        );

    \I__5577\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36703\
        );

    \I__5576\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36698\
        );

    \I__5575\ : InMux
    port map (
            O => \N__36706\,
            I => \N__36698\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__36703\,
            I => \N__36694\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__36698\,
            I => \N__36690\
        );

    \I__5572\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36685\
        );

    \I__5571\ : Span12Mux_v
    port map (
            O => \N__36694\,
            I => \N__36682\
        );

    \I__5570\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36679\
        );

    \I__5569\ : Span4Mux_v
    port map (
            O => \N__36690\,
            I => \N__36676\
        );

    \I__5568\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36673\
        );

    \I__5567\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36670\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__36685\,
            I => \N__36667\
        );

    \I__5565\ : Span12Mux_v
    port map (
            O => \N__36682\,
            I => \N__36664\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__36679\,
            I => \N__36659\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__36676\,
            I => \N__36659\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__36673\,
            I => \N__36652\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__36670\,
            I => \N__36652\
        );

    \I__5560\ : Span4Mux_v
    port map (
            O => \N__36667\,
            I => \N__36652\
        );

    \I__5559\ : Odrv12
    port map (
            O => \N__36664\,
            I => encoder0_position_7
        );

    \I__5558\ : Odrv4
    port map (
            O => \N__36659\,
            I => encoder0_position_7
        );

    \I__5557\ : Odrv4
    port map (
            O => \N__36652\,
            I => encoder0_position_7
        );

    \I__5556\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36642\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__36642\,
            I => \N__36639\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__36639\,
            I => n2350
        );

    \I__5553\ : InMux
    port map (
            O => \N__36636\,
            I => \bfn_14_10_0_\
        );

    \I__5552\ : InMux
    port map (
            O => \N__36633\,
            I => \quad_counter0.n19771\
        );

    \I__5551\ : InMux
    port map (
            O => \N__36630\,
            I => \quad_counter0.n19772\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__36627\,
            I => \N__36624\
        );

    \I__5549\ : InMux
    port map (
            O => \N__36624\,
            I => \N__36619\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__36623\,
            I => \N__36616\
        );

    \I__5547\ : CascadeMux
    port map (
            O => \N__36622\,
            I => \N__36613\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__36619\,
            I => \N__36610\
        );

    \I__5545\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36607\
        );

    \I__5544\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36604\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__36610\,
            I => \N__36599\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__36607\,
            I => \N__36599\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__36604\,
            I => \N__36594\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__36599\,
            I => \N__36591\
        );

    \I__5539\ : InMux
    port map (
            O => \N__36598\,
            I => \N__36586\
        );

    \I__5538\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36586\
        );

    \I__5537\ : Odrv12
    port map (
            O => \N__36594\,
            I => encoder0_position_10
        );

    \I__5536\ : Odrv4
    port map (
            O => \N__36591\,
            I => encoder0_position_10
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__36586\,
            I => encoder0_position_10
        );

    \I__5534\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36576\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__36576\,
            I => \N__36573\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__36573\,
            I => \N__36570\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__36570\,
            I => n2347
        );

    \I__5530\ : InMux
    port map (
            O => \N__36567\,
            I => \quad_counter0.n19773\
        );

    \I__5529\ : CascadeMux
    port map (
            O => \N__36564\,
            I => \N__36561\
        );

    \I__5528\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36558\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__36558\,
            I => \N__36555\
        );

    \I__5526\ : Span4Mux_h
    port map (
            O => \N__36555\,
            I => \N__36551\
        );

    \I__5525\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36548\
        );

    \I__5524\ : Span4Mux_v
    port map (
            O => \N__36551\,
            I => \N__36544\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__36548\,
            I => \N__36541\
        );

    \I__5522\ : InMux
    port map (
            O => \N__36547\,
            I => \N__36537\
        );

    \I__5521\ : Span4Mux_h
    port map (
            O => \N__36544\,
            I => \N__36532\
        );

    \I__5520\ : Span4Mux_h
    port map (
            O => \N__36541\,
            I => \N__36532\
        );

    \I__5519\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36529\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__36537\,
            I => encoder0_position_11
        );

    \I__5517\ : Odrv4
    port map (
            O => \N__36532\,
            I => encoder0_position_11
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__36529\,
            I => encoder0_position_11
        );

    \I__5515\ : InMux
    port map (
            O => \N__36522\,
            I => \N__36519\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__36519\,
            I => \N__36516\
        );

    \I__5513\ : Span4Mux_v
    port map (
            O => \N__36516\,
            I => \N__36513\
        );

    \I__5512\ : Sp12to4
    port map (
            O => \N__36513\,
            I => \N__36510\
        );

    \I__5511\ : Odrv12
    port map (
            O => \N__36510\,
            I => n2346
        );

    \I__5510\ : InMux
    port map (
            O => \N__36507\,
            I => \quad_counter0.n19774\
        );

    \I__5509\ : CascadeMux
    port map (
            O => \N__36504\,
            I => \N__36501\
        );

    \I__5508\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36497\
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__36500\,
            I => \N__36494\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__36497\,
            I => \N__36491\
        );

    \I__5505\ : InMux
    port map (
            O => \N__36494\,
            I => \N__36484\
        );

    \I__5504\ : Span4Mux_h
    port map (
            O => \N__36491\,
            I => \N__36481\
        );

    \I__5503\ : InMux
    port map (
            O => \N__36490\,
            I => \N__36476\
        );

    \I__5502\ : InMux
    port map (
            O => \N__36489\,
            I => \N__36476\
        );

    \I__5501\ : InMux
    port map (
            O => \N__36488\,
            I => \N__36473\
        );

    \I__5500\ : InMux
    port map (
            O => \N__36487\,
            I => \N__36470\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__36484\,
            I => \N__36467\
        );

    \I__5498\ : Sp12to4
    port map (
            O => \N__36481\,
            I => \N__36460\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__36476\,
            I => \N__36460\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__36473\,
            I => \N__36460\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__36470\,
            I => encoder0_position_12
        );

    \I__5494\ : Odrv12
    port map (
            O => \N__36467\,
            I => encoder0_position_12
        );

    \I__5493\ : Odrv12
    port map (
            O => \N__36460\,
            I => encoder0_position_12
        );

    \I__5492\ : InMux
    port map (
            O => \N__36453\,
            I => \N__36450\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__36450\,
            I => \N__36447\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__36447\,
            I => \N__36444\
        );

    \I__5489\ : Span4Mux_v
    port map (
            O => \N__36444\,
            I => \N__36441\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__36441\,
            I => \N__36438\
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__36438\,
            I => n2345
        );

    \I__5486\ : InMux
    port map (
            O => \N__36435\,
            I => \quad_counter0.n19775\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__36432\,
            I => \N__36429\
        );

    \I__5484\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36426\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__36426\,
            I => \N__36423\
        );

    \I__5482\ : Span4Mux_h
    port map (
            O => \N__36423\,
            I => \N__36418\
        );

    \I__5481\ : InMux
    port map (
            O => \N__36422\,
            I => \N__36415\
        );

    \I__5480\ : InMux
    port map (
            O => \N__36421\,
            I => \N__36410\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__36418\,
            I => \N__36405\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__36415\,
            I => \N__36405\
        );

    \I__5477\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36402\
        );

    \I__5476\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36399\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__36410\,
            I => \N__36394\
        );

    \I__5474\ : Span4Mux_v
    port map (
            O => \N__36405\,
            I => \N__36394\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__36402\,
            I => encoder0_position_0
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__36399\,
            I => encoder0_position_0
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__36394\,
            I => encoder0_position_0
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__36387\,
            I => \N__36384\
        );

    \I__5469\ : InMux
    port map (
            O => \N__36384\,
            I => \N__36381\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__36381\,
            I => \N__36378\
        );

    \I__5467\ : Span12Mux_s11_v
    port map (
            O => \N__36378\,
            I => \N__36375\
        );

    \I__5466\ : Odrv12
    port map (
            O => \N__36375\,
            I => \quad_counter0.count_direction\
        );

    \I__5465\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36369\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__36369\,
            I => n2357
        );

    \I__5463\ : InMux
    port map (
            O => \N__36366\,
            I => \quad_counter0.n19763\
        );

    \I__5462\ : CascadeMux
    port map (
            O => \N__36363\,
            I => \N__36360\
        );

    \I__5461\ : InMux
    port map (
            O => \N__36360\,
            I => \N__36357\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__36357\,
            I => \N__36353\
        );

    \I__5459\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36350\
        );

    \I__5458\ : Sp12to4
    port map (
            O => \N__36353\,
            I => \N__36346\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__36350\,
            I => \N__36343\
        );

    \I__5456\ : InMux
    port map (
            O => \N__36349\,
            I => \N__36338\
        );

    \I__5455\ : Span12Mux_v
    port map (
            O => \N__36346\,
            I => \N__36335\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__36343\,
            I => \N__36332\
        );

    \I__5453\ : InMux
    port map (
            O => \N__36342\,
            I => \N__36329\
        );

    \I__5452\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36326\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__36338\,
            I => encoder0_position_1
        );

    \I__5450\ : Odrv12
    port map (
            O => \N__36335\,
            I => encoder0_position_1
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__36332\,
            I => encoder0_position_1
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__36329\,
            I => encoder0_position_1
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__36326\,
            I => encoder0_position_1
        );

    \I__5446\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36312\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__36312\,
            I => \N__36309\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__36309\,
            I => \N__36306\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__36306\,
            I => n2356
        );

    \I__5442\ : InMux
    port map (
            O => \N__36303\,
            I => \quad_counter0.n19764\
        );

    \I__5441\ : InMux
    port map (
            O => \N__36300\,
            I => \N__36297\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__36297\,
            I => n2355
        );

    \I__5439\ : InMux
    port map (
            O => \N__36294\,
            I => \quad_counter0.n19765\
        );

    \I__5438\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36288\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__36288\,
            I => n2354
        );

    \I__5436\ : InMux
    port map (
            O => \N__36285\,
            I => \quad_counter0.n19766\
        );

    \I__5435\ : InMux
    port map (
            O => \N__36282\,
            I => \N__36279\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__36279\,
            I => \N__36276\
        );

    \I__5433\ : Span4Mux_h
    port map (
            O => \N__36276\,
            I => \N__36273\
        );

    \I__5432\ : Odrv4
    port map (
            O => \N__36273\,
            I => n2353
        );

    \I__5431\ : InMux
    port map (
            O => \N__36270\,
            I => \quad_counter0.n19767\
        );

    \I__5430\ : InMux
    port map (
            O => \N__36267\,
            I => \N__36260\
        );

    \I__5429\ : InMux
    port map (
            O => \N__36266\,
            I => \N__36260\
        );

    \I__5428\ : InMux
    port map (
            O => \N__36265\,
            I => \N__36256\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__36260\,
            I => \N__36253\
        );

    \I__5426\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36250\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__36256\,
            I => \N__36246\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__36253\,
            I => \N__36241\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__36250\,
            I => \N__36241\
        );

    \I__5422\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36238\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__36246\,
            I => \N__36235\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__36241\,
            I => \N__36232\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__36238\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__36235\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__36232\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__5416\ : SRMux
    port map (
            O => \N__36225\,
            I => \N__36222\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__36222\,
            I => \N__36219\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__36219\,
            I => \N__36216\
        );

    \I__5413\ : Odrv4
    port map (
            O => \N__36216\,
            I => \c0.n21653\
        );

    \I__5412\ : InMux
    port map (
            O => \N__36213\,
            I => \N__36209\
        );

    \I__5411\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36206\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__36209\,
            I => \N__36202\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__36206\,
            I => \N__36199\
        );

    \I__5408\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36196\
        );

    \I__5407\ : Span4Mux_h
    port map (
            O => \N__36202\,
            I => \N__36193\
        );

    \I__5406\ : Span4Mux_h
    port map (
            O => \N__36199\,
            I => \N__36190\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__36196\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__5404\ : Odrv4
    port map (
            O => \N__36193\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__36190\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__5402\ : SRMux
    port map (
            O => \N__36183\,
            I => \N__36180\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__36180\,
            I => \N__36177\
        );

    \I__5400\ : Span4Mux_v
    port map (
            O => \N__36177\,
            I => \N__36174\
        );

    \I__5399\ : Odrv4
    port map (
            O => \N__36174\,
            I => \c0.n21649\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__36171\,
            I => \N__36167\
        );

    \I__5397\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36163\
        );

    \I__5396\ : InMux
    port map (
            O => \N__36167\,
            I => \N__36160\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__36166\,
            I => \N__36156\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__36163\,
            I => \N__36152\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__36160\,
            I => \N__36149\
        );

    \I__5392\ : InMux
    port map (
            O => \N__36159\,
            I => \N__36144\
        );

    \I__5391\ : InMux
    port map (
            O => \N__36156\,
            I => \N__36144\
        );

    \I__5390\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36141\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__36152\,
            I => \N__36138\
        );

    \I__5388\ : Span4Mux_h
    port map (
            O => \N__36149\,
            I => \N__36133\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__36144\,
            I => \N__36133\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__36141\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__5385\ : Odrv4
    port map (
            O => \N__36138\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__5384\ : Odrv4
    port map (
            O => \N__36133\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__5383\ : SRMux
    port map (
            O => \N__36126\,
            I => \N__36123\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__36123\,
            I => \N__36120\
        );

    \I__5381\ : Span4Mux_v
    port map (
            O => \N__36120\,
            I => \N__36117\
        );

    \I__5380\ : Span4Mux_h
    port map (
            O => \N__36117\,
            I => \N__36114\
        );

    \I__5379\ : Odrv4
    port map (
            O => \N__36114\,
            I => \c0.n21595\
        );

    \I__5378\ : SRMux
    port map (
            O => \N__36111\,
            I => \N__36108\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__36108\,
            I => \N__36105\
        );

    \I__5376\ : Span4Mux_v
    port map (
            O => \N__36105\,
            I => \N__36102\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__36102\,
            I => \c0.n21643\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__36099\,
            I => \N__36096\
        );

    \I__5373\ : InMux
    port map (
            O => \N__36096\,
            I => \N__36093\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__36093\,
            I => \N__36090\
        );

    \I__5371\ : Span4Mux_v
    port map (
            O => \N__36090\,
            I => \N__36087\
        );

    \I__5370\ : Sp12to4
    port map (
            O => \N__36087\,
            I => \N__36084\
        );

    \I__5369\ : Odrv12
    port map (
            O => \N__36084\,
            I => \c0.n6_adj_4583\
        );

    \I__5368\ : InMux
    port map (
            O => \N__36081\,
            I => \N__36077\
        );

    \I__5367\ : InMux
    port map (
            O => \N__36080\,
            I => \N__36073\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__36077\,
            I => \N__36070\
        );

    \I__5365\ : InMux
    port map (
            O => \N__36076\,
            I => \N__36067\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__36073\,
            I => \N__36064\
        );

    \I__5363\ : Span4Mux_h
    port map (
            O => \N__36070\,
            I => \N__36061\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__36067\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__36064\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__5360\ : Odrv4
    port map (
            O => \N__36061\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__5359\ : InMux
    port map (
            O => \N__36054\,
            I => \N__36051\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__36051\,
            I => \N__36048\
        );

    \I__5357\ : Span4Mux_v
    port map (
            O => \N__36048\,
            I => \N__36045\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__36045\,
            I => \c0.n14_adj_4520\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__36042\,
            I => \N__36038\
        );

    \I__5354\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36035\
        );

    \I__5353\ : InMux
    port map (
            O => \N__36038\,
            I => \N__36032\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__36035\,
            I => \N__36026\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__36032\,
            I => \N__36026\
        );

    \I__5350\ : InMux
    port map (
            O => \N__36031\,
            I => \N__36023\
        );

    \I__5349\ : Span4Mux_h
    port map (
            O => \N__36026\,
            I => \N__36020\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__36023\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__5347\ : Odrv4
    port map (
            O => \N__36020\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__5346\ : InMux
    port map (
            O => \N__36015\,
            I => \N__36012\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__36012\,
            I => \c0.n9_adj_4522\
        );

    \I__5344\ : InMux
    port map (
            O => \N__36009\,
            I => \N__36006\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__36006\,
            I => \c0.n20_adj_4265\
        );

    \I__5342\ : InMux
    port map (
            O => \N__36003\,
            I => \N__36000\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__36000\,
            I => \N__35996\
        );

    \I__5340\ : InMux
    port map (
            O => \N__35999\,
            I => \N__35993\
        );

    \I__5339\ : Span4Mux_h
    port map (
            O => \N__35996\,
            I => \N__35990\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__35993\,
            I => \c0.n16919\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__35990\,
            I => \c0.n16919\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__35985\,
            I => \c0.n20_adj_4265_cascade_\
        );

    \I__5335\ : InMux
    port map (
            O => \N__35982\,
            I => \N__35979\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__35979\,
            I => \N__35976\
        );

    \I__5333\ : Span4Mux_h
    port map (
            O => \N__35976\,
            I => \N__35972\
        );

    \I__5332\ : InMux
    port map (
            O => \N__35975\,
            I => \N__35969\
        );

    \I__5331\ : Odrv4
    port map (
            O => \N__35972\,
            I => \c0.n22148\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__35969\,
            I => \c0.n22148\
        );

    \I__5329\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35960\
        );

    \I__5328\ : InMux
    port map (
            O => \N__35963\,
            I => \N__35957\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__35960\,
            I => \N__35954\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__35957\,
            I => \N__35950\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__35954\,
            I => \N__35947\
        );

    \I__5324\ : InMux
    port map (
            O => \N__35953\,
            I => \N__35944\
        );

    \I__5323\ : Span4Mux_v
    port map (
            O => \N__35950\,
            I => \N__35940\
        );

    \I__5322\ : Sp12to4
    port map (
            O => \N__35947\,
            I => \N__35937\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__35944\,
            I => \N__35934\
        );

    \I__5320\ : InMux
    port map (
            O => \N__35943\,
            I => \N__35931\
        );

    \I__5319\ : Odrv4
    port map (
            O => \N__35940\,
            I => \c0.n22145\
        );

    \I__5318\ : Odrv12
    port map (
            O => \N__35937\,
            I => \c0.n22145\
        );

    \I__5317\ : Odrv4
    port map (
            O => \N__35934\,
            I => \c0.n22145\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__35931\,
            I => \c0.n22145\
        );

    \I__5315\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35919\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__35919\,
            I => \c0.n6_adj_4264\
        );

    \I__5313\ : InMux
    port map (
            O => \N__35916\,
            I => \N__35912\
        );

    \I__5312\ : CascadeMux
    port map (
            O => \N__35915\,
            I => \N__35909\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__35912\,
            I => \N__35905\
        );

    \I__5310\ : InMux
    port map (
            O => \N__35909\,
            I => \N__35902\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__35908\,
            I => \N__35898\
        );

    \I__5308\ : Span4Mux_v
    port map (
            O => \N__35905\,
            I => \N__35892\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__35902\,
            I => \N__35892\
        );

    \I__5306\ : InMux
    port map (
            O => \N__35901\,
            I => \N__35889\
        );

    \I__5305\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35886\
        );

    \I__5304\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35883\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__35892\,
            I => \N__35880\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__35889\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__35886\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__35883\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__5299\ : Odrv4
    port map (
            O => \N__35880\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__5298\ : CascadeMux
    port map (
            O => \N__35871\,
            I => \N__35868\
        );

    \I__5297\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35865\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__35865\,
            I => \N__35862\
        );

    \I__5295\ : Span4Mux_h
    port map (
            O => \N__35862\,
            I => \N__35859\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__35859\,
            I => \N__35856\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__35856\,
            I => \c0.n14721\
        );

    \I__5292\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35850\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__35850\,
            I => \N__35846\
        );

    \I__5290\ : InMux
    port map (
            O => \N__35849\,
            I => \N__35843\
        );

    \I__5289\ : Span4Mux_h
    port map (
            O => \N__35846\,
            I => \N__35840\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__35843\,
            I => \N__35837\
        );

    \I__5287\ : Sp12to4
    port map (
            O => \N__35840\,
            I => \N__35834\
        );

    \I__5286\ : Span4Mux_h
    port map (
            O => \N__35837\,
            I => \N__35831\
        );

    \I__5285\ : Odrv12
    port map (
            O => \N__35834\,
            I => \c0.n14530\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__35831\,
            I => \c0.n14530\
        );

    \I__5283\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35823\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__35823\,
            I => \N__35820\
        );

    \I__5281\ : Span12Mux_h
    port map (
            O => \N__35820\,
            I => \N__35817\
        );

    \I__5280\ : Odrv12
    port map (
            O => \N__35817\,
            I => \c0.n7_adj_4741\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__35814\,
            I => \N__35810\
        );

    \I__5278\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35805\
        );

    \I__5277\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35805\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__35805\,
            I => \N__35802\
        );

    \I__5275\ : Odrv4
    port map (
            O => \N__35802\,
            I => \c0.n9683\
        );

    \I__5274\ : InMux
    port map (
            O => \N__35799\,
            I => \N__35796\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__35796\,
            I => \N__35793\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__35793\,
            I => \c0.n9587\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__35790\,
            I => \c0.n9683_cascade_\
        );

    \I__5270\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35770\
        );

    \I__5269\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35770\
        );

    \I__5268\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35770\
        );

    \I__5267\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35770\
        );

    \I__5266\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35761\
        );

    \I__5265\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35761\
        );

    \I__5264\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35761\
        );

    \I__5263\ : InMux
    port map (
            O => \N__35780\,
            I => \N__35761\
        );

    \I__5262\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35758\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__35770\,
            I => \N__35751\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__35761\,
            I => \N__35751\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35748\
        );

    \I__5258\ : InMux
    port map (
            O => \N__35757\,
            I => \N__35745\
        );

    \I__5257\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35742\
        );

    \I__5256\ : Span4Mux_v
    port map (
            O => \N__35751\,
            I => \N__35739\
        );

    \I__5255\ : Span4Mux_v
    port map (
            O => \N__35748\,
            I => \N__35736\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__35745\,
            I => \N__35733\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__35742\,
            I => \N__35730\
        );

    \I__5252\ : Odrv4
    port map (
            O => \N__35739\,
            I => \c0.n10\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__35736\,
            I => \c0.n10\
        );

    \I__5250\ : Odrv12
    port map (
            O => \N__35733\,
            I => \c0.n10\
        );

    \I__5249\ : Odrv4
    port map (
            O => \N__35730\,
            I => \c0.n10\
        );

    \I__5248\ : InMux
    port map (
            O => \N__35721\,
            I => \N__35716\
        );

    \I__5247\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35711\
        );

    \I__5246\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35711\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__35716\,
            I => \N__35708\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__35711\,
            I => \N__35705\
        );

    \I__5243\ : Span4Mux_v
    port map (
            O => \N__35708\,
            I => \N__35702\
        );

    \I__5242\ : Span4Mux_h
    port map (
            O => \N__35705\,
            I => \N__35699\
        );

    \I__5241\ : Odrv4
    port map (
            O => \N__35702\,
            I => \c0.data_out_frame_29_7_N_1482_2\
        );

    \I__5240\ : Odrv4
    port map (
            O => \N__35699\,
            I => \c0.data_out_frame_29_7_N_1482_2\
        );

    \I__5239\ : CascadeMux
    port map (
            O => \N__35694\,
            I => \c0.n14_adj_4727_cascade_\
        );

    \I__5238\ : CascadeMux
    port map (
            O => \N__35691\,
            I => \N__35686\
        );

    \I__5237\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35683\
        );

    \I__5236\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35680\
        );

    \I__5235\ : InMux
    port map (
            O => \N__35686\,
            I => \N__35677\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__35683\,
            I => \N__35674\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__35680\,
            I => \N__35669\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__35677\,
            I => \N__35669\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__35674\,
            I => \c0.n13056\
        );

    \I__5230\ : Odrv12
    port map (
            O => \N__35669\,
            I => \c0.n13056\
        );

    \I__5229\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35659\
        );

    \I__5228\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35654\
        );

    \I__5227\ : InMux
    port map (
            O => \N__35662\,
            I => \N__35654\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__35659\,
            I => \N__35646\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__35654\,
            I => \N__35646\
        );

    \I__5224\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35641\
        );

    \I__5223\ : InMux
    port map (
            O => \N__35652\,
            I => \N__35641\
        );

    \I__5222\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35638\
        );

    \I__5221\ : Span4Mux_v
    port map (
            O => \N__35646\,
            I => \N__35634\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__35641\,
            I => \N__35631\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__35638\,
            I => \N__35628\
        );

    \I__5218\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35625\
        );

    \I__5217\ : Odrv4
    port map (
            O => \N__35634\,
            I => \c0.n63_adj_4235\
        );

    \I__5216\ : Odrv12
    port map (
            O => \N__35631\,
            I => \c0.n63_adj_4235\
        );

    \I__5215\ : Odrv4
    port map (
            O => \N__35628\,
            I => \c0.n63_adj_4235\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__35625\,
            I => \c0.n63_adj_4235\
        );

    \I__5213\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35611\
        );

    \I__5212\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35606\
        );

    \I__5211\ : InMux
    port map (
            O => \N__35614\,
            I => \N__35606\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__35611\,
            I => \N__35597\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__35606\,
            I => \N__35597\
        );

    \I__5208\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35592\
        );

    \I__5207\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35592\
        );

    \I__5206\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35589\
        );

    \I__5205\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35586\
        );

    \I__5204\ : Sp12to4
    port map (
            O => \N__35597\,
            I => \N__35577\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__35592\,
            I => \N__35577\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__35589\,
            I => \N__35577\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__35586\,
            I => \N__35577\
        );

    \I__5200\ : Odrv12
    port map (
            O => \N__35577\,
            I => \c0.n63_adj_4238\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__35574\,
            I => \c0.n2004_cascade_\
        );

    \I__5198\ : CascadeMux
    port map (
            O => \N__35571\,
            I => \N__35568\
        );

    \I__5197\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35565\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__35565\,
            I => \c0.n28_adj_4565\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__35562\,
            I => \N__35558\
        );

    \I__5194\ : CascadeMux
    port map (
            O => \N__35561\,
            I => \N__35555\
        );

    \I__5193\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35551\
        );

    \I__5192\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35546\
        );

    \I__5191\ : InMux
    port map (
            O => \N__35554\,
            I => \N__35546\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__35551\,
            I => \N__35539\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__35546\,
            I => \N__35539\
        );

    \I__5188\ : InMux
    port map (
            O => \N__35545\,
            I => \N__35536\
        );

    \I__5187\ : InMux
    port map (
            O => \N__35544\,
            I => \N__35533\
        );

    \I__5186\ : Span4Mux_v
    port map (
            O => \N__35539\,
            I => \N__35530\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__35536\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__35533\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__35530\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__5182\ : CascadeMux
    port map (
            O => \N__35523\,
            I => \c0.n7570_cascade_\
        );

    \I__5181\ : InMux
    port map (
            O => \N__35520\,
            I => \N__35514\
        );

    \I__5180\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35514\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__35514\,
            I => data_out_frame_6_4
        );

    \I__5178\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35508\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__35508\,
            I => \N__35504\
        );

    \I__5176\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35501\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__35504\,
            I => \N__35498\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__35501\,
            I => data_out_frame_7_4
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__35498\,
            I => data_out_frame_7_4
        );

    \I__5172\ : CascadeMux
    port map (
            O => \N__35493\,
            I => \c0.n13055_cascade_\
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__35490\,
            I => \n13058_cascade_\
        );

    \I__5170\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35483\
        );

    \I__5169\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35480\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__35483\,
            I => \N__35477\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__35480\,
            I => data_out_frame_7_6
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__35477\,
            I => data_out_frame_7_6
        );

    \I__5165\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35467\
        );

    \I__5164\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35464\
        );

    \I__5163\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35460\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__35467\,
            I => \N__35457\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__35464\,
            I => \N__35454\
        );

    \I__5160\ : CascadeMux
    port map (
            O => \N__35463\,
            I => \N__35450\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__35460\,
            I => \N__35443\
        );

    \I__5158\ : Span4Mux_v
    port map (
            O => \N__35457\,
            I => \N__35443\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__35454\,
            I => \N__35443\
        );

    \I__5156\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35438\
        );

    \I__5155\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35438\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__35443\,
            I => \N__35435\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__35438\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__35435\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__5151\ : CascadeMux
    port map (
            O => \N__35430\,
            I => \N__35427\
        );

    \I__5150\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35424\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__35424\,
            I => \N__35421\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__35421\,
            I => \c0.n5_adj_4477\
        );

    \I__5147\ : InMux
    port map (
            O => \N__35418\,
            I => \N__35412\
        );

    \I__5146\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35412\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__35412\,
            I => data_out_frame_13_4
        );

    \I__5144\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35406\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__35406\,
            I => \c0.n11_adj_4669\
        );

    \I__5142\ : InMux
    port map (
            O => \N__35403\,
            I => \N__35400\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__35400\,
            I => \N__35396\
        );

    \I__5140\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35393\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__35396\,
            I => \N__35390\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__35393\,
            I => data_out_frame_8_5
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__35390\,
            I => data_out_frame_8_5
        );

    \I__5136\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35382\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__35382\,
            I => \N__35378\
        );

    \I__5134\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35375\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__35378\,
            I => \N__35372\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__35375\,
            I => data_out_frame_7_5
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__35372\,
            I => data_out_frame_7_5
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__35367\,
            I => \N__35364\
        );

    \I__5129\ : InMux
    port map (
            O => \N__35364\,
            I => \N__35361\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__35361\,
            I => \N__35357\
        );

    \I__5127\ : InMux
    port map (
            O => \N__35360\,
            I => \N__35354\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__35357\,
            I => \N__35348\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__35354\,
            I => \N__35348\
        );

    \I__5124\ : InMux
    port map (
            O => \N__35353\,
            I => \N__35345\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__35348\,
            I => \N__35341\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__35345\,
            I => \N__35338\
        );

    \I__5121\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35335\
        );

    \I__5120\ : Span4Mux_v
    port map (
            O => \N__35341\,
            I => \N__35330\
        );

    \I__5119\ : Span4Mux_h
    port map (
            O => \N__35338\,
            I => \N__35330\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__35335\,
            I => encoder1_position_25
        );

    \I__5117\ : Odrv4
    port map (
            O => \N__35330\,
            I => encoder1_position_25
        );

    \I__5116\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35322\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__35322\,
            I => n2262
        );

    \I__5114\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35315\
        );

    \I__5113\ : CascadeMux
    port map (
            O => \N__35318\,
            I => \N__35312\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__35315\,
            I => \N__35309\
        );

    \I__5111\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35306\
        );

    \I__5110\ : Span4Mux_h
    port map (
            O => \N__35309\,
            I => \N__35303\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__35306\,
            I => data_out_frame_10_6
        );

    \I__5108\ : Odrv4
    port map (
            O => \N__35303\,
            I => data_out_frame_10_6
        );

    \I__5107\ : CascadeMux
    port map (
            O => \N__35298\,
            I => \N__35294\
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__35297\,
            I => \N__35291\
        );

    \I__5105\ : InMux
    port map (
            O => \N__35294\,
            I => \N__35288\
        );

    \I__5104\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35280\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__35288\,
            I => \N__35277\
        );

    \I__5102\ : InMux
    port map (
            O => \N__35287\,
            I => \N__35274\
        );

    \I__5101\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35269\
        );

    \I__5100\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35269\
        );

    \I__5099\ : InMux
    port map (
            O => \N__35284\,
            I => \N__35265\
        );

    \I__5098\ : CascadeMux
    port map (
            O => \N__35283\,
            I => \N__35262\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__35280\,
            I => \N__35258\
        );

    \I__5096\ : Span4Mux_v
    port map (
            O => \N__35277\,
            I => \N__35251\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__35274\,
            I => \N__35251\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__35269\,
            I => \N__35251\
        );

    \I__5093\ : InMux
    port map (
            O => \N__35268\,
            I => \N__35248\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__35265\,
            I => \N__35245\
        );

    \I__5091\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35240\
        );

    \I__5090\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35240\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__35258\,
            I => \N__35235\
        );

    \I__5088\ : Span4Mux_v
    port map (
            O => \N__35251\,
            I => \N__35235\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__35248\,
            I => encoder1_position_4
        );

    \I__5086\ : Odrv12
    port map (
            O => \N__35245\,
            I => encoder1_position_4
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__35240\,
            I => encoder1_position_4
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__35235\,
            I => encoder1_position_4
        );

    \I__5083\ : InMux
    port map (
            O => \N__35226\,
            I => \N__35222\
        );

    \I__5082\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35219\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__35222\,
            I => \N__35216\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__35219\,
            I => data_out_frame_8_0
        );

    \I__5079\ : Odrv4
    port map (
            O => \N__35216\,
            I => data_out_frame_8_0
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__35211\,
            I => \N__35208\
        );

    \I__5077\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35204\
        );

    \I__5076\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35201\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__35204\,
            I => \N__35198\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__35201\,
            I => \N__35195\
        );

    \I__5073\ : Span4Mux_v
    port map (
            O => \N__35198\,
            I => \N__35189\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__35195\,
            I => \N__35189\
        );

    \I__5071\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35185\
        );

    \I__5070\ : Span4Mux_v
    port map (
            O => \N__35189\,
            I => \N__35182\
        );

    \I__5069\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35179\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__35185\,
            I => encoder1_position_17
        );

    \I__5067\ : Odrv4
    port map (
            O => \N__35182\,
            I => encoder1_position_17
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__35179\,
            I => encoder1_position_17
        );

    \I__5065\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35169\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__35169\,
            I => \c0.n16_adj_4233\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__35166\,
            I => \N__35163\
        );

    \I__5062\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35159\
        );

    \I__5061\ : InMux
    port map (
            O => \N__35162\,
            I => \N__35156\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__35159\,
            I => \N__35153\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__35156\,
            I => data_out_frame_11_7
        );

    \I__5058\ : Odrv12
    port map (
            O => \N__35153\,
            I => data_out_frame_11_7
        );

    \I__5057\ : InMux
    port map (
            O => \N__35148\,
            I => \N__35144\
        );

    \I__5056\ : InMux
    port map (
            O => \N__35147\,
            I => \N__35141\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__35144\,
            I => \N__35138\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__35141\,
            I => data_out_frame_13_5
        );

    \I__5053\ : Odrv12
    port map (
            O => \N__35138\,
            I => data_out_frame_13_5
        );

    \I__5052\ : InMux
    port map (
            O => \N__35133\,
            I => \N__35129\
        );

    \I__5051\ : InMux
    port map (
            O => \N__35132\,
            I => \N__35126\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__35129\,
            I => \N__35123\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__35126\,
            I => \N__35120\
        );

    \I__5048\ : Span4Mux_v
    port map (
            O => \N__35123\,
            I => \N__35117\
        );

    \I__5047\ : Span4Mux_v
    port map (
            O => \N__35120\,
            I => \N__35113\
        );

    \I__5046\ : Span4Mux_v
    port map (
            O => \N__35117\,
            I => \N__35108\
        );

    \I__5045\ : InMux
    port map (
            O => \N__35116\,
            I => \N__35105\
        );

    \I__5044\ : Span4Mux_v
    port map (
            O => \N__35113\,
            I => \N__35102\
        );

    \I__5043\ : InMux
    port map (
            O => \N__35112\,
            I => \N__35099\
        );

    \I__5042\ : InMux
    port map (
            O => \N__35111\,
            I => \N__35096\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__35108\,
            I => encoder1_position_11
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__35105\,
            I => encoder1_position_11
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__35102\,
            I => encoder1_position_11
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__35099\,
            I => encoder1_position_11
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__35096\,
            I => encoder1_position_11
        );

    \I__5036\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35082\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__35082\,
            I => \N__35079\
        );

    \I__5034\ : Span4Mux_v
    port map (
            O => \N__35079\,
            I => \N__35075\
        );

    \I__5033\ : InMux
    port map (
            O => \N__35078\,
            I => \N__35072\
        );

    \I__5032\ : Span4Mux_h
    port map (
            O => \N__35075\,
            I => \N__35069\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__35072\,
            I => data_out_frame_12_3
        );

    \I__5030\ : Odrv4
    port map (
            O => \N__35069\,
            I => data_out_frame_12_3
        );

    \I__5029\ : CascadeMux
    port map (
            O => \N__35064\,
            I => \N__35061\
        );

    \I__5028\ : InMux
    port map (
            O => \N__35061\,
            I => \N__35057\
        );

    \I__5027\ : InMux
    port map (
            O => \N__35060\,
            I => \N__35054\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__35057\,
            I => \N__35051\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__35054\,
            I => data_out_frame_12_2
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__35051\,
            I => data_out_frame_12_2
        );

    \I__5023\ : InMux
    port map (
            O => \N__35046\,
            I => \N__35043\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__35043\,
            I => n2281
        );

    \I__5021\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35035\
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__35039\,
            I => \N__35029\
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__35038\,
            I => \N__35026\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__35035\,
            I => \N__35023\
        );

    \I__5017\ : InMux
    port map (
            O => \N__35034\,
            I => \N__35018\
        );

    \I__5016\ : InMux
    port map (
            O => \N__35033\,
            I => \N__35018\
        );

    \I__5015\ : InMux
    port map (
            O => \N__35032\,
            I => \N__35013\
        );

    \I__5014\ : InMux
    port map (
            O => \N__35029\,
            I => \N__35013\
        );

    \I__5013\ : InMux
    port map (
            O => \N__35026\,
            I => \N__35010\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__35023\,
            I => \N__35007\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__35018\,
            I => \N__35004\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__35013\,
            I => encoder1_position_10
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__35010\,
            I => encoder1_position_10
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__35007\,
            I => encoder1_position_10
        );

    \I__5007\ : Odrv12
    port map (
            O => \N__35004\,
            I => encoder1_position_10
        );

    \I__5006\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34992\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__34992\,
            I => \N__34988\
        );

    \I__5004\ : InMux
    port map (
            O => \N__34991\,
            I => \N__34985\
        );

    \I__5003\ : Span4Mux_h
    port map (
            O => \N__34988\,
            I => \N__34982\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__34985\,
            I => data_out_frame_5_6
        );

    \I__5001\ : Odrv4
    port map (
            O => \N__34982\,
            I => data_out_frame_5_6
        );

    \I__5000\ : InMux
    port map (
            O => \N__34977\,
            I => \N__34970\
        );

    \I__4999\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34970\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__34975\,
            I => \N__34967\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__34970\,
            I => \N__34964\
        );

    \I__4996\ : InMux
    port map (
            O => \N__34967\,
            I => \N__34960\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__34964\,
            I => \N__34956\
        );

    \I__4994\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34953\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__34960\,
            I => \N__34950\
        );

    \I__4992\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34947\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__34956\,
            I => \N__34944\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__34953\,
            I => encoder1_position_15
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__34950\,
            I => encoder1_position_15
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__34947\,
            I => encoder1_position_15
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__34944\,
            I => encoder1_position_15
        );

    \I__4986\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34932\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__34932\,
            I => \N__34929\
        );

    \I__4984\ : Span4Mux_v
    port map (
            O => \N__34929\,
            I => \N__34925\
        );

    \I__4983\ : InMux
    port map (
            O => \N__34928\,
            I => \N__34922\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__34925\,
            I => \N__34919\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__34922\,
            I => data_out_frame_12_7
        );

    \I__4980\ : Odrv4
    port map (
            O => \N__34919\,
            I => data_out_frame_12_7
        );

    \I__4979\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34911\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__34911\,
            I => n2263
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__34908\,
            I => \N__34905\
        );

    \I__4976\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34902\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__34902\,
            I => n2264
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__34899\,
            I => \N__34896\
        );

    \I__4973\ : InMux
    port map (
            O => \N__34896\,
            I => \N__34892\
        );

    \I__4972\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34889\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__34892\,
            I => \N__34885\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__34889\,
            I => \N__34881\
        );

    \I__4969\ : InMux
    port map (
            O => \N__34888\,
            I => \N__34878\
        );

    \I__4968\ : Span4Mux_v
    port map (
            O => \N__34885\,
            I => \N__34875\
        );

    \I__4967\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34872\
        );

    \I__4966\ : Span4Mux_v
    port map (
            O => \N__34881\,
            I => \N__34869\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__34878\,
            I => encoder1_position_27
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__34875\,
            I => encoder1_position_27
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__34872\,
            I => encoder1_position_27
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__34869\,
            I => encoder1_position_27
        );

    \I__4961\ : CascadeMux
    port map (
            O => \N__34860\,
            I => \N__34857\
        );

    \I__4960\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34853\
        );

    \I__4959\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34850\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34847\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__34850\,
            I => data_out_frame_5_3
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__34847\,
            I => data_out_frame_5_3
        );

    \I__4955\ : InMux
    port map (
            O => \N__34842\,
            I => \N__34838\
        );

    \I__4954\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34835\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__34838\,
            I => \N__34832\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__34835\,
            I => data_out_frame_7_1
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__34832\,
            I => data_out_frame_7_1
        );

    \I__4950\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34824\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__34824\,
            I => n2270
        );

    \I__4948\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34818\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__34818\,
            I => \N__34811\
        );

    \I__4946\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34806\
        );

    \I__4945\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34806\
        );

    \I__4944\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34800\
        );

    \I__4943\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34800\
        );

    \I__4942\ : Span4Mux_v
    port map (
            O => \N__34811\,
            I => \N__34795\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__34806\,
            I => \N__34795\
        );

    \I__4940\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34792\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__34800\,
            I => \c0.n13395\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__34795\,
            I => \c0.n13395\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__34792\,
            I => \c0.n13395\
        );

    \I__4936\ : CascadeMux
    port map (
            O => \N__34785\,
            I => \N__34782\
        );

    \I__4935\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34777\
        );

    \I__4934\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34772\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__34780\,
            I => \N__34769\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__34777\,
            I => \N__34766\
        );

    \I__4931\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34762\
        );

    \I__4930\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34759\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__34772\,
            I => \N__34756\
        );

    \I__4928\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34753\
        );

    \I__4927\ : Span4Mux_h
    port map (
            O => \N__34766\,
            I => \N__34750\
        );

    \I__4926\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34747\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34741\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__34759\,
            I => \N__34741\
        );

    \I__4923\ : Span4Mux_v
    port map (
            O => \N__34756\,
            I => \N__34738\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__34753\,
            I => \N__34734\
        );

    \I__4921\ : Span4Mux_v
    port map (
            O => \N__34750\,
            I => \N__34729\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__34747\,
            I => \N__34729\
        );

    \I__4919\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34726\
        );

    \I__4918\ : Span4Mux_v
    port map (
            O => \N__34741\,
            I => \N__34721\
        );

    \I__4917\ : Span4Mux_h
    port map (
            O => \N__34738\,
            I => \N__34721\
        );

    \I__4916\ : InMux
    port map (
            O => \N__34737\,
            I => \N__34718\
        );

    \I__4915\ : Span4Mux_h
    port map (
            O => \N__34734\,
            I => \N__34715\
        );

    \I__4914\ : Span4Mux_v
    port map (
            O => \N__34729\,
            I => \N__34712\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__34726\,
            I => \N__34709\
        );

    \I__4912\ : Span4Mux_h
    port map (
            O => \N__34721\,
            I => \N__34706\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__34718\,
            I => encoder1_position_1
        );

    \I__4910\ : Odrv4
    port map (
            O => \N__34715\,
            I => encoder1_position_1
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__34712\,
            I => encoder1_position_1
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__34709\,
            I => encoder1_position_1
        );

    \I__4907\ : Odrv4
    port map (
            O => \N__34706\,
            I => encoder1_position_1
        );

    \I__4906\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34692\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__34692\,
            I => \N__34688\
        );

    \I__4904\ : InMux
    port map (
            O => \N__34691\,
            I => \N__34685\
        );

    \I__4903\ : Span4Mux_h
    port map (
            O => \N__34688\,
            I => \N__34682\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__34685\,
            I => data_out_frame_9_0
        );

    \I__4901\ : Odrv4
    port map (
            O => \N__34682\,
            I => data_out_frame_9_0
        );

    \I__4900\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34674\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__34674\,
            I => \N__34670\
        );

    \I__4898\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34667\
        );

    \I__4897\ : Span4Mux_v
    port map (
            O => \N__34670\,
            I => \N__34664\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__34667\,
            I => data_out_frame_5_4
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__34664\,
            I => data_out_frame_5_4
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__34659\,
            I => \N__34656\
        );

    \I__4893\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34651\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__34655\,
            I => \N__34646\
        );

    \I__4891\ : InMux
    port map (
            O => \N__34654\,
            I => \N__34643\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__34651\,
            I => \N__34640\
        );

    \I__4889\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34637\
        );

    \I__4888\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34634\
        );

    \I__4887\ : InMux
    port map (
            O => \N__34646\,
            I => \N__34631\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__34643\,
            I => \N__34628\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__34640\,
            I => \N__34623\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__34637\,
            I => \N__34623\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__34634\,
            I => encoder1_position_22
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__34631\,
            I => encoder1_position_22
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__34628\,
            I => encoder1_position_22
        );

    \I__4880\ : Odrv4
    port map (
            O => \N__34623\,
            I => encoder1_position_22
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__34614\,
            I => \N__34611\
        );

    \I__4878\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34606\
        );

    \I__4877\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34603\
        );

    \I__4876\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34599\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__34606\,
            I => \N__34596\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__34603\,
            I => \N__34590\
        );

    \I__4873\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34587\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__34599\,
            I => \N__34584\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__34596\,
            I => \N__34581\
        );

    \I__4870\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34578\
        );

    \I__4869\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34575\
        );

    \I__4868\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34572\
        );

    \I__4867\ : Span12Mux_s7_v
    port map (
            O => \N__34590\,
            I => \N__34569\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__34587\,
            I => \N__34566\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__34584\,
            I => \N__34561\
        );

    \I__4864\ : Span4Mux_h
    port map (
            O => \N__34581\,
            I => \N__34561\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__34578\,
            I => encoder1_position_7
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__34575\,
            I => encoder1_position_7
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__34572\,
            I => encoder1_position_7
        );

    \I__4860\ : Odrv12
    port map (
            O => \N__34569\,
            I => encoder1_position_7
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__34566\,
            I => encoder1_position_7
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__34561\,
            I => encoder1_position_7
        );

    \I__4857\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34545\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__34545\,
            I => \N__34541\
        );

    \I__4855\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34538\
        );

    \I__4854\ : Span4Mux_h
    port map (
            O => \N__34541\,
            I => \N__34535\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__34538\,
            I => data_out_frame_7_2
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__34535\,
            I => data_out_frame_7_2
        );

    \I__4851\ : InMux
    port map (
            O => \N__34530\,
            I => \N__34527\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__34527\,
            I => \N__34524\
        );

    \I__4849\ : Span4Mux_v
    port map (
            O => \N__34524\,
            I => \N__34521\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__34521\,
            I => \c0.data_out_frame_29_0\
        );

    \I__4847\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34515\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__34515\,
            I => \c0.data_out_frame_28_0\
        );

    \I__4845\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34509\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__34509\,
            I => \N__34506\
        );

    \I__4843\ : Span12Mux_v
    port map (
            O => \N__34506\,
            I => \N__34503\
        );

    \I__4842\ : Odrv12
    port map (
            O => \N__34503\,
            I => \c0.n26_adj_4570\
        );

    \I__4841\ : CascadeMux
    port map (
            O => \N__34500\,
            I => \c0.n10529_cascade_\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__34497\,
            I => \c0.n22489_cascade_\
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__34494\,
            I => \c0.n21416_cascade_\
        );

    \I__4838\ : InMux
    port map (
            O => \N__34491\,
            I => \N__34488\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__34488\,
            I => \N__34485\
        );

    \I__4836\ : Span4Mux_v
    port map (
            O => \N__34485\,
            I => \N__34482\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__34482\,
            I => \c0.n24530\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__34479\,
            I => \c0.n22671_cascade_\
        );

    \I__4833\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34473\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__34473\,
            I => \c0.n20230\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__34470\,
            I => \c0.n20230_cascade_\
        );

    \I__4830\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34464\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__34464\,
            I => \N__34461\
        );

    \I__4828\ : Sp12to4
    port map (
            O => \N__34461\,
            I => \N__34458\
        );

    \I__4827\ : Odrv12
    port map (
            O => \N__34458\,
            I => \c0.data_out_frame_29_5\
        );

    \I__4826\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34452\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__34452\,
            I => \c0.n21457\
        );

    \I__4824\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34445\
        );

    \I__4823\ : InMux
    port map (
            O => \N__34448\,
            I => \N__34442\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__34445\,
            I => \c0.n21489\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__34442\,
            I => \c0.n21489\
        );

    \I__4820\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34434\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34429\
        );

    \I__4818\ : InMux
    port map (
            O => \N__34433\,
            I => \N__34426\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__34432\,
            I => \N__34422\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__34429\,
            I => \N__34416\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__34426\,
            I => \N__34416\
        );

    \I__4814\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34413\
        );

    \I__4813\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34410\
        );

    \I__4812\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34407\
        );

    \I__4811\ : Span4Mux_v
    port map (
            O => \N__34416\,
            I => \N__34404\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__34413\,
            I => \N__34401\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__34410\,
            I => \N__34398\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__34407\,
            I => encoder1_position_6
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__34404\,
            I => encoder1_position_6
        );

    \I__4806\ : Odrv4
    port map (
            O => \N__34401\,
            I => encoder1_position_6
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__34398\,
            I => encoder1_position_6
        );

    \I__4804\ : InMux
    port map (
            O => \N__34389\,
            I => \N__34386\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__34386\,
            I => \N__34383\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__34383\,
            I => \c0.n20461\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__34380\,
            I => \c0.n21330_cascade_\
        );

    \I__4800\ : InMux
    port map (
            O => \N__34377\,
            I => \N__34374\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__34374\,
            I => \c0.n6_adj_4331\
        );

    \I__4798\ : InMux
    port map (
            O => \N__34371\,
            I => \N__34368\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__34368\,
            I => \N__34364\
        );

    \I__4796\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34361\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__34364\,
            I => \c0.n22414\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__34361\,
            I => \c0.n22414\
        );

    \I__4793\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34353\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__34353\,
            I => \N__34349\
        );

    \I__4791\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34346\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__34349\,
            I => \N__34339\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__34346\,
            I => \N__34339\
        );

    \I__4788\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34336\
        );

    \I__4787\ : InMux
    port map (
            O => \N__34344\,
            I => \N__34333\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__34339\,
            I => \N__34330\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__34336\,
            I => n21307
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__34333\,
            I => n21307
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__34330\,
            I => n21307
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__34323\,
            I => \c0.n6_adj_4215_cascade_\
        );

    \I__4781\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34317\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__34317\,
            I => \N__34313\
        );

    \I__4779\ : InMux
    port map (
            O => \N__34316\,
            I => \N__34310\
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__34313\,
            I => \c0.n22268\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__34310\,
            I => \c0.n22268\
        );

    \I__4776\ : CascadeMux
    port map (
            O => \N__34305\,
            I => \N__34302\
        );

    \I__4775\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34299\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__34299\,
            I => \N__34296\
        );

    \I__4773\ : Span4Mux_h
    port map (
            O => \N__34296\,
            I => \N__34293\
        );

    \I__4772\ : Span4Mux_h
    port map (
            O => \N__34293\,
            I => \N__34290\
        );

    \I__4771\ : Odrv4
    port map (
            O => \N__34290\,
            I => \c0.n5_adj_4660\
        );

    \I__4770\ : InMux
    port map (
            O => \N__34287\,
            I => \N__34284\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__34284\,
            I => \N__34281\
        );

    \I__4768\ : Span12Mux_v
    port map (
            O => \N__34281\,
            I => \N__34278\
        );

    \I__4767\ : Odrv12
    port map (
            O => \N__34278\,
            I => \c0.n6_adj_4659\
        );

    \I__4766\ : InMux
    port map (
            O => \N__34275\,
            I => \N__34272\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__34272\,
            I => \N__34269\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__34269\,
            I => \N__34266\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__34266\,
            I => \c0.n24755\
        );

    \I__4762\ : InMux
    port map (
            O => \N__34263\,
            I => \N__34259\
        );

    \I__4761\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34256\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__34259\,
            I => \N__34251\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__34256\,
            I => \N__34251\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__34251\,
            I => \N__34248\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__34248\,
            I => \c0.n22330\
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__34245\,
            I => \c0.n19_adj_4693_cascade_\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__34242\,
            I => \c0.n6_adj_4691_cascade_\
        );

    \I__4754\ : InMux
    port map (
            O => \N__34239\,
            I => \N__34236\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__34236\,
            I => \c0.n21_adj_4692\
        );

    \I__4752\ : InMux
    port map (
            O => \N__34233\,
            I => \N__34230\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__34230\,
            I => \N__34227\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__34227\,
            I => \N__34224\
        );

    \I__4749\ : Span4Mux_v
    port map (
            O => \N__34224\,
            I => \N__34221\
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__34221\,
            I => n2274
        );

    \I__4747\ : InMux
    port map (
            O => \N__34218\,
            I => \N__34215\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__34215\,
            I => \N__34212\
        );

    \I__4745\ : Span4Mux_v
    port map (
            O => \N__34212\,
            I => \N__34209\
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__34209\,
            I => n2283
        );

    \I__4743\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34202\
        );

    \I__4742\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34199\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__34202\,
            I => \N__34196\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__34199\,
            I => \c0.n22656\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__34196\,
            I => \c0.n22656\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__34191\,
            I => \N__34188\
        );

    \I__4737\ : InMux
    port map (
            O => \N__34188\,
            I => \N__34185\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__34185\,
            I => \N__34182\
        );

    \I__4735\ : Span4Mux_h
    port map (
            O => \N__34182\,
            I => \N__34178\
        );

    \I__4734\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34175\
        );

    \I__4733\ : Odrv4
    port map (
            O => \N__34178\,
            I => \c0.n22800\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__34175\,
            I => \c0.n22800\
        );

    \I__4731\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34167\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34164\
        );

    \I__4729\ : Odrv12
    port map (
            O => \N__34164\,
            I => \c0.n10_adj_4339\
        );

    \I__4728\ : CascadeMux
    port map (
            O => \N__34161\,
            I => \c0.n14_adj_4338_cascade_\
        );

    \I__4727\ : CascadeMux
    port map (
            O => \N__34158\,
            I => \c0.n20461_cascade_\
        );

    \I__4726\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34151\
        );

    \I__4725\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34147\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__34151\,
            I => \N__34144\
        );

    \I__4723\ : InMux
    port map (
            O => \N__34150\,
            I => \N__34141\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__34147\,
            I => \N__34138\
        );

    \I__4721\ : Span4Mux_v
    port map (
            O => \N__34144\,
            I => \N__34133\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__34141\,
            I => \N__34130\
        );

    \I__4719\ : Span4Mux_h
    port map (
            O => \N__34138\,
            I => \N__34127\
        );

    \I__4718\ : InMux
    port map (
            O => \N__34137\,
            I => \N__34122\
        );

    \I__4717\ : InMux
    port map (
            O => \N__34136\,
            I => \N__34122\
        );

    \I__4716\ : Odrv4
    port map (
            O => \N__34133\,
            I => \c0.n20388\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__34130\,
            I => \c0.n20388\
        );

    \I__4714\ : Odrv4
    port map (
            O => \N__34127\,
            I => \c0.n20388\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__34122\,
            I => \c0.n20388\
        );

    \I__4712\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34110\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__34110\,
            I => \N__34106\
        );

    \I__4710\ : InMux
    port map (
            O => \N__34109\,
            I => \N__34103\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__34106\,
            I => \c0.n22408\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__34103\,
            I => \c0.n22408\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__34098\,
            I => \N__34095\
        );

    \I__4706\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34092\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__34087\
        );

    \I__4704\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34084\
        );

    \I__4703\ : InMux
    port map (
            O => \N__34090\,
            I => \N__34080\
        );

    \I__4702\ : Span4Mux_v
    port map (
            O => \N__34087\,
            I => \N__34075\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__34084\,
            I => \N__34075\
        );

    \I__4700\ : CascadeMux
    port map (
            O => \N__34083\,
            I => \N__34070\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__34080\,
            I => \N__34067\
        );

    \I__4698\ : Span4Mux_h
    port map (
            O => \N__34075\,
            I => \N__34064\
        );

    \I__4697\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34061\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__34073\,
            I => \N__34058\
        );

    \I__4695\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34055\
        );

    \I__4694\ : Sp12to4
    port map (
            O => \N__34067\,
            I => \N__34050\
        );

    \I__4693\ : Sp12to4
    port map (
            O => \N__34064\,
            I => \N__34050\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__34061\,
            I => \N__34047\
        );

    \I__4691\ : InMux
    port map (
            O => \N__34058\,
            I => \N__34044\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__34055\,
            I => \N__34041\
        );

    \I__4689\ : Span12Mux_v
    port map (
            O => \N__34050\,
            I => \N__34038\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__34047\,
            I => encoder1_position_16
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__34044\,
            I => encoder1_position_16
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__34041\,
            I => encoder1_position_16
        );

    \I__4685\ : Odrv12
    port map (
            O => \N__34038\,
            I => encoder1_position_16
        );

    \I__4684\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34024\
        );

    \I__4683\ : InMux
    port map (
            O => \N__34028\,
            I => \N__34021\
        );

    \I__4682\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34018\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__34024\,
            I => \c0.n20449\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__34021\,
            I => \c0.n20449\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__34018\,
            I => \c0.n20449\
        );

    \I__4678\ : InMux
    port map (
            O => \N__34011\,
            I => \N__34008\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__34005\,
            I => \c0.n10_adj_4374\
        );

    \I__4675\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33999\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__33999\,
            I => \c0.data_out_frame_29__7__N_855\
        );

    \I__4673\ : CascadeMux
    port map (
            O => \N__33996\,
            I => \N__33990\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__33995\,
            I => \N__33987\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__33994\,
            I => \N__33984\
        );

    \I__4670\ : InMux
    port map (
            O => \N__33993\,
            I => \N__33981\
        );

    \I__4669\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33978\
        );

    \I__4668\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33973\
        );

    \I__4667\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33973\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__33981\,
            I => \N__33970\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__33978\,
            I => \N__33967\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__33973\,
            I => \N__33964\
        );

    \I__4663\ : Span4Mux_h
    port map (
            O => \N__33970\,
            I => \N__33961\
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__33967\,
            I => \c0.n13384\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__33964\,
            I => \c0.n13384\
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__33961\,
            I => \c0.n13384\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__33954\,
            I => \N__33950\
        );

    \I__4658\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33947\
        );

    \I__4657\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33943\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__33947\,
            I => \N__33939\
        );

    \I__4655\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33936\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__33943\,
            I => \N__33933\
        );

    \I__4653\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33930\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__33939\,
            I => \N__33925\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__33936\,
            I => \N__33925\
        );

    \I__4650\ : Span4Mux_h
    port map (
            O => \N__33933\,
            I => \N__33922\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__33930\,
            I => encoder1_position_0
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__33925\,
            I => encoder1_position_0
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__33922\,
            I => encoder1_position_0
        );

    \I__4646\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33912\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__33912\,
            I => \N__33908\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__33911\,
            I => \N__33905\
        );

    \I__4643\ : Span4Mux_v
    port map (
            O => \N__33908\,
            I => \N__33902\
        );

    \I__4642\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33899\
        );

    \I__4641\ : Sp12to4
    port map (
            O => \N__33902\,
            I => \N__33896\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__33899\,
            I => \c0.n22611\
        );

    \I__4639\ : Odrv12
    port map (
            O => \N__33896\,
            I => \c0.n22611\
        );

    \I__4638\ : InMux
    port map (
            O => \N__33891\,
            I => \N__33888\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__33888\,
            I => \c0.n10_adj_4274\
        );

    \I__4636\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \N__33881\
        );

    \I__4635\ : InMux
    port map (
            O => \N__33884\,
            I => \N__33878\
        );

    \I__4634\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33875\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__33878\,
            I => \c0.n22791\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__33875\,
            I => \c0.n22791\
        );

    \I__4631\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33866\
        );

    \I__4630\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33863\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__33866\,
            I => \N__33860\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__33863\,
            I => \c0.n22466\
        );

    \I__4627\ : Odrv4
    port map (
            O => \N__33860\,
            I => \c0.n22466\
        );

    \I__4626\ : InMux
    port map (
            O => \N__33855\,
            I => \N__33847\
        );

    \I__4625\ : InMux
    port map (
            O => \N__33854\,
            I => \N__33847\
        );

    \I__4624\ : InMux
    port map (
            O => \N__33853\,
            I => \N__33844\
        );

    \I__4623\ : InMux
    port map (
            O => \N__33852\,
            I => \N__33841\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__33847\,
            I => \N__33838\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__33844\,
            I => \N__33835\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__33841\,
            I => \c0.n13121\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__33838\,
            I => \c0.n13121\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__33835\,
            I => \c0.n13121\
        );

    \I__4617\ : InMux
    port map (
            O => \N__33828\,
            I => \N__33825\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__33825\,
            I => \N__33822\
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__33822\,
            I => \c0.n34_adj_4328\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__33819\,
            I => \c0.n30_adj_4326_cascade_\
        );

    \I__4613\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33813\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__33813\,
            I => \c0.n29_adj_4329\
        );

    \I__4611\ : CascadeMux
    port map (
            O => \N__33810\,
            I => \N__33807\
        );

    \I__4610\ : InMux
    port map (
            O => \N__33807\,
            I => \N__33803\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__33806\,
            I => \N__33800\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__33803\,
            I => \N__33795\
        );

    \I__4607\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33792\
        );

    \I__4606\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33789\
        );

    \I__4605\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33786\
        );

    \I__4604\ : Span12Mux_v
    port map (
            O => \N__33795\,
            I => \N__33781\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__33792\,
            I => \N__33781\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__33789\,
            I => \N__33778\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__33786\,
            I => encoder1_position_20
        );

    \I__4600\ : Odrv12
    port map (
            O => \N__33781\,
            I => encoder1_position_20
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__33778\,
            I => encoder1_position_20
        );

    \I__4598\ : CascadeMux
    port map (
            O => \N__33771\,
            I => \N__33768\
        );

    \I__4597\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33765\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__33765\,
            I => \c0.n22788\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__33762\,
            I => \c0.n22788_cascade_\
        );

    \I__4594\ : SRMux
    port map (
            O => \N__33759\,
            I => \N__33756\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__33756\,
            I => \N__33753\
        );

    \I__4592\ : Span4Mux_h
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__33750\,
            I => \c0.n21637\
        );

    \I__4590\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33744\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__33744\,
            I => \c0.n22638\
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__33741\,
            I => \c0.n22831_cascade_\
        );

    \I__4587\ : InMux
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33732\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__33732\,
            I => \c0.n20_adj_4321\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__33729\,
            I => \c0.n13_adj_4320_cascade_\
        );

    \I__4583\ : InMux
    port map (
            O => \N__33726\,
            I => \N__33723\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__33723\,
            I => \c0.n14_adj_4319\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__33720\,
            I => \c0.n28_adj_4322_cascade_\
        );

    \I__4580\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33712\
        );

    \I__4579\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33707\
        );

    \I__4578\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33707\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__33712\,
            I => \c0.n12488\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__33707\,
            I => \c0.n12488\
        );

    \I__4575\ : InMux
    port map (
            O => \N__33702\,
            I => \N__33697\
        );

    \I__4574\ : CascadeMux
    port map (
            O => \N__33701\,
            I => \N__33694\
        );

    \I__4573\ : CascadeMux
    port map (
            O => \N__33700\,
            I => \N__33690\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__33697\,
            I => \N__33687\
        );

    \I__4571\ : InMux
    port map (
            O => \N__33694\,
            I => \N__33683\
        );

    \I__4570\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33678\
        );

    \I__4569\ : InMux
    port map (
            O => \N__33690\,
            I => \N__33678\
        );

    \I__4568\ : Span4Mux_v
    port map (
            O => \N__33687\,
            I => \N__33675\
        );

    \I__4567\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33672\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__33683\,
            I => \N__33668\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__33678\,
            I => \N__33665\
        );

    \I__4564\ : Span4Mux_v
    port map (
            O => \N__33675\,
            I => \N__33662\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__33672\,
            I => \N__33659\
        );

    \I__4562\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33656\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__33668\,
            I => \N__33653\
        );

    \I__4560\ : Span4Mux_h
    port map (
            O => \N__33665\,
            I => \N__33650\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__33662\,
            I => \N__33645\
        );

    \I__4558\ : Span4Mux_v
    port map (
            O => \N__33659\,
            I => \N__33645\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__33656\,
            I => encoder1_position_14
        );

    \I__4556\ : Odrv4
    port map (
            O => \N__33653\,
            I => encoder1_position_14
        );

    \I__4555\ : Odrv4
    port map (
            O => \N__33650\,
            I => encoder1_position_14
        );

    \I__4554\ : Odrv4
    port map (
            O => \N__33645\,
            I => encoder1_position_14
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__33636\,
            I => \c0.n20318_cascade_\
        );

    \I__4552\ : SRMux
    port map (
            O => \N__33633\,
            I => \N__33630\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33627\
        );

    \I__4550\ : Span4Mux_h
    port map (
            O => \N__33627\,
            I => \N__33624\
        );

    \I__4549\ : Odrv4
    port map (
            O => \N__33624\,
            I => \c0.n21579\
        );

    \I__4548\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33615\
        );

    \I__4547\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33615\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__33615\,
            I => \c0.n4_adj_4678\
        );

    \I__4545\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33607\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__33611\,
            I => \N__33604\
        );

    \I__4543\ : CascadeMux
    port map (
            O => \N__33610\,
            I => \N__33601\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33597\
        );

    \I__4541\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33594\
        );

    \I__4540\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33589\
        );

    \I__4539\ : InMux
    port map (
            O => \N__33600\,
            I => \N__33586\
        );

    \I__4538\ : Span4Mux_h
    port map (
            O => \N__33597\,
            I => \N__33581\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__33594\,
            I => \N__33581\
        );

    \I__4536\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33578\
        );

    \I__4535\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33575\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33572\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__33586\,
            I => \N__33569\
        );

    \I__4532\ : Span4Mux_v
    port map (
            O => \N__33581\,
            I => \N__33566\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__33578\,
            I => \N__33563\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__33575\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__4529\ : Odrv12
    port map (
            O => \N__33572\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__4528\ : Odrv12
    port map (
            O => \N__33569\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__4527\ : Odrv4
    port map (
            O => \N__33566\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__33563\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__4525\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33548\
        );

    \I__4524\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33545\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__33548\,
            I => \N__33538\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__33545\,
            I => \N__33538\
        );

    \I__4521\ : InMux
    port map (
            O => \N__33544\,
            I => \N__33535\
        );

    \I__4520\ : InMux
    port map (
            O => \N__33543\,
            I => \N__33532\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__33538\,
            I => \c0.n22131\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__33535\,
            I => \c0.n22131\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__33532\,
            I => \c0.n22131\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__33525\,
            I => \N__33520\
        );

    \I__4515\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33517\
        );

    \I__4514\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33514\
        );

    \I__4513\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33511\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__33517\,
            I => \N__33508\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__33514\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__33511\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__33508\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__4508\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33496\
        );

    \I__4507\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33491\
        );

    \I__4506\ : InMux
    port map (
            O => \N__33499\,
            I => \N__33491\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__33496\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__33491\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__4503\ : SRMux
    port map (
            O => \N__33486\,
            I => \N__33483\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__33483\,
            I => \c0.n21625\
        );

    \I__4501\ : SRMux
    port map (
            O => \N__33480\,
            I => \N__33477\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__33477\,
            I => \N__33474\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__33474\,
            I => \c0.n8_adj_4561\
        );

    \I__4498\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33467\
        );

    \I__4497\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33463\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__33467\,
            I => \N__33460\
        );

    \I__4495\ : InMux
    port map (
            O => \N__33466\,
            I => \N__33457\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__33463\,
            I => \N__33454\
        );

    \I__4493\ : Span4Mux_h
    port map (
            O => \N__33460\,
            I => \N__33451\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__33457\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__4491\ : Odrv12
    port map (
            O => \N__33454\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__33451\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__4489\ : SRMux
    port map (
            O => \N__33444\,
            I => \N__33441\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__33441\,
            I => \N__33438\
        );

    \I__4487\ : Odrv12
    port map (
            O => \N__33438\,
            I => \c0.n8_adj_4558\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__33435\,
            I => \c0.data_out_frame_29_7_N_1482_0_cascade_\
        );

    \I__4485\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33429\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__33429\,
            I => \c0.n6_adj_4495\
        );

    \I__4483\ : InMux
    port map (
            O => \N__33426\,
            I => \N__33423\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__33423\,
            I => \c0.n14784\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__33420\,
            I => \c0.n9706_cascade_\
        );

    \I__4480\ : CascadeMux
    port map (
            O => \N__33417\,
            I => \c0.n6_cascade_\
        );

    \I__4479\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33410\
        );

    \I__4478\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33407\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__33410\,
            I => \N__33402\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__33407\,
            I => \N__33402\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__33402\,
            I => data_out_frame_9_6
        );

    \I__4474\ : InMux
    port map (
            O => \N__33399\,
            I => \N__33395\
        );

    \I__4473\ : InMux
    port map (
            O => \N__33398\,
            I => \N__33392\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__33395\,
            I => data_out_frame_6_6
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__33392\,
            I => data_out_frame_6_6
        );

    \I__4470\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33384\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__4468\ : Span4Mux_h
    port map (
            O => \N__33381\,
            I => \N__33377\
        );

    \I__4467\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33374\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__33377\,
            I => n14247
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__33374\,
            I => n14247
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__33369\,
            I => \N__33366\
        );

    \I__4463\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33363\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__33363\,
            I => \N__33359\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__33362\,
            I => \N__33356\
        );

    \I__4460\ : Span4Mux_v
    port map (
            O => \N__33359\,
            I => \N__33353\
        );

    \I__4459\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33350\
        );

    \I__4458\ : Span4Mux_v
    port map (
            O => \N__33353\,
            I => \N__33347\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__33350\,
            I => data_out_frame_0_4
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__33347\,
            I => data_out_frame_0_4
        );

    \I__4455\ : InMux
    port map (
            O => \N__33342\,
            I => \N__33338\
        );

    \I__4454\ : InMux
    port map (
            O => \N__33341\,
            I => \N__33335\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__33338\,
            I => \N__33332\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__33335\,
            I => data_out_frame_9_2
        );

    \I__4451\ : Odrv4
    port map (
            O => \N__33332\,
            I => data_out_frame_9_2
        );

    \I__4450\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33323\
        );

    \I__4449\ : InMux
    port map (
            O => \N__33326\,
            I => \N__33320\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__33323\,
            I => data_out_frame_11_4
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__33320\,
            I => data_out_frame_11_4
        );

    \I__4446\ : InMux
    port map (
            O => \N__33315\,
            I => \N__33312\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__33312\,
            I => \N__33308\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__33311\,
            I => \N__33305\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__33308\,
            I => \N__33302\
        );

    \I__4442\ : InMux
    port map (
            O => \N__33305\,
            I => \N__33299\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__33302\,
            I => \N__33296\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__33299\,
            I => data_out_frame_13_2
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__33296\,
            I => data_out_frame_13_2
        );

    \I__4438\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__33288\,
            I => \c0.n12976\
        );

    \I__4436\ : CascadeMux
    port map (
            O => \N__33285\,
            I => \c0.n12976_cascade_\
        );

    \I__4435\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33279\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__33279\,
            I => \N__33276\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__33276\,
            I => \N__33273\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__33273\,
            I => n2275
        );

    \I__4431\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33266\
        );

    \I__4430\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33263\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__33266\,
            I => data_out_frame_10_0
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__33263\,
            I => data_out_frame_10_0
        );

    \I__4427\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33255\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33251\
        );

    \I__4425\ : InMux
    port map (
            O => \N__33254\,
            I => \N__33248\
        );

    \I__4424\ : Span4Mux_h
    port map (
            O => \N__33251\,
            I => \N__33245\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__33248\,
            I => data_out_frame_10_4
        );

    \I__4422\ : Odrv4
    port map (
            O => \N__33245\,
            I => data_out_frame_10_4
        );

    \I__4421\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33237\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__33237\,
            I => \c0.n24783\
        );

    \I__4419\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33230\
        );

    \I__4418\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33227\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__33230\,
            I => \N__33224\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__33227\,
            I => data_out_frame_6_0
        );

    \I__4415\ : Odrv12
    port map (
            O => \N__33224\,
            I => data_out_frame_6_0
        );

    \I__4414\ : CascadeMux
    port map (
            O => \N__33219\,
            I => \N__33216\
        );

    \I__4413\ : InMux
    port map (
            O => \N__33216\,
            I => \N__33212\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__33215\,
            I => \N__33209\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__33212\,
            I => \N__33206\
        );

    \I__4410\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33203\
        );

    \I__4409\ : Odrv12
    port map (
            O => \N__33206\,
            I => \c0.tx_transmit_N_3650\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__33203\,
            I => \c0.tx_transmit_N_3650\
        );

    \I__4407\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33195\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__33195\,
            I => \N__33192\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__33192\,
            I => \N__33189\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__33189\,
            I => \c0.n24888\
        );

    \I__4403\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33182\
        );

    \I__4402\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33179\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__33182\,
            I => \N__33174\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__33179\,
            I => \N__33174\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__33174\,
            I => data_out_frame_12_0
        );

    \I__4398\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33168\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__33168\,
            I => \N__33165\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__33165\,
            I => \N__33161\
        );

    \I__4395\ : InMux
    port map (
            O => \N__33164\,
            I => \N__33158\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__33161\,
            I => \N__33155\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__33158\,
            I => data_out_frame_12_1
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__33155\,
            I => data_out_frame_12_1
        );

    \I__4391\ : InMux
    port map (
            O => \N__33150\,
            I => \quad_counter1.n19759\
        );

    \I__4390\ : InMux
    port map (
            O => \N__33147\,
            I => \quad_counter1.n19760\
        );

    \I__4389\ : InMux
    port map (
            O => \N__33144\,
            I => \quad_counter1.n19761\
        );

    \I__4388\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33126\
        );

    \I__4387\ : CascadeMux
    port map (
            O => \N__33140\,
            I => \N__33122\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__33139\,
            I => \N__33118\
        );

    \I__4385\ : CascadeMux
    port map (
            O => \N__33138\,
            I => \N__33114\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__33137\,
            I => \N__33110\
        );

    \I__4383\ : CascadeMux
    port map (
            O => \N__33136\,
            I => \N__33106\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__33135\,
            I => \N__33102\
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__33134\,
            I => \N__33098\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__33133\,
            I => \N__33094\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__33132\,
            I => \N__33090\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__33131\,
            I => \N__33086\
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__33130\,
            I => \N__33082\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__33129\,
            I => \N__33078\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__33126\,
            I => \N__33068\
        );

    \I__4374\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33051\
        );

    \I__4373\ : InMux
    port map (
            O => \N__33122\,
            I => \N__33051\
        );

    \I__4372\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33051\
        );

    \I__4371\ : InMux
    port map (
            O => \N__33118\,
            I => \N__33051\
        );

    \I__4370\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33051\
        );

    \I__4369\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33051\
        );

    \I__4368\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33051\
        );

    \I__4367\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33051\
        );

    \I__4366\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33034\
        );

    \I__4365\ : InMux
    port map (
            O => \N__33106\,
            I => \N__33034\
        );

    \I__4364\ : InMux
    port map (
            O => \N__33105\,
            I => \N__33034\
        );

    \I__4363\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33034\
        );

    \I__4362\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33034\
        );

    \I__4361\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33034\
        );

    \I__4360\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33034\
        );

    \I__4359\ : InMux
    port map (
            O => \N__33094\,
            I => \N__33034\
        );

    \I__4358\ : InMux
    port map (
            O => \N__33093\,
            I => \N__33017\
        );

    \I__4357\ : InMux
    port map (
            O => \N__33090\,
            I => \N__33017\
        );

    \I__4356\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33017\
        );

    \I__4355\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33017\
        );

    \I__4354\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33017\
        );

    \I__4353\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33017\
        );

    \I__4352\ : InMux
    port map (
            O => \N__33081\,
            I => \N__33017\
        );

    \I__4351\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33017\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__33077\,
            I => \N__33014\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__33076\,
            I => \N__33011\
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__33075\,
            I => \N__33008\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__33074\,
            I => \N__33005\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__33073\,
            I => \N__33002\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__33072\,
            I => \N__32999\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__33071\,
            I => \N__32996\
        );

    \I__4343\ : Span4Mux_v
    port map (
            O => \N__33068\,
            I => \N__32990\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__32990\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__33034\,
            I => \N__32987\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__33017\,
            I => \N__32984\
        );

    \I__4339\ : InMux
    port map (
            O => \N__33014\,
            I => \N__32975\
        );

    \I__4338\ : InMux
    port map (
            O => \N__33011\,
            I => \N__32975\
        );

    \I__4337\ : InMux
    port map (
            O => \N__33008\,
            I => \N__32975\
        );

    \I__4336\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32975\
        );

    \I__4335\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32966\
        );

    \I__4334\ : InMux
    port map (
            O => \N__32999\,
            I => \N__32966\
        );

    \I__4333\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32966\
        );

    \I__4332\ : InMux
    port map (
            O => \N__32995\,
            I => \N__32966\
        );

    \I__4331\ : Span4Mux_v
    port map (
            O => \N__32990\,
            I => \N__32963\
        );

    \I__4330\ : Span4Mux_h
    port map (
            O => \N__32987\,
            I => \N__32960\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__32984\,
            I => \N__32957\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32952\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__32966\,
            I => \N__32952\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__32963\,
            I => \N__32949\
        );

    \I__4325\ : Span4Mux_v
    port map (
            O => \N__32960\,
            I => \N__32946\
        );

    \I__4324\ : Sp12to4
    port map (
            O => \N__32957\,
            I => \N__32941\
        );

    \I__4323\ : Span12Mux_h
    port map (
            O => \N__32952\,
            I => \N__32941\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__32949\,
            I => \quad_counter1.n2226\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__32946\,
            I => \quad_counter1.n2226\
        );

    \I__4320\ : Odrv12
    port map (
            O => \N__32941\,
            I => \quad_counter1.n2226\
        );

    \I__4319\ : InMux
    port map (
            O => \N__32934\,
            I => \bfn_12_19_0_\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__32931\,
            I => \c0.n24784_cascade_\
        );

    \I__4317\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__32919\,
            I => \N__32916\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__32916\,
            I => n25019
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__32913\,
            I => \N__32909\
        );

    \I__4311\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32906\
        );

    \I__4310\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32903\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__32906\,
            I => data_out_frame_11_2
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__32903\,
            I => data_out_frame_11_2
        );

    \I__4307\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32895\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__32895\,
            I => \N__32892\
        );

    \I__4305\ : Odrv4
    port map (
            O => \N__32892\,
            I => n2273
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__32889\,
            I => \N__32885\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__32888\,
            I => \N__32881\
        );

    \I__4302\ : InMux
    port map (
            O => \N__32885\,
            I => \N__32878\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__32884\,
            I => \N__32874\
        );

    \I__4300\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32871\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__32878\,
            I => \N__32868\
        );

    \I__4298\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32863\
        );

    \I__4297\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32863\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__32871\,
            I => \N__32858\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__32868\,
            I => \N__32858\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__32863\,
            I => encoder1_position_18
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__32858\,
            I => encoder1_position_18
        );

    \I__4292\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32850\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__32850\,
            I => \N__32844\
        );

    \I__4290\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32841\
        );

    \I__4289\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32838\
        );

    \I__4288\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32835\
        );

    \I__4287\ : Sp12to4
    port map (
            O => \N__32844\,
            I => \N__32830\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__32841\,
            I => \N__32830\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__32838\,
            I => \N__32827\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__32835\,
            I => encoder1_position_19
        );

    \I__4283\ : Odrv12
    port map (
            O => \N__32830\,
            I => encoder1_position_19
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__32827\,
            I => encoder1_position_19
        );

    \I__4281\ : InMux
    port map (
            O => \N__32820\,
            I => \N__32817\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__32817\,
            I => \N__32814\
        );

    \I__4279\ : Span4Mux_v
    port map (
            O => \N__32814\,
            I => \N__32811\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__32811\,
            I => n2272
        );

    \I__4277\ : InMux
    port map (
            O => \N__32808\,
            I => \quad_counter1.n19750\
        );

    \I__4276\ : InMux
    port map (
            O => \N__32805\,
            I => \N__32802\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__32802\,
            I => \N__32799\
        );

    \I__4274\ : Odrv12
    port map (
            O => \N__32799\,
            I => n2271
        );

    \I__4273\ : InMux
    port map (
            O => \N__32796\,
            I => \quad_counter1.n19751\
        );

    \I__4272\ : InMux
    port map (
            O => \N__32793\,
            I => \quad_counter1.n19752\
        );

    \I__4271\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32787\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__32787\,
            I => \N__32784\
        );

    \I__4269\ : Span4Mux_h
    port map (
            O => \N__32784\,
            I => \N__32781\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__32781\,
            I => n2269
        );

    \I__4267\ : InMux
    port map (
            O => \N__32778\,
            I => \quad_counter1.n19753\
        );

    \I__4266\ : InMux
    port map (
            O => \N__32775\,
            I => \bfn_12_18_0_\
        );

    \I__4265\ : InMux
    port map (
            O => \N__32772\,
            I => \quad_counter1.n19755\
        );

    \I__4264\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32766\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__32766\,
            I => \N__32763\
        );

    \I__4262\ : Span4Mux_h
    port map (
            O => \N__32763\,
            I => \N__32760\
        );

    \I__4261\ : Span4Mux_v
    port map (
            O => \N__32760\,
            I => \N__32757\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__32757\,
            I => n2266
        );

    \I__4259\ : InMux
    port map (
            O => \N__32754\,
            I => \quad_counter1.n19756\
        );

    \I__4258\ : InMux
    port map (
            O => \N__32751\,
            I => \quad_counter1.n19757\
        );

    \I__4257\ : InMux
    port map (
            O => \N__32748\,
            I => \quad_counter1.n19758\
        );

    \I__4256\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32742\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__32742\,
            I => \N__32739\
        );

    \I__4254\ : Span4Mux_v
    port map (
            O => \N__32739\,
            I => \N__32736\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__32736\,
            I => n2280
        );

    \I__4252\ : InMux
    port map (
            O => \N__32733\,
            I => \quad_counter1.n19742\
        );

    \I__4251\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32727\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32724\
        );

    \I__4249\ : Span4Mux_v
    port map (
            O => \N__32724\,
            I => \N__32721\
        );

    \I__4248\ : Odrv4
    port map (
            O => \N__32721\,
            I => n2279
        );

    \I__4247\ : InMux
    port map (
            O => \N__32718\,
            I => \quad_counter1.n19743\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__32715\,
            I => \N__32712\
        );

    \I__4245\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32708\
        );

    \I__4244\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32703\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32700\
        );

    \I__4242\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32695\
        );

    \I__4241\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32695\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__32703\,
            I => \N__32691\
        );

    \I__4239\ : Span4Mux_v
    port map (
            O => \N__32700\,
            I => \N__32688\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__32695\,
            I => \N__32685\
        );

    \I__4237\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32681\
        );

    \I__4236\ : Span12Mux_h
    port map (
            O => \N__32691\,
            I => \N__32678\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__32688\,
            I => \N__32673\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__32685\,
            I => \N__32673\
        );

    \I__4233\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32670\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__32681\,
            I => encoder1_position_13
        );

    \I__4231\ : Odrv12
    port map (
            O => \N__32678\,
            I => encoder1_position_13
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__32673\,
            I => encoder1_position_13
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__32670\,
            I => encoder1_position_13
        );

    \I__4228\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32658\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32655\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__32655\,
            I => \N__32652\
        );

    \I__4225\ : Span4Mux_v
    port map (
            O => \N__32652\,
            I => \N__32649\
        );

    \I__4224\ : Odrv4
    port map (
            O => \N__32649\,
            I => n2278
        );

    \I__4223\ : InMux
    port map (
            O => \N__32646\,
            I => \quad_counter1.n19744\
        );

    \I__4222\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32640\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__32640\,
            I => \N__32637\
        );

    \I__4220\ : Span4Mux_h
    port map (
            O => \N__32637\,
            I => \N__32634\
        );

    \I__4219\ : Span4Mux_v
    port map (
            O => \N__32634\,
            I => \N__32631\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__32631\,
            I => n2277
        );

    \I__4217\ : InMux
    port map (
            O => \N__32628\,
            I => \quad_counter1.n19745\
        );

    \I__4216\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32622\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__32622\,
            I => n2276
        );

    \I__4214\ : InMux
    port map (
            O => \N__32619\,
            I => \bfn_12_17_0_\
        );

    \I__4213\ : InMux
    port map (
            O => \N__32616\,
            I => \quad_counter1.n19747\
        );

    \I__4212\ : InMux
    port map (
            O => \N__32613\,
            I => \quad_counter1.n19748\
        );

    \I__4211\ : InMux
    port map (
            O => \N__32610\,
            I => \quad_counter1.n19749\
        );

    \I__4210\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32604\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__32604\,
            I => \N__32601\
        );

    \I__4208\ : Odrv4
    port map (
            O => \N__32601\,
            I => n2289
        );

    \I__4207\ : InMux
    port map (
            O => \N__32598\,
            I => \quad_counter1.n19733\
        );

    \I__4206\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32592\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__32592\,
            I => \N__32589\
        );

    \I__4204\ : Sp12to4
    port map (
            O => \N__32589\,
            I => \N__32586\
        );

    \I__4203\ : Odrv12
    port map (
            O => \N__32586\,
            I => n2288
        );

    \I__4202\ : InMux
    port map (
            O => \N__32583\,
            I => \quad_counter1.n19734\
        );

    \I__4201\ : InMux
    port map (
            O => \N__32580\,
            I => \N__32577\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__32577\,
            I => \N__32574\
        );

    \I__4199\ : Odrv12
    port map (
            O => \N__32574\,
            I => n2287
        );

    \I__4198\ : InMux
    port map (
            O => \N__32571\,
            I => \quad_counter1.n19735\
        );

    \I__4197\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32565\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__32565\,
            I => \N__32562\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__32562\,
            I => \N__32559\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__32559\,
            I => \N__32556\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__32556\,
            I => n2286
        );

    \I__4192\ : InMux
    port map (
            O => \N__32553\,
            I => \quad_counter1.n19736\
        );

    \I__4191\ : InMux
    port map (
            O => \N__32550\,
            I => \N__32547\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__32547\,
            I => \N__32544\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__32544\,
            I => \N__32541\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__32541\,
            I => n2285
        );

    \I__4187\ : InMux
    port map (
            O => \N__32538\,
            I => \quad_counter1.n19737\
        );

    \I__4186\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32532\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__32532\,
            I => n2284
        );

    \I__4184\ : InMux
    port map (
            O => \N__32529\,
            I => \bfn_12_16_0_\
        );

    \I__4183\ : InMux
    port map (
            O => \N__32526\,
            I => \quad_counter1.n19739\
        );

    \I__4182\ : InMux
    port map (
            O => \N__32523\,
            I => \N__32520\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__32520\,
            I => \N__32517\
        );

    \I__4180\ : Span4Mux_h
    port map (
            O => \N__32517\,
            I => \N__32514\
        );

    \I__4179\ : Span4Mux_v
    port map (
            O => \N__32514\,
            I => \N__32511\
        );

    \I__4178\ : Odrv4
    port map (
            O => \N__32511\,
            I => n2282
        );

    \I__4177\ : InMux
    port map (
            O => \N__32508\,
            I => \quad_counter1.n19740\
        );

    \I__4176\ : InMux
    port map (
            O => \N__32505\,
            I => \quad_counter1.n19741\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__32502\,
            I => \N__32499\
        );

    \I__4174\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32495\
        );

    \I__4173\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32492\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__32495\,
            I => data_out_frame_7_0
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__32492\,
            I => data_out_frame_7_0
        );

    \I__4170\ : InMux
    port map (
            O => \N__32487\,
            I => \N__32484\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__32484\,
            I => \N__32481\
        );

    \I__4168\ : Span4Mux_v
    port map (
            O => \N__32481\,
            I => \N__32478\
        );

    \I__4167\ : Odrv4
    port map (
            O => \N__32478\,
            I => \c0.n5_adj_4567\
        );

    \I__4166\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32472\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__32472\,
            I => \N__32469\
        );

    \I__4164\ : Span4Mux_v
    port map (
            O => \N__32469\,
            I => \N__32465\
        );

    \I__4163\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32462\
        );

    \I__4162\ : Span4Mux_h
    port map (
            O => \N__32465\,
            I => \N__32459\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__32462\,
            I => data_out_frame_13_1
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__32459\,
            I => data_out_frame_13_1
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__4158\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32448\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32445\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__32445\,
            I => \N__32442\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__32442\,
            I => \N__32439\
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__32439\,
            I => \c0.n11_adj_4646\
        );

    \I__4153\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32433\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__32433\,
            I => \N__32430\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__32430\,
            I => \c0.n5_adj_4644\
        );

    \I__4150\ : InMux
    port map (
            O => \N__32427\,
            I => \N__32424\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__32424\,
            I => \N__32421\
        );

    \I__4148\ : Span4Mux_v
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__32418\,
            I => \c0.n11_adj_4652\
        );

    \I__4146\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32412\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__32412\,
            I => \c0.data_out_frame_28_2\
        );

    \I__4144\ : InMux
    port map (
            O => \N__32409\,
            I => \N__32406\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__32406\,
            I => \N__32403\
        );

    \I__4142\ : Span4Mux_v
    port map (
            O => \N__32403\,
            I => \N__32400\
        );

    \I__4141\ : Span4Mux_v
    port map (
            O => \N__32400\,
            I => \N__32397\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__32397\,
            I => \c0.n26_adj_4651\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__32394\,
            I => \N__32391\
        );

    \I__4138\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32388\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__32388\,
            I => \N__32385\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__32385\,
            I => \quad_counter1.count_direction\
        );

    \I__4135\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32379\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__32379\,
            I => \N__32376\
        );

    \I__4133\ : Span4Mux_h
    port map (
            O => \N__32376\,
            I => \N__32373\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__32373\,
            I => n2291
        );

    \I__4131\ : InMux
    port map (
            O => \N__32370\,
            I => \quad_counter1.n19731\
        );

    \I__4130\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__32364\,
            I => \N__32361\
        );

    \I__4128\ : Span4Mux_v
    port map (
            O => \N__32361\,
            I => \N__32358\
        );

    \I__4127\ : Span4Mux_h
    port map (
            O => \N__32358\,
            I => \N__32355\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__32355\,
            I => n2290
        );

    \I__4125\ : InMux
    port map (
            O => \N__32352\,
            I => \quad_counter1.n19732\
        );

    \I__4124\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32346\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__32346\,
            I => \N__32341\
        );

    \I__4122\ : InMux
    port map (
            O => \N__32345\,
            I => \N__32338\
        );

    \I__4121\ : InMux
    port map (
            O => \N__32344\,
            I => \N__32335\
        );

    \I__4120\ : Span4Mux_h
    port map (
            O => \N__32341\,
            I => \N__32330\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__32338\,
            I => \N__32330\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__32335\,
            I => \N__32327\
        );

    \I__4117\ : Span4Mux_v
    port map (
            O => \N__32330\,
            I => \N__32324\
        );

    \I__4116\ : Odrv12
    port map (
            O => \N__32327\,
            I => \c0.n13531\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__32324\,
            I => \c0.n13531\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__32319\,
            I => \N__32315\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__32318\,
            I => \N__32312\
        );

    \I__4112\ : InMux
    port map (
            O => \N__32315\,
            I => \N__32309\
        );

    \I__4111\ : InMux
    port map (
            O => \N__32312\,
            I => \N__32306\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__32309\,
            I => \c0.n20415\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__32306\,
            I => \c0.n20415\
        );

    \I__4108\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32298\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__32298\,
            I => \N__32294\
        );

    \I__4106\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32291\
        );

    \I__4105\ : Odrv4
    port map (
            O => \N__32294\,
            I => \c0.n22452\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__32291\,
            I => \c0.n22452\
        );

    \I__4103\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32283\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__32283\,
            I => \N__32280\
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__32280\,
            I => \c0.n9_adj_4562\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__32277\,
            I => \c0.n10_adj_4690_cascade_\
        );

    \I__4099\ : InMux
    port map (
            O => \N__32274\,
            I => \N__32271\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__32271\,
            I => \c0.n22710\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__32268\,
            I => \c0.n22710_cascade_\
        );

    \I__4096\ : InMux
    port map (
            O => \N__32265\,
            I => \N__32262\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32256\
        );

    \I__4094\ : InMux
    port map (
            O => \N__32261\,
            I => \N__32253\
        );

    \I__4093\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32248\
        );

    \I__4092\ : InMux
    port map (
            O => \N__32259\,
            I => \N__32248\
        );

    \I__4091\ : Span4Mux_h
    port map (
            O => \N__32256\,
            I => \N__32245\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__32253\,
            I => \N__32240\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__32248\,
            I => \N__32240\
        );

    \I__4088\ : Odrv4
    port map (
            O => \N__32245\,
            I => \c0.n12539\
        );

    \I__4087\ : Odrv12
    port map (
            O => \N__32240\,
            I => \c0.n12539\
        );

    \I__4086\ : InMux
    port map (
            O => \N__32235\,
            I => \N__32227\
        );

    \I__4085\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32227\
        );

    \I__4084\ : InMux
    port map (
            O => \N__32233\,
            I => \N__32224\
        );

    \I__4083\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32221\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__32227\,
            I => \N__32218\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__32224\,
            I => \N__32215\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__32221\,
            I => \c0.n21309\
        );

    \I__4079\ : Odrv12
    port map (
            O => \N__32218\,
            I => \c0.n21309\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__32215\,
            I => \c0.n21309\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__32208\,
            I => \c0.n6_adj_4683_cascade_\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__32205\,
            I => \N__32202\
        );

    \I__4075\ : InMux
    port map (
            O => \N__32202\,
            I => \N__32197\
        );

    \I__4074\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32192\
        );

    \I__4073\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32192\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__32197\,
            I => \N__32189\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__32192\,
            I => \N__32186\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__32189\,
            I => \c0.n13938\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__32186\,
            I => \c0.n13938\
        );

    \I__4068\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32178\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__32178\,
            I => \c0.n12_adj_4688\
        );

    \I__4066\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32172\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__32172\,
            I => \c0.n20360\
        );

    \I__4064\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32163\
        );

    \I__4063\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32163\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__32163\,
            I => \c0.n22668\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__32160\,
            I => \c0.n20360_cascade_\
        );

    \I__4060\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32154\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__32154\,
            I => \c0.data_out_frame_29_7\
        );

    \I__4058\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__32148\,
            I => \N__32145\
        );

    \I__4056\ : Odrv12
    port map (
            O => \N__32145\,
            I => \c0.n26_adj_4713\
        );

    \I__4055\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32131\
        );

    \I__4054\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32131\
        );

    \I__4053\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32131\
        );

    \I__4052\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32128\
        );

    \I__4051\ : InMux
    port map (
            O => \N__32138\,
            I => \N__32125\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__32131\,
            I => \N__32122\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__32128\,
            I => \N__32119\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__32125\,
            I => \c0.n20367\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__32122\,
            I => \c0.n20367\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__32119\,
            I => \c0.n20367\
        );

    \I__4045\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32109\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__32109\,
            I => \N__32106\
        );

    \I__4043\ : Odrv12
    port map (
            O => \N__32106\,
            I => \c0.n6_adj_4336\
        );

    \I__4042\ : InMux
    port map (
            O => \N__32103\,
            I => \N__32100\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__32100\,
            I => \N__32096\
        );

    \I__4040\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32093\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__32096\,
            I => \c0.n22531\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__32093\,
            I => \c0.n22531\
        );

    \I__4037\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32085\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__32085\,
            I => \N__32082\
        );

    \I__4035\ : Span4Mux_v
    port map (
            O => \N__32082\,
            I => \N__32079\
        );

    \I__4034\ : Sp12to4
    port map (
            O => \N__32079\,
            I => \N__32076\
        );

    \I__4033\ : Odrv12
    port map (
            O => \N__32076\,
            I => n25065
        );

    \I__4032\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32070\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__32070\,
            I => \c0.n13741\
        );

    \I__4030\ : CascadeMux
    port map (
            O => \N__32067\,
            I => \c0.n14_adj_4317_cascade_\
        );

    \I__4029\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32061\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__32061\,
            I => \c0.n15_adj_4318\
        );

    \I__4027\ : InMux
    port map (
            O => \N__32058\,
            I => \N__32055\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__32055\,
            I => \c0.n6_adj_4330\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__32052\,
            I => \c0.n21323_cascade_\
        );

    \I__4024\ : InMux
    port map (
            O => \N__32049\,
            I => \N__32046\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__32046\,
            I => \c0.n14_adj_4368\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__32043\,
            I => \c0.n12488_cascade_\
        );

    \I__4021\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__32034\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__32034\,
            I => \c0.n20379\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__32031\,
            I => \c0.n13531_cascade_\
        );

    \I__4017\ : InMux
    port map (
            O => \N__32028\,
            I => \N__32025\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__32025\,
            I => \N__32022\
        );

    \I__4015\ : Span4Mux_v
    port map (
            O => \N__32022\,
            I => \N__32018\
        );

    \I__4014\ : InMux
    port map (
            O => \N__32021\,
            I => \N__32015\
        );

    \I__4013\ : Odrv4
    port map (
            O => \N__32018\,
            I => \c0.n22294\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__32015\,
            I => \c0.n22294\
        );

    \I__4011\ : InMux
    port map (
            O => \N__32010\,
            I => \c0.rx.n19718\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__32007\,
            I => \N__32004\
        );

    \I__4009\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31996\
        );

    \I__4008\ : InMux
    port map (
            O => \N__32003\,
            I => \N__31996\
        );

    \I__4007\ : InMux
    port map (
            O => \N__32002\,
            I => \N__31993\
        );

    \I__4006\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31990\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__31996\,
            I => \N__31987\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__31993\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__31990\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__31987\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__4001\ : InMux
    port map (
            O => \N__31980\,
            I => \c0.rx.n19719\
        );

    \I__4000\ : InMux
    port map (
            O => \N__31977\,
            I => \N__31967\
        );

    \I__3999\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31967\
        );

    \I__3998\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31967\
        );

    \I__3997\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31964\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__31967\,
            I => \N__31961\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__31964\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__31961\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__3993\ : InMux
    port map (
            O => \N__31956\,
            I => \c0.rx.n19720\
        );

    \I__3992\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31950\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__31950\,
            I => \N__31944\
        );

    \I__3990\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31939\
        );

    \I__3989\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31939\
        );

    \I__3988\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31936\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__31944\,
            I => \N__31933\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__31939\,
            I => \N__31930\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__31936\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__31933\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__31930\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__3982\ : InMux
    port map (
            O => \N__31923\,
            I => \c0.rx.n19721\
        );

    \I__3981\ : InMux
    port map (
            O => \N__31920\,
            I => \c0.rx.n19722\
        );

    \I__3980\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31914\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__31914\,
            I => \N__31911\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__31911\,
            I => \N__31908\
        );

    \I__3977\ : Span4Mux_v
    port map (
            O => \N__31908\,
            I => \N__31904\
        );

    \I__3976\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31901\
        );

    \I__3975\ : Sp12to4
    port map (
            O => \N__31904\,
            I => \N__31895\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__31901\,
            I => \N__31891\
        );

    \I__3973\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31888\
        );

    \I__3972\ : InMux
    port map (
            O => \N__31899\,
            I => \N__31885\
        );

    \I__3971\ : InMux
    port map (
            O => \N__31898\,
            I => \N__31882\
        );

    \I__3970\ : Span12Mux_v
    port map (
            O => \N__31895\,
            I => \N__31879\
        );

    \I__3969\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31876\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__31891\,
            I => \N__31871\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__31888\,
            I => \N__31871\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__31885\,
            I => \N__31868\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__31882\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__3964\ : Odrv12
    port map (
            O => \N__31879\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__31876\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__31871\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__31868\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__3960\ : SRMux
    port map (
            O => \N__31857\,
            I => \N__31854\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__31854\,
            I => \N__31851\
        );

    \I__3958\ : Span4Mux_h
    port map (
            O => \N__31851\,
            I => \N__31848\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__31848\,
            I => n14895
        );

    \I__3956\ : SRMux
    port map (
            O => \N__31845\,
            I => \N__31842\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__31842\,
            I => \N__31839\
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__31839\,
            I => \c0.n21645\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__31836\,
            I => \c0.n22638_cascade_\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__31833\,
            I => \n14895_cascade_\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__31830\,
            I => \n24921_cascade_\
        );

    \I__3950\ : InMux
    port map (
            O => \N__31827\,
            I => \N__31824\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__31824\,
            I => \N__31821\
        );

    \I__3948\ : Odrv12
    port map (
            O => \N__31821\,
            I => n24922
        );

    \I__3947\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31815\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__31815\,
            I => \c0.rx.n24916\
        );

    \I__3945\ : InMux
    port map (
            O => \N__31812\,
            I => \N__31809\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__31809\,
            I => \c0.rx.n8\
        );

    \I__3943\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31800\
        );

    \I__3942\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31797\
        );

    \I__3941\ : InMux
    port map (
            O => \N__31804\,
            I => \N__31792\
        );

    \I__3940\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31792\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__31800\,
            I => \r_Clock_Count_0\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__31797\,
            I => \r_Clock_Count_0\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__31792\,
            I => \r_Clock_Count_0\
        );

    \I__3936\ : InMux
    port map (
            O => \N__31785\,
            I => \N__31782\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__31782\,
            I => n226
        );

    \I__3934\ : InMux
    port map (
            O => \N__31779\,
            I => \bfn_11_26_0_\
        );

    \I__3933\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31768\
        );

    \I__3932\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31768\
        );

    \I__3931\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31765\
        );

    \I__3930\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31762\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__31768\,
            I => \N__31759\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__31765\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__31762\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__31759\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__3925\ : InMux
    port map (
            O => \N__31752\,
            I => \c0.rx.n19716\
        );

    \I__3924\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31743\
        );

    \I__3923\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31740\
        );

    \I__3922\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31735\
        );

    \I__3921\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31735\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__31743\,
            I => \N__31732\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__31740\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__31735\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__31732\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__3916\ : InMux
    port map (
            O => \N__31725\,
            I => \c0.rx.n19717\
        );

    \I__3915\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31717\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__31721\,
            I => \N__31714\
        );

    \I__3913\ : InMux
    port map (
            O => \N__31720\,
            I => \N__31710\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__31717\,
            I => \N__31707\
        );

    \I__3911\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31702\
        );

    \I__3910\ : InMux
    port map (
            O => \N__31713\,
            I => \N__31702\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__31710\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__3908\ : Odrv4
    port map (
            O => \N__31707\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__31702\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__31695\,
            I => \c0.rx.n9_cascade_\
        );

    \I__3905\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31688\
        );

    \I__3904\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31684\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__31688\,
            I => \N__31681\
        );

    \I__3902\ : InMux
    port map (
            O => \N__31687\,
            I => \N__31678\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__31684\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__31681\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__31678\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__31671\,
            I => \c0.rx.n17531_cascade_\
        );

    \I__3897\ : InMux
    port map (
            O => \N__31668\,
            I => \N__31665\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__31665\,
            I => \c0.rx.n17590\
        );

    \I__3895\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31659\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__31659\,
            I => \N__31655\
        );

    \I__3893\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31651\
        );

    \I__3892\ : Sp12to4
    port map (
            O => \N__31655\,
            I => \N__31648\
        );

    \I__3891\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31645\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__31651\,
            I => \N__31642\
        );

    \I__3889\ : Span12Mux_v
    port map (
            O => \N__31648\,
            I => \N__31639\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__31645\,
            I => \N__31636\
        );

    \I__3887\ : Span4Mux_h
    port map (
            O => \N__31642\,
            I => \N__31633\
        );

    \I__3886\ : Odrv12
    port map (
            O => \N__31639\,
            I => \c0.rx.n17848\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__31636\,
            I => \c0.rx.n17848\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__31633\,
            I => \c0.rx.n17848\
        );

    \I__3883\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31623\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__31623\,
            I => \c0.rx.n14\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__31620\,
            I => \c0.rx.n24697_cascade_\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__31617\,
            I => \c0.rx.n24914_cascade_\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__31614\,
            I => \N__31611\
        );

    \I__3878\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31608\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__31608\,
            I => \c0.n24255\
        );

    \I__3876\ : SRMux
    port map (
            O => \N__31605\,
            I => \N__31602\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__31602\,
            I => \N__31599\
        );

    \I__3874\ : Sp12to4
    port map (
            O => \N__31599\,
            I => \N__31596\
        );

    \I__3873\ : Odrv12
    port map (
            O => \N__31596\,
            I => \c0.n21583\
        );

    \I__3872\ : InMux
    port map (
            O => \N__31593\,
            I => \N__31589\
        );

    \I__3871\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31586\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__31589\,
            I => \N__31582\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__31586\,
            I => \N__31579\
        );

    \I__3868\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31576\
        );

    \I__3867\ : Span4Mux_h
    port map (
            O => \N__31582\,
            I => \N__31573\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__31579\,
            I => \N__31570\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__31576\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__31573\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__31570\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__3862\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31560\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__31560\,
            I => \N__31555\
        );

    \I__3860\ : InMux
    port map (
            O => \N__31559\,
            I => \N__31552\
        );

    \I__3859\ : InMux
    port map (
            O => \N__31558\,
            I => \N__31549\
        );

    \I__3858\ : Span4Mux_h
    port map (
            O => \N__31555\,
            I => \N__31546\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__31552\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__31549\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__31546\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__31539\,
            I => \c0.n14530_cascade_\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__31536\,
            I => \N__31533\
        );

    \I__3852\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31529\
        );

    \I__3851\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31526\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31523\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__31526\,
            I => data_out_frame_11_6
        );

    \I__3848\ : Odrv12
    port map (
            O => \N__31523\,
            I => data_out_frame_11_6
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__31518\,
            I => \c0.n25098_cascade_\
        );

    \I__3846\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__31512\,
            I => \c0.n25101\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__31509\,
            I => \N__31506\
        );

    \I__3843\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31500\
        );

    \I__3842\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31500\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__31500\,
            I => data_out_frame_6_5
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__31497\,
            I => \N__31494\
        );

    \I__3839\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31490\
        );

    \I__3838\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31487\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__31490\,
            I => data_out_frame_5_5
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__31487\,
            I => data_out_frame_5_5
        );

    \I__3835\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31479\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__31479\,
            I => \c0.n5_adj_4679\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__31476\,
            I => \c0.n25016_cascade_\
        );

    \I__3832\ : InMux
    port map (
            O => \N__31473\,
            I => \N__31470\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__31470\,
            I => \N__31467\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__31467\,
            I => \c0.n24794\
        );

    \I__3829\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31461\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__31461\,
            I => \c0.n5_adj_4700\
        );

    \I__3827\ : InMux
    port map (
            O => \N__31458\,
            I => \N__31454\
        );

    \I__3826\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31451\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__31454\,
            I => data_out_frame_10_2
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__31451\,
            I => data_out_frame_10_2
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__31446\,
            I => \N__31442\
        );

    \I__3822\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31437\
        );

    \I__3821\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31437\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__31437\,
            I => data_out_frame_11_0
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__31434\,
            I => \N__31431\
        );

    \I__3818\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31428\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__31428\,
            I => \N__31425\
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__31425\,
            I => \c0.n11_adj_4703\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__31422\,
            I => \c0.n24945_cascade_\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__31419\,
            I => \N__31412\
        );

    \I__3813\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31409\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__31417\,
            I => \N__31406\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__31416\,
            I => \N__31402\
        );

    \I__3810\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31396\
        );

    \I__3809\ : InMux
    port map (
            O => \N__31412\,
            I => \N__31396\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__31409\,
            I => \N__31392\
        );

    \I__3807\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31389\
        );

    \I__3806\ : InMux
    port map (
            O => \N__31405\,
            I => \N__31386\
        );

    \I__3805\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31381\
        );

    \I__3804\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31381\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__31396\,
            I => \N__31378\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__31395\,
            I => \N__31375\
        );

    \I__3801\ : Span4Mux_v
    port map (
            O => \N__31392\,
            I => \N__31372\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__31389\,
            I => \N__31369\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31366\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__31381\,
            I => \N__31363\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__31378\,
            I => \N__31360\
        );

    \I__3796\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31357\
        );

    \I__3795\ : Span4Mux_h
    port map (
            O => \N__31372\,
            I => \N__31352\
        );

    \I__3794\ : Span4Mux_v
    port map (
            O => \N__31369\,
            I => \N__31352\
        );

    \I__3793\ : Span4Mux_v
    port map (
            O => \N__31366\,
            I => \N__31347\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__31363\,
            I => \N__31347\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__31360\,
            I => \N__31344\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__31357\,
            I => \N__31341\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__31352\,
            I => n24682
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__31347\,
            I => n24682
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__31344\,
            I => n24682
        );

    \I__3786\ : Odrv12
    port map (
            O => \N__31341\,
            I => n24682
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__31332\,
            I => \c0.n24797_cascade_\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__31329\,
            I => \N__31325\
        );

    \I__3783\ : InMux
    port map (
            O => \N__31328\,
            I => \N__31320\
        );

    \I__3782\ : InMux
    port map (
            O => \N__31325\,
            I => \N__31305\
        );

    \I__3781\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31305\
        );

    \I__3780\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31305\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__31320\,
            I => \N__31300\
        );

    \I__3778\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31297\
        );

    \I__3777\ : CascadeMux
    port map (
            O => \N__31318\,
            I => \N__31294\
        );

    \I__3776\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31291\
        );

    \I__3775\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31286\
        );

    \I__3774\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31286\
        );

    \I__3773\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31281\
        );

    \I__3772\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31281\
        );

    \I__3771\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31278\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__31305\,
            I => \N__31275\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__31304\,
            I => \N__31272\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__31303\,
            I => \N__31267\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__31300\,
            I => \N__31261\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31261\
        );

    \I__3765\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31258\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31255\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__31286\,
            I => \N__31248\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31248\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__31278\,
            I => \N__31248\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__31275\,
            I => \N__31245\
        );

    \I__3759\ : InMux
    port map (
            O => \N__31272\,
            I => \N__31242\
        );

    \I__3758\ : InMux
    port map (
            O => \N__31271\,
            I => \N__31237\
        );

    \I__3757\ : InMux
    port map (
            O => \N__31270\,
            I => \N__31237\
        );

    \I__3756\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31234\
        );

    \I__3755\ : InMux
    port map (
            O => \N__31266\,
            I => \N__31231\
        );

    \I__3754\ : Span4Mux_v
    port map (
            O => \N__31261\,
            I => \N__31226\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__31258\,
            I => \N__31226\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__31255\,
            I => \N__31219\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__31248\,
            I => \N__31219\
        );

    \I__3750\ : Span4Mux_v
    port map (
            O => \N__31245\,
            I => \N__31219\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__31242\,
            I => \N__31214\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__31237\,
            I => \N__31214\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__31234\,
            I => \N__31211\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__31231\,
            I => byte_transmit_counter_4
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__31226\,
            I => byte_transmit_counter_4
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__31219\,
            I => byte_transmit_counter_4
        );

    \I__3743\ : Odrv12
    port map (
            O => \N__31214\,
            I => byte_transmit_counter_4
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__31211\,
            I => byte_transmit_counter_4
        );

    \I__3741\ : InMux
    port map (
            O => \N__31200\,
            I => \N__31194\
        );

    \I__3740\ : InMux
    port map (
            O => \N__31199\,
            I => \N__31191\
        );

    \I__3739\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31186\
        );

    \I__3738\ : InMux
    port map (
            O => \N__31197\,
            I => \N__31183\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31178\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__31191\,
            I => \N__31178\
        );

    \I__3735\ : InMux
    port map (
            O => \N__31190\,
            I => \N__31173\
        );

    \I__3734\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31170\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__31186\,
            I => \N__31167\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31162\
        );

    \I__3731\ : Span4Mux_h
    port map (
            O => \N__31178\,
            I => \N__31162\
        );

    \I__3730\ : InMux
    port map (
            O => \N__31177\,
            I => \N__31159\
        );

    \I__3729\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31153\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__31173\,
            I => \N__31150\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__31170\,
            I => \N__31147\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__31167\,
            I => \N__31140\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__31162\,
            I => \N__31140\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__31159\,
            I => \N__31140\
        );

    \I__3723\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31137\
        );

    \I__3722\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31134\
        );

    \I__3721\ : InMux
    port map (
            O => \N__31156\,
            I => \N__31131\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__31153\,
            I => \N__31128\
        );

    \I__3719\ : Span4Mux_h
    port map (
            O => \N__31150\,
            I => \N__31125\
        );

    \I__3718\ : Span4Mux_v
    port map (
            O => \N__31147\,
            I => \N__31120\
        );

    \I__3717\ : Span4Mux_v
    port map (
            O => \N__31140\,
            I => \N__31120\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__31137\,
            I => \N__31115\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31115\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__31131\,
            I => byte_transmit_counter_3
        );

    \I__3713\ : Odrv12
    port map (
            O => \N__31128\,
            I => byte_transmit_counter_3
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__31125\,
            I => byte_transmit_counter_3
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__31120\,
            I => byte_transmit_counter_3
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__31115\,
            I => byte_transmit_counter_3
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__31104\,
            I => \n24799_cascade_\
        );

    \I__3708\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31098\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__31098\,
            I => n25012
        );

    \I__3706\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31092\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__31092\,
            I => \N__31089\
        );

    \I__3704\ : Span4Mux_h
    port map (
            O => \N__31089\,
            I => \N__31086\
        );

    \I__3703\ : Odrv4
    port map (
            O => \N__31086\,
            I => n10_adj_4775
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__3701\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31077\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__31077\,
            I => \N__31074\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__31074\,
            I => \c0.n24953\
        );

    \I__3698\ : InMux
    port map (
            O => \N__31071\,
            I => \N__31068\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__3696\ : Span4Mux_h
    port map (
            O => \N__31065\,
            I => \N__31062\
        );

    \I__3695\ : Odrv4
    port map (
            O => \N__31062\,
            I => \c0.n24803\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__31059\,
            I => \N__31055\
        );

    \I__3693\ : InMux
    port map (
            O => \N__31058\,
            I => \N__31052\
        );

    \I__3692\ : InMux
    port map (
            O => \N__31055\,
            I => \N__31049\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__31052\,
            I => data_out_frame_8_2
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__31049\,
            I => data_out_frame_8_2
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__31044\,
            I => \c0.n25059_cascade_\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__31041\,
            I => \n25004_cascade_\
        );

    \I__3687\ : InMux
    port map (
            O => \N__31038\,
            I => \N__31035\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__31035\,
            I => \N__31032\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__31032\,
            I => n10_adj_4778
        );

    \I__3684\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__31026\,
            I => \c0.n24809\
        );

    \I__3682\ : InMux
    port map (
            O => \N__31023\,
            I => \N__31020\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__31020\,
            I => n24811
        );

    \I__3680\ : InMux
    port map (
            O => \N__31017\,
            I => \N__31014\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__31014\,
            I => \N__31011\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__31011\,
            I => \N__31008\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__31008\,
            I => n24904
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__31005\,
            I => \N__31001\
        );

    \I__3675\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30998\
        );

    \I__3674\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30995\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__30998\,
            I => \N__30992\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__30995\,
            I => \N__30989\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__30992\,
            I => \N__30986\
        );

    \I__3670\ : Odrv12
    port map (
            O => \N__30989\,
            I => data_out_frame_28_3
        );

    \I__3669\ : Odrv4
    port map (
            O => \N__30986\,
            I => data_out_frame_28_3
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__30981\,
            I => \c0.n25110_cascade_\
        );

    \I__3667\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__30975\,
            I => \c0.n25113\
        );

    \I__3665\ : InMux
    port map (
            O => \N__30972\,
            I => \N__30969\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__30969\,
            I => \c0.n25056\
        );

    \I__3663\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30963\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__30963\,
            I => \N__30959\
        );

    \I__3661\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30956\
        );

    \I__3660\ : Span12Mux_s10_h
    port map (
            O => \N__30959\,
            I => \N__30953\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__30956\,
            I => data_out_frame_10_3
        );

    \I__3658\ : Odrv12
    port map (
            O => \N__30953\,
            I => data_out_frame_10_3
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__30948\,
            I => \N__30945\
        );

    \I__3656\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30942\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__30942\,
            I => \N__30938\
        );

    \I__3654\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30935\
        );

    \I__3653\ : Span4Mux_v
    port map (
            O => \N__30938\,
            I => \N__30932\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__30935\,
            I => \c0.n21362\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__30932\,
            I => \c0.n21362\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__30927\,
            I => \N__30924\
        );

    \I__3649\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30921\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__30921\,
            I => \N__30918\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__30918\,
            I => \c0.n11_adj_4572\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__30915\,
            I => \N__30912\
        );

    \I__3645\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30906\
        );

    \I__3644\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30906\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__30906\,
            I => data_out_frame_13_0
        );

    \I__3642\ : InMux
    port map (
            O => \N__30903\,
            I => \N__30899\
        );

    \I__3641\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30896\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__30899\,
            I => \N__30893\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__30896\,
            I => data_out_frame_6_2
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__30893\,
            I => data_out_frame_6_2
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__30888\,
            I => \c0.n5_adj_4650_cascade_\
        );

    \I__3636\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30882\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__30882\,
            I => \N__30879\
        );

    \I__3634\ : Odrv12
    port map (
            O => \N__30879\,
            I => \c0.n6_adj_4649\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__30876\,
            I => \n22735_cascade_\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__30873\,
            I => \N__30870\
        );

    \I__3631\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30867\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__30867\,
            I => \c0.n22757\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__30864\,
            I => \c0.n20_adj_4699_cascade_\
        );

    \I__3628\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__30858\,
            I => n22285
        );

    \I__3626\ : InMux
    port map (
            O => \N__30855\,
            I => \N__30852\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__30852\,
            I => \N__30849\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__30849\,
            I => \c0.n6_adj_4210\
        );

    \I__3623\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30839\
        );

    \I__3622\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30839\
        );

    \I__3621\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30836\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__30839\,
            I => \c0.n13683\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__30836\,
            I => \c0.n13683\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__30831\,
            I => \c0.n22534_cascade_\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__30828\,
            I => \c0.n20415_cascade_\
        );

    \I__3616\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30820\
        );

    \I__3615\ : InMux
    port map (
            O => \N__30824\,
            I => \N__30815\
        );

    \I__3614\ : InMux
    port map (
            O => \N__30823\,
            I => \N__30815\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__30820\,
            I => \c0.n20384\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__30815\,
            I => \c0.n20384\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__30810\,
            I => \N__30806\
        );

    \I__3610\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30803\
        );

    \I__3609\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30800\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__30803\,
            I => \c0.n22544\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__30800\,
            I => \c0.n22544\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__30795\,
            I => \N__30792\
        );

    \I__3605\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30789\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__30789\,
            I => \c0.data_out_frame_28_5\
        );

    \I__3603\ : InMux
    port map (
            O => \N__30786\,
            I => \N__30783\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__30783\,
            I => \N__30780\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__30780\,
            I => \N__30777\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__30777\,
            I => \c0.n26_adj_4680\
        );

    \I__3599\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30767\
        );

    \I__3598\ : InMux
    port map (
            O => \N__30773\,
            I => \N__30767\
        );

    \I__3597\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30764\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__30767\,
            I => \c0.n22478\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__30764\,
            I => \c0.n22478\
        );

    \I__3594\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30756\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__30756\,
            I => n22735
        );

    \I__3592\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30750\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__30750\,
            I => \c0.n6_adj_4456\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__30747\,
            I => \n21484_cascade_\
        );

    \I__3589\ : InMux
    port map (
            O => \N__30744\,
            I => \N__30740\
        );

    \I__3588\ : InMux
    port map (
            O => \N__30743\,
            I => \N__30737\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__30740\,
            I => \c0.n22246\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__30737\,
            I => \c0.n22246\
        );

    \I__3585\ : InMux
    port map (
            O => \N__30732\,
            I => \N__30728\
        );

    \I__3584\ : InMux
    port map (
            O => \N__30731\,
            I => \N__30725\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__30728\,
            I => \N__30722\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__30725\,
            I => data_out_frame_7_3
        );

    \I__3581\ : Odrv4
    port map (
            O => \N__30722\,
            I => data_out_frame_7_3
        );

    \I__3580\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30714\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__30714\,
            I => \c0.n10_adj_4313\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__30711\,
            I => \N__30708\
        );

    \I__3577\ : InMux
    port map (
            O => \N__30708\,
            I => \N__30705\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__30705\,
            I => \N__30701\
        );

    \I__3575\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30698\
        );

    \I__3574\ : Span4Mux_v
    port map (
            O => \N__30701\,
            I => \N__30695\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__30698\,
            I => data_out_frame_11_3
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__30695\,
            I => data_out_frame_11_3
        );

    \I__3571\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30687\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__30687\,
            I => \c0.n22534\
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__30684\,
            I => \c0.n22246_cascade_\
        );

    \I__3568\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30677\
        );

    \I__3567\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30674\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__30677\,
            I => \N__30671\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__30674\,
            I => \c0.n22846\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__30671\,
            I => \c0.n22846\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__30666\,
            I => \c0.n20379_cascade_\
        );

    \I__3562\ : InMux
    port map (
            O => \N__30663\,
            I => \N__30660\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__30660\,
            I => \N__30653\
        );

    \I__3560\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30646\
        );

    \I__3559\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30646\
        );

    \I__3558\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30646\
        );

    \I__3557\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30643\
        );

    \I__3556\ : Span4Mux_v
    port map (
            O => \N__30653\,
            I => \N__30640\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__30646\,
            I => \N__30637\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__30643\,
            I => \A_filtered_adj_4763\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__30640\,
            I => \A_filtered_adj_4763\
        );

    \I__3552\ : Odrv12
    port map (
            O => \N__30637\,
            I => \A_filtered_adj_4763\
        );

    \I__3551\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30627\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__30627\,
            I => \N__30624\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__30624\,
            I => \N__30619\
        );

    \I__3548\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30614\
        );

    \I__3547\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30614\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__30619\,
            I => \quad_counter1.B_delayed\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__30614\,
            I => \quad_counter1.B_delayed\
        );

    \I__3544\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30603\
        );

    \I__3543\ : InMux
    port map (
            O => \N__30608\,
            I => \N__30603\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__30603\,
            I => \c0.data_out_frame_29__7__N_849\
        );

    \I__3541\ : SRMux
    port map (
            O => \N__30600\,
            I => \N__30597\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__30597\,
            I => \c0.n21597\
        );

    \I__3539\ : SRMux
    port map (
            O => \N__30594\,
            I => \N__30591\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__30591\,
            I => \N__30588\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__30588\,
            I => \c0.n21587\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__30585\,
            I => \c0.n10_adj_4303_cascade_\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__30582\,
            I => \N__30578\
        );

    \I__3534\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30574\
        );

    \I__3533\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30569\
        );

    \I__3532\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30569\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__30574\,
            I => \N__30566\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__30569\,
            I => \N__30562\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__30566\,
            I => \N__30559\
        );

    \I__3528\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30556\
        );

    \I__3527\ : Span12Mux_v
    port map (
            O => \N__30562\,
            I => \N__30551\
        );

    \I__3526\ : Span4Mux_v
    port map (
            O => \N__30559\,
            I => \N__30548\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__30556\,
            I => \N__30545\
        );

    \I__3524\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30542\
        );

    \I__3523\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30539\
        );

    \I__3522\ : Odrv12
    port map (
            O => \N__30551\,
            I => \c0.r_SM_Main_2_N_3754_0\
        );

    \I__3521\ : Odrv4
    port map (
            O => \N__30548\,
            I => \c0.r_SM_Main_2_N_3754_0\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__30545\,
            I => \c0.r_SM_Main_2_N_3754_0\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__30542\,
            I => \c0.r_SM_Main_2_N_3754_0\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__30539\,
            I => \c0.r_SM_Main_2_N_3754_0\
        );

    \I__3517\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30521\
        );

    \I__3516\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30521\
        );

    \I__3515\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30517\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30514\
        );

    \I__3513\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30511\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__30517\,
            I => \N__30508\
        );

    \I__3511\ : Span4Mux_v
    port map (
            O => \N__30514\,
            I => \N__30505\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__30511\,
            I => \c0.tx_active\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__30508\,
            I => \c0.tx_active\
        );

    \I__3508\ : Odrv4
    port map (
            O => \N__30505\,
            I => \c0.tx_active\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__30498\,
            I => \c0.n5_cascade_\
        );

    \I__3506\ : SRMux
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__3504\ : Span4Mux_h
    port map (
            O => \N__30489\,
            I => \N__30486\
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__30486\,
            I => \c0.n21585\
        );

    \I__3502\ : InMux
    port map (
            O => \N__30483\,
            I => \N__30480\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__30480\,
            I => \c0.n3\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__30477\,
            I => \c0.n8_adj_4740_cascade_\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__30474\,
            I => \c0.n22952_cascade_\
        );

    \I__3498\ : CEMux
    port map (
            O => \N__30471\,
            I => \N__30468\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__30468\,
            I => \c0.n14380\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__30465\,
            I => \c0.n14380_cascade_\
        );

    \I__3495\ : SRMux
    port map (
            O => \N__30462\,
            I => \N__30459\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__30459\,
            I => \c0.n14942\
        );

    \I__3493\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30453\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__30453\,
            I => \c0.n4728\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__30450\,
            I => \c0.n4728_cascade_\
        );

    \I__3490\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30444\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__30444\,
            I => \c0.n58_adj_4742\
        );

    \I__3488\ : SRMux
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30434\
        );

    \I__3486\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30431\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__30434\,
            I => \c0.n22952\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__30431\,
            I => \c0.n22952\
        );

    \I__3483\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30423\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__30423\,
            I => n25008
        );

    \I__3481\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30417\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__30417\,
            I => \c0.n11_adj_4681\
        );

    \I__3479\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30411\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30408\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__30408\,
            I => \c0.n24897\
        );

    \I__3476\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30399\
        );

    \I__3475\ : InMux
    port map (
            O => \N__30404\,
            I => \N__30399\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__30399\,
            I => data_out_frame_5_0
        );

    \I__3473\ : InMux
    port map (
            O => \N__30396\,
            I => \N__30390\
        );

    \I__3472\ : InMux
    port map (
            O => \N__30395\,
            I => \N__30390\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__30390\,
            I => data_out_frame_0_2
        );

    \I__3470\ : InMux
    port map (
            O => \N__30387\,
            I => \N__30383\
        );

    \I__3469\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30380\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__30383\,
            I => \N__30377\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__30380\,
            I => data_out_frame_12_5
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__30377\,
            I => data_out_frame_12_5
        );

    \I__3465\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30369\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__30369\,
            I => \N__30366\
        );

    \I__3463\ : Odrv12
    port map (
            O => \N__30366\,
            I => \c0.n24900\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__30363\,
            I => \n14247_cascade_\
        );

    \I__3461\ : InMux
    port map (
            O => \N__30360\,
            I => \N__30354\
        );

    \I__3460\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30354\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__30354\,
            I => data_out_frame_0_3
        );

    \I__3458\ : InMux
    port map (
            O => \N__30351\,
            I => \N__30348\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__30345\,
            I => \N__30342\
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__30342\,
            I => n24796
        );

    \I__3454\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30336\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__30336\,
            I => \N__30332\
        );

    \I__3452\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30329\
        );

    \I__3451\ : Span4Mux_h
    port map (
            O => \N__30332\,
            I => \N__30326\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__30329\,
            I => data_out_frame_7_7
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__30326\,
            I => data_out_frame_7_7
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__30321\,
            I => \n24805_cascade_\
        );

    \I__3447\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__30315\,
            I => n10_adj_4780
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__30312\,
            I => \N__30309\
        );

    \I__3444\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30305\
        );

    \I__3443\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30302\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__30305\,
            I => \N__30299\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__30302\,
            I => data_out_frame_11_5
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__30299\,
            I => data_out_frame_11_5
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__30294\,
            I => \c0.n25092_cascade_\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__30291\,
            I => \c0.n25095_cascade_\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__30288\,
            I => \N__30285\
        );

    \I__3436\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30282\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__30282\,
            I => \N__30279\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__30279\,
            I => \N__30276\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__30276\,
            I => n25014
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__30273\,
            I => \N__30270\
        );

    \I__3431\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30264\
        );

    \I__3430\ : InMux
    port map (
            O => \N__30269\,
            I => \N__30264\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__30264\,
            I => data_out_frame_9_5
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__30261\,
            I => \c0.n20341_cascade_\
        );

    \I__3427\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30255\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__30255\,
            I => \N__30251\
        );

    \I__3425\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30248\
        );

    \I__3424\ : Span4Mux_v
    port map (
            O => \N__30251\,
            I => \N__30245\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__30248\,
            I => data_out_frame_13_7
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__30245\,
            I => data_out_frame_13_7
        );

    \I__3421\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30237\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__30237\,
            I => \N__30233\
        );

    \I__3419\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30230\
        );

    \I__3418\ : Span4Mux_v
    port map (
            O => \N__30233\,
            I => \N__30227\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__30230\,
            I => data_out_frame_10_7
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__30227\,
            I => data_out_frame_10_7
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__30222\,
            I => \N__30218\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__30221\,
            I => \N__30214\
        );

    \I__3413\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30210\
        );

    \I__3412\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30207\
        );

    \I__3411\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30204\
        );

    \I__3410\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30198\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__30210\,
            I => \N__30195\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__30207\,
            I => \N__30192\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__30204\,
            I => \N__30189\
        );

    \I__3406\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30184\
        );

    \I__3405\ : InMux
    port map (
            O => \N__30202\,
            I => \N__30184\
        );

    \I__3404\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30181\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__30198\,
            I => \N__30178\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__30195\,
            I => \N__30175\
        );

    \I__3401\ : Span4Mux_v
    port map (
            O => \N__30192\,
            I => \N__30168\
        );

    \I__3400\ : Span4Mux_h
    port map (
            O => \N__30189\,
            I => \N__30168\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__30184\,
            I => \N__30168\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__30181\,
            I => \N__30165\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__30178\,
            I => \N__30162\
        );

    \I__3396\ : Span4Mux_v
    port map (
            O => \N__30175\,
            I => \N__30159\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__30168\,
            I => \N__30156\
        );

    \I__3394\ : Odrv12
    port map (
            O => \N__30165\,
            I => n9603
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__30162\,
            I => n9603
        );

    \I__3392\ : Odrv4
    port map (
            O => \N__30159\,
            I => n9603
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__30156\,
            I => n9603
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__30147\,
            I => \N__30143\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__30146\,
            I => \N__30140\
        );

    \I__3388\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30135\
        );

    \I__3387\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30132\
        );

    \I__3386\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30126\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__30138\,
            I => \N__30122\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__30135\,
            I => \N__30119\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__30132\,
            I => \N__30116\
        );

    \I__3382\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30113\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__30130\,
            I => \N__30110\
        );

    \I__3380\ : InMux
    port map (
            O => \N__30129\,
            I => \N__30107\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__30126\,
            I => \N__30104\
        );

    \I__3378\ : InMux
    port map (
            O => \N__30125\,
            I => \N__30099\
        );

    \I__3377\ : InMux
    port map (
            O => \N__30122\,
            I => \N__30099\
        );

    \I__3376\ : Span4Mux_h
    port map (
            O => \N__30119\,
            I => \N__30096\
        );

    \I__3375\ : Span4Mux_v
    port map (
            O => \N__30116\,
            I => \N__30091\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__30113\,
            I => \N__30091\
        );

    \I__3373\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30087\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__30107\,
            I => \N__30084\
        );

    \I__3371\ : Span4Mux_h
    port map (
            O => \N__30104\,
            I => \N__30081\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__30099\,
            I => \N__30078\
        );

    \I__3369\ : Sp12to4
    port map (
            O => \N__30096\,
            I => \N__30073\
        );

    \I__3368\ : Sp12to4
    port map (
            O => \N__30091\,
            I => \N__30073\
        );

    \I__3367\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30069\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__30087\,
            I => \N__30064\
        );

    \I__3365\ : Span4Mux_h
    port map (
            O => \N__30084\,
            I => \N__30064\
        );

    \I__3364\ : Span4Mux_v
    port map (
            O => \N__30081\,
            I => \N__30061\
        );

    \I__3363\ : Span12Mux_v
    port map (
            O => \N__30078\,
            I => \N__30058\
        );

    \I__3362\ : Span12Mux_v
    port map (
            O => \N__30073\,
            I => \N__30055\
        );

    \I__3361\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30052\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__30069\,
            I => byte_transmit_counter_5
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__30064\,
            I => byte_transmit_counter_5
        );

    \I__3358\ : Odrv4
    port map (
            O => \N__30061\,
            I => byte_transmit_counter_5
        );

    \I__3357\ : Odrv12
    port map (
            O => \N__30058\,
            I => byte_transmit_counter_5
        );

    \I__3356\ : Odrv12
    port map (
            O => \N__30055\,
            I => byte_transmit_counter_5
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__30052\,
            I => byte_transmit_counter_5
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__30039\,
            I => \N__30036\
        );

    \I__3353\ : InMux
    port map (
            O => \N__30036\,
            I => \N__30033\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__30033\,
            I => \N__30029\
        );

    \I__3351\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30026\
        );

    \I__3350\ : Span4Mux_h
    port map (
            O => \N__30029\,
            I => \N__30023\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__30026\,
            I => \r_Tx_Data_0\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__30023\,
            I => \r_Tx_Data_0\
        );

    \I__3347\ : InMux
    port map (
            O => \N__30018\,
            I => \N__30014\
        );

    \I__3346\ : InMux
    port map (
            O => \N__30017\,
            I => \N__30011\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__30014\,
            I => \N__30008\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__30011\,
            I => data_out_frame_13_6
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__30008\,
            I => data_out_frame_13_6
        );

    \I__3342\ : InMux
    port map (
            O => \N__30003\,
            I => \N__30000\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__30000\,
            I => \N__29996\
        );

    \I__3340\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29993\
        );

    \I__3339\ : Span4Mux_h
    port map (
            O => \N__29996\,
            I => \N__29990\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__29993\,
            I => data_out_frame_8_3
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__29990\,
            I => data_out_frame_8_3
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__29985\,
            I => \c0.n24033_cascade_\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__29982\,
            I => \n21307_cascade_\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__29979\,
            I => \c0.n7_cascade_\
        );

    \I__3333\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__29973\,
            I => \c0.n23918\
        );

    \I__3331\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29967\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__29967\,
            I => \N__29963\
        );

    \I__3329\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29960\
        );

    \I__3328\ : Span4Mux_v
    port map (
            O => \N__29963\,
            I => \N__29957\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__29960\,
            I => \r_Tx_Data_2\
        );

    \I__3326\ : Odrv4
    port map (
            O => \N__29957\,
            I => \r_Tx_Data_2\
        );

    \I__3325\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29949\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__29949\,
            I => \c0.n22163\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__29946\,
            I => \c0.n6_adj_4297_cascade_\
        );

    \I__3322\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29940\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__29940\,
            I => \c0.data_out_frame_28_4\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__29937\,
            I => \n26_cascade_\
        );

    \I__3319\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29931\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29928\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__29928\,
            I => n25021
        );

    \I__3316\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29922\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__29922\,
            I => \N__29919\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__29919\,
            I => n25022
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__29916\,
            I => \c0.n21391_cascade_\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__29913\,
            I => \c0.n21362_cascade_\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__29910\,
            I => \c0.n21244_cascade_\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__29907\,
            I => \N__29903\
        );

    \I__3309\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29900\
        );

    \I__3308\ : InMux
    port map (
            O => \N__29903\,
            I => \N__29897\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__29900\,
            I => \N__29892\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__29897\,
            I => \N__29892\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__29892\,
            I => \N__29888\
        );

    \I__3304\ : InMux
    port map (
            O => \N__29891\,
            I => \N__29885\
        );

    \I__3303\ : Span4Mux_h
    port map (
            O => \N__29888\,
            I => \N__29882\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__29885\,
            I => \B_filtered_adj_4764\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__29882\,
            I => \B_filtered_adj_4764\
        );

    \I__3300\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29874\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__29874\,
            I => \quad_counter1.A_delayed\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__29871\,
            I => \N__29867\
        );

    \I__3297\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29864\
        );

    \I__3296\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29861\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__29864\,
            I => \r_Tx_Data_4\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__29861\,
            I => \r_Tx_Data_4\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__29856\,
            I => \n9806_cascade_\
        );

    \I__3292\ : InMux
    port map (
            O => \N__29853\,
            I => \N__29847\
        );

    \I__3291\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29847\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__29847\,
            I => \N__29842\
        );

    \I__3289\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29837\
        );

    \I__3288\ : InMux
    port map (
            O => \N__29845\,
            I => \N__29837\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__29842\,
            I => \N__29834\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__29837\,
            I => \N__29831\
        );

    \I__3285\ : Span4Mux_h
    port map (
            O => \N__29834\,
            I => \N__29828\
        );

    \I__3284\ : Span12Mux_h
    port map (
            O => \N__29831\,
            I => \N__29825\
        );

    \I__3283\ : Span4Mux_v
    port map (
            O => \N__29828\,
            I => \N__29822\
        );

    \I__3282\ : Odrv12
    port map (
            O => \N__29825\,
            I => \PIN_12_c\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__29822\,
            I => \PIN_12_c\
        );

    \I__3280\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29810\
        );

    \I__3279\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29810\
        );

    \I__3278\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29807\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__29810\,
            I => \quadA_delayed_adj_4767\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__29807\,
            I => \quadA_delayed_adj_4767\
        );

    \I__3275\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29799\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__29799\,
            I => n9806
        );

    \I__3273\ : CEMux
    port map (
            O => \N__29796\,
            I => \N__29793\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__29790\,
            I => \N__29786\
        );

    \I__3270\ : CEMux
    port map (
            O => \N__29789\,
            I => \N__29783\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__29786\,
            I => n14345
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__29783\,
            I => n14345
        );

    \I__3267\ : SRMux
    port map (
            O => \N__29778\,
            I => \N__29774\
        );

    \I__3266\ : SRMux
    port map (
            O => \N__29777\,
            I => \N__29771\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__29774\,
            I => \N__29767\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__29771\,
            I => \N__29764\
        );

    \I__3263\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29761\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__29767\,
            I => \N__29758\
        );

    \I__3261\ : Span4Mux_h
    port map (
            O => \N__29764\,
            I => \N__29755\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__29761\,
            I => \a_delay_counter_15__N_4123_adj_4772\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__29758\,
            I => \a_delay_counter_15__N_4123_adj_4772\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__29755\,
            I => \a_delay_counter_15__N_4123_adj_4772\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__29748\,
            I => \n14345_cascade_\
        );

    \I__3256\ : InMux
    port map (
            O => \N__29745\,
            I => \N__29742\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__29742\,
            I => n39_adj_4770
        );

    \I__3254\ : InMux
    port map (
            O => \N__29739\,
            I => \N__29735\
        );

    \I__3253\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29732\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__29735\,
            I => \quad_counter1.a_delay_counter_5\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__29732\,
            I => \quad_counter1.a_delay_counter_5\
        );

    \I__3250\ : InMux
    port map (
            O => \N__29727\,
            I => \N__29723\
        );

    \I__3249\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29720\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__29723\,
            I => \quad_counter1.a_delay_counter_11\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__29720\,
            I => \quad_counter1.a_delay_counter_11\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__29715\,
            I => \N__29711\
        );

    \I__3245\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29708\
        );

    \I__3244\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29705\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__29708\,
            I => \quad_counter1.a_delay_counter_4\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__29705\,
            I => \quad_counter1.a_delay_counter_4\
        );

    \I__3241\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29695\
        );

    \I__3240\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29690\
        );

    \I__3239\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29690\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__29695\,
            I => a_delay_counter_0_adj_4765
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__29690\,
            I => a_delay_counter_0_adj_4765
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__29685\,
            I => \N__29682\
        );

    \I__3235\ : InMux
    port map (
            O => \N__29682\,
            I => \N__29679\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__29679\,
            I => \quad_counter1.n25\
        );

    \I__3233\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29672\
        );

    \I__3232\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29669\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__29672\,
            I => \quad_counter1.a_delay_counter_9\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__29669\,
            I => \quad_counter1.a_delay_counter_9\
        );

    \I__3229\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29660\
        );

    \I__3228\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29657\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__29660\,
            I => \quad_counter1.a_delay_counter_6\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__29657\,
            I => \quad_counter1.a_delay_counter_6\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__29652\,
            I => \N__29648\
        );

    \I__3224\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29645\
        );

    \I__3223\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29642\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__29645\,
            I => \quad_counter1.a_delay_counter_12\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__29642\,
            I => \quad_counter1.a_delay_counter_12\
        );

    \I__3220\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29633\
        );

    \I__3219\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29630\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__29633\,
            I => \quad_counter1.a_delay_counter_13\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__29630\,
            I => \quad_counter1.a_delay_counter_13\
        );

    \I__3216\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29622\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__29622\,
            I => \quad_counter1.n26\
        );

    \I__3214\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29615\
        );

    \I__3213\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29612\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__29615\,
            I => \quad_counter1.a_delay_counter_8\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__29612\,
            I => \quad_counter1.a_delay_counter_8\
        );

    \I__3210\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29603\
        );

    \I__3209\ : InMux
    port map (
            O => \N__29606\,
            I => \N__29600\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__29603\,
            I => \quad_counter1.a_delay_counter_1\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__29600\,
            I => \quad_counter1.a_delay_counter_1\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__29595\,
            I => \N__29591\
        );

    \I__3205\ : InMux
    port map (
            O => \N__29594\,
            I => \N__29588\
        );

    \I__3204\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29585\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__29588\,
            I => \quad_counter1.a_delay_counter_2\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__29585\,
            I => \quad_counter1.a_delay_counter_2\
        );

    \I__3201\ : InMux
    port map (
            O => \N__29580\,
            I => \N__29576\
        );

    \I__3200\ : InMux
    port map (
            O => \N__29579\,
            I => \N__29573\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__29576\,
            I => \quad_counter1.a_delay_counter_3\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__29573\,
            I => \quad_counter1.a_delay_counter_3\
        );

    \I__3197\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__29565\,
            I => \quad_counter1.n28\
        );

    \I__3195\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29558\
        );

    \I__3194\ : InMux
    port map (
            O => \N__29561\,
            I => \N__29555\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__29558\,
            I => \quad_counter1.a_delay_counter_14\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__29555\,
            I => \quad_counter1.a_delay_counter_14\
        );

    \I__3191\ : InMux
    port map (
            O => \N__29550\,
            I => \N__29546\
        );

    \I__3190\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29543\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__29546\,
            I => \quad_counter1.a_delay_counter_7\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__29543\,
            I => \quad_counter1.a_delay_counter_7\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__29538\,
            I => \N__29534\
        );

    \I__3186\ : InMux
    port map (
            O => \N__29537\,
            I => \N__29531\
        );

    \I__3185\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29528\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__29531\,
            I => \quad_counter1.a_delay_counter_10\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__29528\,
            I => \quad_counter1.a_delay_counter_10\
        );

    \I__3182\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29519\
        );

    \I__3181\ : InMux
    port map (
            O => \N__29522\,
            I => \N__29516\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__29519\,
            I => \quad_counter1.a_delay_counter_15\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__29516\,
            I => \quad_counter1.a_delay_counter_15\
        );

    \I__3178\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29508\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__29508\,
            I => \quad_counter1.n27\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__29505\,
            I => \N__29502\
        );

    \I__3175\ : InMux
    port map (
            O => \N__29502\,
            I => \N__29498\
        );

    \I__3174\ : InMux
    port map (
            O => \N__29501\,
            I => \N__29495\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__29498\,
            I => \N__29491\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29488\
        );

    \I__3171\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29485\
        );

    \I__3170\ : Span12Mux_v
    port map (
            O => \N__29491\,
            I => \N__29482\
        );

    \I__3169\ : Span4Mux_h
    port map (
            O => \N__29488\,
            I => \N__29479\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__29485\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__3167\ : Odrv12
    port map (
            O => \N__29482\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__29479\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__3165\ : SRMux
    port map (
            O => \N__29472\,
            I => \N__29469\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__29469\,
            I => \N__29466\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__29466\,
            I => \N__29463\
        );

    \I__3162\ : Span4Mux_v
    port map (
            O => \N__29463\,
            I => \N__29460\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__29460\,
            I => \c0.n21573\
        );

    \I__3160\ : SRMux
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29451\
        );

    \I__3158\ : Span4Mux_h
    port map (
            O => \N__29451\,
            I => \N__29448\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__29448\,
            I => \c0.n21581\
        );

    \I__3156\ : SRMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__3154\ : Span4Mux_h
    port map (
            O => \N__29439\,
            I => \N__29436\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__29436\,
            I => \c0.n21575\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__3151\ : InMux
    port map (
            O => \N__29430\,
            I => \N__29426\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__29429\,
            I => \N__29423\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__29426\,
            I => \N__29420\
        );

    \I__3148\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29416\
        );

    \I__3147\ : Span4Mux_v
    port map (
            O => \N__29420\,
            I => \N__29413\
        );

    \I__3146\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29410\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__29416\,
            I => \N__29405\
        );

    \I__3144\ : Span4Mux_v
    port map (
            O => \N__29413\,
            I => \N__29405\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__29410\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__29405\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__3141\ : SRMux
    port map (
            O => \N__29400\,
            I => \N__29397\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__29397\,
            I => \N__29394\
        );

    \I__3139\ : Span4Mux_h
    port map (
            O => \N__29394\,
            I => \N__29391\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__29391\,
            I => \c0.n21577\
        );

    \I__3137\ : InMux
    port map (
            O => \N__29388\,
            I => \c0.n19796\
        );

    \I__3136\ : InMux
    port map (
            O => \N__29385\,
            I => \c0.n19797\
        );

    \I__3135\ : InMux
    port map (
            O => \N__29382\,
            I => \c0.n19798\
        );

    \I__3134\ : InMux
    port map (
            O => \N__29379\,
            I => \c0.n19799\
        );

    \I__3133\ : InMux
    port map (
            O => \N__29376\,
            I => \N__29372\
        );

    \I__3132\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29369\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__29372\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__29369\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__3129\ : InMux
    port map (
            O => \N__29364\,
            I => \c0.n19800\
        );

    \I__3128\ : InMux
    port map (
            O => \N__29361\,
            I => \c0.n19801\
        );

    \I__3127\ : InMux
    port map (
            O => \N__29358\,
            I => \N__29354\
        );

    \I__3126\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29351\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__29354\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__29351\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__3123\ : SRMux
    port map (
            O => \N__29346\,
            I => \N__29343\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__29343\,
            I => \N__29340\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__29340\,
            I => \N__29337\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__29337\,
            I => \c0.n21611\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__3118\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29327\
        );

    \I__3117\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29324\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__29327\,
            I => data_out_frame_12_6
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__29324\,
            I => data_out_frame_12_6
        );

    \I__3114\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29316\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__29316\,
            I => \c0.n5_adj_4334\
        );

    \I__3112\ : InMux
    port map (
            O => \N__29313\,
            I => \N__29310\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__29310\,
            I => \c0.n4_adj_4332\
        );

    \I__3110\ : InMux
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__29304\,
            I => \N__29301\
        );

    \I__3108\ : Span4Mux_v
    port map (
            O => \N__29301\,
            I => \N__29298\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__29298\,
            I => \c0.n26_adj_4662\
        );

    \I__3106\ : InMux
    port map (
            O => \N__29295\,
            I => \c0.n19795\
        );

    \I__3105\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29288\
        );

    \I__3104\ : InMux
    port map (
            O => \N__29291\,
            I => \N__29285\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__29288\,
            I => \N__29282\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__29285\,
            I => \r_Tx_Data_6\
        );

    \I__3101\ : Odrv12
    port map (
            O => \N__29282\,
            I => \r_Tx_Data_6\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__29277\,
            I => \N__29274\
        );

    \I__3099\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29270\
        );

    \I__3098\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29267\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__29270\,
            I => \N__29264\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__29267\,
            I => data_out_frame_5_2
        );

    \I__3095\ : Odrv12
    port map (
            O => \N__29264\,
            I => data_out_frame_5_2
        );

    \I__3094\ : InMux
    port map (
            O => \N__29259\,
            I => \N__29253\
        );

    \I__3093\ : InMux
    port map (
            O => \N__29258\,
            I => \N__29253\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__29250\,
            I => n17951
        );

    \I__3090\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29232\
        );

    \I__3089\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29232\
        );

    \I__3088\ : InMux
    port map (
            O => \N__29245\,
            I => \N__29232\
        );

    \I__3087\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29227\
        );

    \I__3086\ : InMux
    port map (
            O => \N__29243\,
            I => \N__29227\
        );

    \I__3085\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29224\
        );

    \I__3084\ : InMux
    port map (
            O => \N__29241\,
            I => \N__29221\
        );

    \I__3083\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29215\
        );

    \I__3082\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29215\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__29232\,
            I => \N__29209\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__29227\,
            I => \N__29206\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__29224\,
            I => \N__29203\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__29221\,
            I => \N__29200\
        );

    \I__3077\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29197\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__29215\,
            I => \N__29194\
        );

    \I__3075\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29187\
        );

    \I__3074\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29187\
        );

    \I__3073\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29187\
        );

    \I__3072\ : Span12Mux_s8_h
    port map (
            O => \N__29209\,
            I => \N__29180\
        );

    \I__3071\ : Sp12to4
    port map (
            O => \N__29206\,
            I => \N__29180\
        );

    \I__3070\ : Span12Mux_s11_v
    port map (
            O => \N__29203\,
            I => \N__29180\
        );

    \I__3069\ : Span4Mux_v
    port map (
            O => \N__29200\,
            I => \N__29175\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29175\
        );

    \I__3067\ : Span4Mux_h
    port map (
            O => \N__29194\,
            I => \N__29172\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__29187\,
            I => \r_SM_Main_1_adj_4774\
        );

    \I__3065\ : Odrv12
    port map (
            O => \N__29180\,
            I => \r_SM_Main_1_adj_4774\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__29175\,
            I => \r_SM_Main_1_adj_4774\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__29172\,
            I => \r_SM_Main_1_adj_4774\
        );

    \I__3062\ : InMux
    port map (
            O => \N__29163\,
            I => \N__29160\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__29160\,
            I => \N__29157\
        );

    \I__3060\ : Odrv12
    port map (
            O => \N__29157\,
            I => n25006
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__29154\,
            I => \N__29151\
        );

    \I__3058\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29148\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__29148\,
            I => \N__29145\
        );

    \I__3056\ : Span4Mux_h
    port map (
            O => \N__29145\,
            I => \N__29142\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__29142\,
            I => \c0.n11_adj_4663\
        );

    \I__3054\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29136\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__29136\,
            I => \N__29132\
        );

    \I__3052\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29129\
        );

    \I__3051\ : Span4Mux_v
    port map (
            O => \N__29132\,
            I => \N__29126\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__29129\,
            I => data_out_frame_5_1
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__29126\,
            I => data_out_frame_5_1
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__29121\,
            I => \N__29118\
        );

    \I__3047\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29112\
        );

    \I__3046\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29112\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__29112\,
            I => data_out_frame_13_3
        );

    \I__3044\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29105\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__29108\,
            I => \N__29102\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29099\
        );

    \I__3041\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29096\
        );

    \I__3040\ : Span4Mux_h
    port map (
            O => \N__29099\,
            I => \N__29093\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__29096\,
            I => data_out_frame_8_7
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__29093\,
            I => data_out_frame_8_7
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__29088\,
            I => \N__29085\
        );

    \I__3036\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29081\
        );

    \I__3035\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29078\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__29081\,
            I => \N__29075\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__29078\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__3032\ : Odrv12
    port map (
            O => \N__29075\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__3031\ : InMux
    port map (
            O => \N__29070\,
            I => \c0.tx.n19725\
        );

    \I__3030\ : InMux
    port map (
            O => \N__29067\,
            I => \N__29063\
        );

    \I__3029\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29060\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__29063\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__29060\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__3026\ : InMux
    port map (
            O => \N__29055\,
            I => \c0.tx.n19726\
        );

    \I__3025\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29048\
        );

    \I__3024\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29045\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__29048\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__29045\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__3021\ : InMux
    port map (
            O => \N__29040\,
            I => \c0.tx.n19727\
        );

    \I__3020\ : InMux
    port map (
            O => \N__29037\,
            I => \N__29033\
        );

    \I__3019\ : InMux
    port map (
            O => \N__29036\,
            I => \N__29030\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__29033\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__29030\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__3016\ : InMux
    port map (
            O => \N__29025\,
            I => \c0.tx.n19728\
        );

    \I__3015\ : InMux
    port map (
            O => \N__29022\,
            I => \N__29018\
        );

    \I__3014\ : InMux
    port map (
            O => \N__29021\,
            I => \N__29015\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__29018\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__29015\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__3011\ : InMux
    port map (
            O => \N__29010\,
            I => \c0.tx.n19729\
        );

    \I__3010\ : InMux
    port map (
            O => \N__29007\,
            I => \bfn_9_17_0_\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__29004\,
            I => \N__29000\
        );

    \I__3008\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28993\
        );

    \I__3007\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28993\
        );

    \I__3006\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28988\
        );

    \I__3005\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28988\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28984\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28981\
        );

    \I__3002\ : InMux
    port map (
            O => \N__28987\,
            I => \N__28978\
        );

    \I__3001\ : Span4Mux_v
    port map (
            O => \N__28984\,
            I => \N__28975\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__28981\,
            I => \N__28972\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__28978\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__28975\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__28972\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__2996\ : SRMux
    port map (
            O => \N__28965\,
            I => \N__28961\
        );

    \I__2995\ : SRMux
    port map (
            O => \N__28964\,
            I => \N__28958\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__28961\,
            I => \N__28955\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__28958\,
            I => \N__28952\
        );

    \I__2992\ : Span4Mux_h
    port map (
            O => \N__28955\,
            I => \N__28948\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__28952\,
            I => \N__28945\
        );

    \I__2990\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28942\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__28948\,
            I => \c0.tx.n17199\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__28945\,
            I => \c0.tx.n17199\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__28942\,
            I => \c0.tx.n17199\
        );

    \I__2986\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28932\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__28932\,
            I => \N__28929\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__28929\,
            I => \N__28926\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__28926\,
            I => \c0.tx.n4\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__28923\,
            I => \c0.tx.n14290_cascade_\
        );

    \I__2981\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28917\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__28917\,
            I => \N__28913\
        );

    \I__2979\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28910\
        );

    \I__2978\ : Span4Mux_h
    port map (
            O => \N__28913\,
            I => \N__28907\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__28910\,
            I => data_out_frame_6_7
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__28907\,
            I => data_out_frame_6_7
        );

    \I__2975\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28899\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__28899\,
            I => \c0.n26_adj_4645\
        );

    \I__2973\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28893\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__28893\,
            I => n24808
        );

    \I__2971\ : InMux
    port map (
            O => \N__28890\,
            I => \N__28887\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28884\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__28884\,
            I => n10_adj_4779
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__28881\,
            I => \c0.tx.n5_cascade_\
        );

    \I__2967\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28872\
        );

    \I__2966\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28865\
        );

    \I__2965\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28865\
        );

    \I__2964\ : InMux
    port map (
            O => \N__28875\,
            I => \N__28865\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__28872\,
            I => \N__28862\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__28865\,
            I => \N__28859\
        );

    \I__2961\ : Span4Mux_h
    port map (
            O => \N__28862\,
            I => \N__28856\
        );

    \I__2960\ : Span4Mux_h
    port map (
            O => \N__28859\,
            I => \N__28853\
        );

    \I__2959\ : Odrv4
    port map (
            O => \N__28856\,
            I => \c0.tx.n17904\
        );

    \I__2958\ : Odrv4
    port map (
            O => \N__28853\,
            I => \c0.tx.n17904\
        );

    \I__2957\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28845\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__28845\,
            I => \N__28842\
        );

    \I__2955\ : Odrv12
    port map (
            O => \N__28842\,
            I => \c0.tx.n25051\
        );

    \I__2954\ : InMux
    port map (
            O => \N__28839\,
            I => \bfn_9_16_0_\
        );

    \I__2953\ : InMux
    port map (
            O => \N__28836\,
            I => \N__28832\
        );

    \I__2952\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28829\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__28832\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__28829\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__2949\ : InMux
    port map (
            O => \N__28824\,
            I => \c0.tx.n19723\
        );

    \I__2948\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28817\
        );

    \I__2947\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28814\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__28817\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__28814\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__2944\ : InMux
    port map (
            O => \N__28809\,
            I => \c0.tx.n19724\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__28806\,
            I => \n10_adj_4776_cascade_\
        );

    \I__2942\ : InMux
    port map (
            O => \N__28803\,
            I => \N__28797\
        );

    \I__2941\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28797\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__28797\,
            I => \r_Tx_Data_5\
        );

    \I__2939\ : InMux
    port map (
            O => \N__28794\,
            I => \N__28791\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__28791\,
            I => \c0.tx.n25077\
        );

    \I__2937\ : InMux
    port map (
            O => \N__28788\,
            I => \N__28782\
        );

    \I__2936\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28782\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__28782\,
            I => \r_Tx_Data_7\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__28779\,
            I => \N__28775\
        );

    \I__2933\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28771\
        );

    \I__2932\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28768\
        );

    \I__2931\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28763\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__28771\,
            I => \N__28758\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28758\
        );

    \I__2928\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28752\
        );

    \I__2927\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28752\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__28763\,
            I => \N__28749\
        );

    \I__2925\ : Span4Mux_v
    port map (
            O => \N__28758\,
            I => \N__28746\
        );

    \I__2924\ : InMux
    port map (
            O => \N__28757\,
            I => \N__28743\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28740\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__28749\,
            I => \N__28735\
        );

    \I__2921\ : Span4Mux_h
    port map (
            O => \N__28746\,
            I => \N__28735\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__28743\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__28740\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__28735\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__28728\,
            I => \N__28723\
        );

    \I__2916\ : InMux
    port map (
            O => \N__28727\,
            I => \N__28716\
        );

    \I__2915\ : InMux
    port map (
            O => \N__28726\,
            I => \N__28713\
        );

    \I__2914\ : InMux
    port map (
            O => \N__28723\,
            I => \N__28710\
        );

    \I__2913\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28701\
        );

    \I__2912\ : InMux
    port map (
            O => \N__28721\,
            I => \N__28701\
        );

    \I__2911\ : InMux
    port map (
            O => \N__28720\,
            I => \N__28701\
        );

    \I__2910\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28701\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__28716\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__28713\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__28710\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__28701\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__2905\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__28689\,
            I => \c0.tx.n25074\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__28686\,
            I => \N__28680\
        );

    \I__2902\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28676\
        );

    \I__2901\ : InMux
    port map (
            O => \N__28684\,
            I => \N__28673\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__28683\,
            I => \N__28670\
        );

    \I__2899\ : InMux
    port map (
            O => \N__28680\,
            I => \N__28663\
        );

    \I__2898\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28660\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__28676\,
            I => \N__28655\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__28673\,
            I => \N__28655\
        );

    \I__2895\ : InMux
    port map (
            O => \N__28670\,
            I => \N__28652\
        );

    \I__2894\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28649\
        );

    \I__2893\ : InMux
    port map (
            O => \N__28668\,
            I => \N__28644\
        );

    \I__2892\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28644\
        );

    \I__2891\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28641\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28636\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__28660\,
            I => \N__28636\
        );

    \I__2888\ : Span4Mux_v
    port map (
            O => \N__28655\,
            I => \N__28633\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__28652\,
            I => \N__28626\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__28649\,
            I => \N__28626\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__28644\,
            I => \N__28626\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__28641\,
            I => \r_SM_Main_0\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__28636\,
            I => \r_SM_Main_0\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__28633\,
            I => \r_SM_Main_0\
        );

    \I__2881\ : Odrv12
    port map (
            O => \N__28626\,
            I => \r_SM_Main_0\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__28617\,
            I => \c0.n24960_cascade_\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__28614\,
            I => \c0.n24806_cascade_\
        );

    \I__2878\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__28608\,
            I => \N__28605\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__28605\,
            I => n24757
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__28602\,
            I => \n3_cascade_\
        );

    \I__2874\ : IoInMux
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__28596\,
            I => \N__28593\
        );

    \I__2872\ : IoSpan4Mux
    port map (
            O => \N__28593\,
            I => \N__28589\
        );

    \I__2871\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28586\
        );

    \I__2870\ : Span4Mux_s0_h
    port map (
            O => \N__28589\,
            I => \N__28581\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__28586\,
            I => \N__28581\
        );

    \I__2868\ : Span4Mux_h
    port map (
            O => \N__28581\,
            I => \N__28578\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__2866\ : Span4Mux_h
    port map (
            O => \N__28575\,
            I => \N__28571\
        );

    \I__2865\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28568\
        );

    \I__2864\ : Odrv4
    port map (
            O => \N__28571\,
            I => tx_o
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__28568\,
            I => tx_o
        );

    \I__2862\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28560\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__28560\,
            I => \N__28556\
        );

    \I__2860\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28553\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__28556\,
            I => \N__28550\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__28553\,
            I => \r_Tx_Data_3\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__28550\,
            I => \r_Tx_Data_3\
        );

    \I__2856\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28542\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__28542\,
            I => \c0.tx.n19492\
        );

    \I__2854\ : InMux
    port map (
            O => \N__28539\,
            I => \N__28536\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__2852\ : Span4Mux_v
    port map (
            O => \N__28533\,
            I => \N__28527\
        );

    \I__2851\ : InMux
    port map (
            O => \N__28532\,
            I => \N__28520\
        );

    \I__2850\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28520\
        );

    \I__2849\ : InMux
    port map (
            O => \N__28530\,
            I => \N__28520\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__28527\,
            I => \c0.tx.n22949\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__28520\,
            I => \c0.tx.n22949\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__28515\,
            I => \c0.tx.n19492_cascade_\
        );

    \I__2845\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28509\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__28509\,
            I => \N__28505\
        );

    \I__2843\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28502\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__28505\,
            I => \N__28499\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__28502\,
            I => \r_Tx_Data_1\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__28499\,
            I => \r_Tx_Data_1\
        );

    \I__2839\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28491\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__28491\,
            I => \c0.tx.n25080\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__28488\,
            I => \c0.tx.n25083_cascade_\
        );

    \I__2836\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__28482\,
            I => \c0.tx.o_Tx_Serial_N_3782\
        );

    \I__2834\ : InMux
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__28476\,
            I => \N__28473\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__28473\,
            I => \N__28470\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__28470\,
            I => n10
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__28467\,
            I => \N__28464\
        );

    \I__2829\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28459\
        );

    \I__2828\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28454\
        );

    \I__2827\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28454\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__28459\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__28454\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__28449\,
            I => \N__28446\
        );

    \I__2823\ : InMux
    port map (
            O => \N__28446\,
            I => \N__28443\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__28443\,
            I => \N__28440\
        );

    \I__2821\ : Span4Mux_v
    port map (
            O => \N__28440\,
            I => \N__28436\
        );

    \I__2820\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28433\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__28436\,
            I => \c0.tx.n17832\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__28433\,
            I => \c0.tx.n17832\
        );

    \I__2817\ : InMux
    port map (
            O => \N__28428\,
            I => \quad_counter1.n19714\
        );

    \I__2816\ : InMux
    port map (
            O => \N__28425\,
            I => \quad_counter1.n19715\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__28422\,
            I => \N__28419\
        );

    \I__2814\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28415\
        );

    \I__2813\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28411\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__28415\,
            I => \N__28407\
        );

    \I__2811\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28402\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__28411\,
            I => \N__28399\
        );

    \I__2809\ : InMux
    port map (
            O => \N__28410\,
            I => \N__28396\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__28407\,
            I => \N__28393\
        );

    \I__2807\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28390\
        );

    \I__2806\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28387\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__28402\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__28399\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__28396\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__28393\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__28390\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__28387\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__2799\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28369\
        );

    \I__2798\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28366\
        );

    \I__2797\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28363\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__28369\,
            I => \N__28358\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__28366\,
            I => \N__28358\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__28363\,
            I => \N__28352\
        );

    \I__2793\ : Span4Mux_h
    port map (
            O => \N__28358\,
            I => \N__28352\
        );

    \I__2792\ : InMux
    port map (
            O => \N__28357\,
            I => \N__28349\
        );

    \I__2791\ : Span4Mux_v
    port map (
            O => \N__28352\,
            I => \N__28346\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__28349\,
            I => \r_SM_Main_2_N_3751_1\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__28346\,
            I => \r_SM_Main_2_N_3751_1\
        );

    \I__2788\ : InMux
    port map (
            O => \N__28341\,
            I => \N__28338\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__28338\,
            I => \c0.tx.n3843\
        );

    \I__2786\ : InMux
    port map (
            O => \N__28335\,
            I => \quad_counter1.n19705\
        );

    \I__2785\ : InMux
    port map (
            O => \N__28332\,
            I => \quad_counter1.n19706\
        );

    \I__2784\ : InMux
    port map (
            O => \N__28329\,
            I => \quad_counter1.n19707\
        );

    \I__2783\ : InMux
    port map (
            O => \N__28326\,
            I => \bfn_9_8_0_\
        );

    \I__2782\ : InMux
    port map (
            O => \N__28323\,
            I => \quad_counter1.n19709\
        );

    \I__2781\ : InMux
    port map (
            O => \N__28320\,
            I => \quad_counter1.n19710\
        );

    \I__2780\ : InMux
    port map (
            O => \N__28317\,
            I => \quad_counter1.n19711\
        );

    \I__2779\ : InMux
    port map (
            O => \N__28314\,
            I => \quad_counter1.n19712\
        );

    \I__2778\ : InMux
    port map (
            O => \N__28311\,
            I => \quad_counter1.n19713\
        );

    \I__2777\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28304\
        );

    \I__2776\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28301\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__28304\,
            I => \N__28298\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__28301\,
            I => data_out_frame_9_7
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__28298\,
            I => data_out_frame_9_7
        );

    \I__2772\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28290\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__28290\,
            I => \N__28287\
        );

    \I__2770\ : Odrv12
    port map (
            O => \N__28287\,
            I => \c0.rx.n24875\
        );

    \I__2769\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28281\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__28281\,
            I => \c0.rx.n25068\
        );

    \I__2767\ : InMux
    port map (
            O => \N__28278\,
            I => \bfn_9_7_0_\
        );

    \I__2766\ : InMux
    port map (
            O => \N__28275\,
            I => \quad_counter1.n19701\
        );

    \I__2765\ : InMux
    port map (
            O => \N__28272\,
            I => \quad_counter1.n19702\
        );

    \I__2764\ : InMux
    port map (
            O => \N__28269\,
            I => \quad_counter1.n19703\
        );

    \I__2763\ : InMux
    port map (
            O => \N__28266\,
            I => \quad_counter1.n19704\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__28263\,
            I => \c0.n25104_cascade_\
        );

    \I__2761\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28254\
        );

    \I__2759\ : Odrv12
    port map (
            O => \N__28254\,
            I => \c0.n25107\
        );

    \I__2758\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28247\
        );

    \I__2757\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28244\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__28247\,
            I => \N__28241\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__28244\,
            I => data_out_frame_5_7
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__28241\,
            I => data_out_frame_5_7
        );

    \I__2753\ : InMux
    port map (
            O => \N__28236\,
            I => \N__28233\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__28233\,
            I => n25071
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__28230\,
            I => \n3821_cascade_\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__28227\,
            I => \c0.tx.n6_cascade_\
        );

    \I__2749\ : InMux
    port map (
            O => \N__28224\,
            I => \N__28221\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__28221\,
            I => \N__28218\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__28218\,
            I => \c0.n25089\
        );

    \I__2746\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__28212\,
            I => \N__28209\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__28209\,
            I => n25018
        );

    \I__2743\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28203\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__28203\,
            I => \c0.tx.n23980\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__28200\,
            I => \c0.n5_adj_4712_cascade_\
        );

    \I__2740\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28194\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__28194\,
            I => \N__28191\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__28191\,
            I => \c0.n24800\
        );

    \I__2737\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28185\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__28185\,
            I => \N__28182\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__28182\,
            I => \c0.tx.n5_adj_4207\
        );

    \I__2734\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28176\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__28176\,
            I => \c0.n24949\
        );

    \I__2732\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__28170\,
            I => \N__28167\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__28167\,
            I => n10_adj_4777
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__28164\,
            I => \c0.n25086_cascade_\
        );

    \I__2728\ : InMux
    port map (
            O => \N__28161\,
            I => \N__28157\
        );

    \I__2727\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28154\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__28157\,
            I => data_out_frame_9_3
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__28154\,
            I => data_out_frame_9_3
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__28149\,
            I => \n24802_cascade_\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \c0.n11_adj_4715_cascade_\
        );

    \I__2722\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28140\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__28140\,
            I => n25010
        );

    \I__2720\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28130\
        );

    \I__2719\ : InMux
    port map (
            O => \N__28136\,
            I => \N__28125\
        );

    \I__2718\ : InMux
    port map (
            O => \N__28135\,
            I => \N__28125\
        );

    \I__2717\ : InMux
    port map (
            O => \N__28134\,
            I => \N__28122\
        );

    \I__2716\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28119\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__28130\,
            I => \N__28114\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__28125\,
            I => \N__28114\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__28122\,
            I => \N__28111\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28106\
        );

    \I__2711\ : Span4Mux_h
    port map (
            O => \N__28114\,
            I => \N__28106\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__28111\,
            I => \A_filtered\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__28106\,
            I => \A_filtered\
        );

    \I__2708\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28098\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__28098\,
            I => n8628
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__28095\,
            I => \n9603_cascade_\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__28092\,
            I => \N__28087\
        );

    \I__2704\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28084\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__28090\,
            I => \N__28081\
        );

    \I__2702\ : InMux
    port map (
            O => \N__28087\,
            I => \N__28078\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__28084\,
            I => \N__28075\
        );

    \I__2700\ : InMux
    port map (
            O => \N__28081\,
            I => \N__28072\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__28078\,
            I => \B_filtered\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__28075\,
            I => \B_filtered\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__28072\,
            I => \B_filtered\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__28065\,
            I => \N__28061\
        );

    \I__2695\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28057\
        );

    \I__2694\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28052\
        );

    \I__2693\ : InMux
    port map (
            O => \N__28060\,
            I => \N__28052\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28047\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__28052\,
            I => \N__28047\
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__28047\,
            I => \quad_counter0.B_delayed\
        );

    \I__2689\ : InMux
    port map (
            O => \N__28044\,
            I => \quad_counter0.n19685\
        );

    \I__2688\ : InMux
    port map (
            O => \N__28041\,
            I => \N__28037\
        );

    \I__2687\ : InMux
    port map (
            O => \N__28040\,
            I => \N__28034\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__28037\,
            I => \quad_counter0.a_delay_counter_15\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__28034\,
            I => \quad_counter0.a_delay_counter_15\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__28029\,
            I => \N__28026\
        );

    \I__2683\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28021\
        );

    \I__2682\ : CEMux
    port map (
            O => \N__28025\,
            I => \N__28018\
        );

    \I__2681\ : CEMux
    port map (
            O => \N__28024\,
            I => \N__28015\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__28021\,
            I => n14469
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__28018\,
            I => n14469
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__28015\,
            I => n14469
        );

    \I__2677\ : SRMux
    port map (
            O => \N__28008\,
            I => \N__28004\
        );

    \I__2676\ : InMux
    port map (
            O => \N__28007\,
            I => \N__28000\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__28004\,
            I => \N__27997\
        );

    \I__2674\ : SRMux
    port map (
            O => \N__28003\,
            I => \N__27994\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__28000\,
            I => \N__27991\
        );

    \I__2672\ : Odrv12
    port map (
            O => \N__27997\,
            I => \a_delay_counter_15__N_4123\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__27994\,
            I => \a_delay_counter_15__N_4123\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__27991\,
            I => \a_delay_counter_15__N_4123\
        );

    \I__2669\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27980\
        );

    \I__2668\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27977\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__27980\,
            I => \N__27974\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__27977\,
            I => \quad_counter1.b_delay_counter_13\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__27974\,
            I => \quad_counter1.b_delay_counter_13\
        );

    \I__2664\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27965\
        );

    \I__2663\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27962\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__27965\,
            I => \quad_counter1.b_delay_counter_1\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__27962\,
            I => \quad_counter1.b_delay_counter_1\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__27957\,
            I => \N__27953\
        );

    \I__2659\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27950\
        );

    \I__2658\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27947\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__27950\,
            I => \quad_counter1.b_delay_counter_2\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__27947\,
            I => \quad_counter1.b_delay_counter_2\
        );

    \I__2655\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27938\
        );

    \I__2654\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27935\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__27938\,
            I => \quad_counter1.b_delay_counter_5\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__27935\,
            I => \quad_counter1.b_delay_counter_5\
        );

    \I__2651\ : InMux
    port map (
            O => \N__27930\,
            I => \N__27927\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__27927\,
            I => \N__27924\
        );

    \I__2649\ : Odrv4
    port map (
            O => \N__27924\,
            I => \quad_counter1.n28_adj_4199\
        );

    \I__2648\ : InMux
    port map (
            O => \N__27921\,
            I => \N__27916\
        );

    \I__2647\ : InMux
    port map (
            O => \N__27920\,
            I => \N__27913\
        );

    \I__2646\ : InMux
    port map (
            O => \N__27919\,
            I => \N__27910\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27904\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__27913\,
            I => \N__27904\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__27910\,
            I => \N__27901\
        );

    \I__2642\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27898\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__27904\,
            I => \N__27891\
        );

    \I__2640\ : Span4Mux_h
    port map (
            O => \N__27901\,
            I => \N__27891\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__27898\,
            I => \N__27891\
        );

    \I__2638\ : Span4Mux_h
    port map (
            O => \N__27891\,
            I => \N__27888\
        );

    \I__2637\ : Span4Mux_v
    port map (
            O => \N__27888\,
            I => \N__27885\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__27885\,
            I => \PIN_7_c\
        );

    \I__2635\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27878\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__27881\,
            I => \N__27875\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__27878\,
            I => \N__27872\
        );

    \I__2632\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27868\
        );

    \I__2631\ : Span4Mux_h
    port map (
            O => \N__27872\,
            I => \N__27865\
        );

    \I__2630\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27862\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__27868\,
            I => \quadA_delayed\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__27865\,
            I => \quadA_delayed\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__27862\,
            I => \quadA_delayed\
        );

    \I__2626\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27851\
        );

    \I__2625\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27848\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__27851\,
            I => \quad_counter1.b_delay_counter_14\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__27848\,
            I => \quad_counter1.b_delay_counter_14\
        );

    \I__2622\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27839\
        );

    \I__2621\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27836\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__27839\,
            I => \quad_counter1.b_delay_counter_7\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__27836\,
            I => \quad_counter1.b_delay_counter_7\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__27831\,
            I => \N__27827\
        );

    \I__2617\ : InMux
    port map (
            O => \N__27830\,
            I => \N__27824\
        );

    \I__2616\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27821\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__27824\,
            I => \quad_counter1.b_delay_counter_12\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__27821\,
            I => \quad_counter1.b_delay_counter_12\
        );

    \I__2613\ : InMux
    port map (
            O => \N__27816\,
            I => \N__27812\
        );

    \I__2612\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27809\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__27812\,
            I => \quad_counter1.b_delay_counter_15\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__27809\,
            I => \quad_counter1.b_delay_counter_15\
        );

    \I__2609\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27801\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__27801\,
            I => \quad_counter1.n27_adj_4201\
        );

    \I__2607\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27794\
        );

    \I__2606\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27791\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__27794\,
            I => \quad_counter0.a_delay_counter_7\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__27791\,
            I => \quad_counter0.a_delay_counter_7\
        );

    \I__2603\ : InMux
    port map (
            O => \N__27786\,
            I => \quad_counter0.n19677\
        );

    \I__2602\ : InMux
    port map (
            O => \N__27783\,
            I => \N__27779\
        );

    \I__2601\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27776\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__27779\,
            I => \quad_counter0.a_delay_counter_8\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__27776\,
            I => \quad_counter0.a_delay_counter_8\
        );

    \I__2598\ : InMux
    port map (
            O => \N__27771\,
            I => \bfn_6_14_0_\
        );

    \I__2597\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27764\
        );

    \I__2596\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27761\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__27764\,
            I => \quad_counter0.a_delay_counter_9\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__27761\,
            I => \quad_counter0.a_delay_counter_9\
        );

    \I__2593\ : InMux
    port map (
            O => \N__27756\,
            I => \quad_counter0.n19679\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__27753\,
            I => \N__27749\
        );

    \I__2591\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27746\
        );

    \I__2590\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27743\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__27746\,
            I => \quad_counter0.a_delay_counter_10\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__27743\,
            I => \quad_counter0.a_delay_counter_10\
        );

    \I__2587\ : InMux
    port map (
            O => \N__27738\,
            I => \quad_counter0.n19680\
        );

    \I__2586\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27731\
        );

    \I__2585\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27728\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__27731\,
            I => \quad_counter0.a_delay_counter_11\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__27728\,
            I => \quad_counter0.a_delay_counter_11\
        );

    \I__2582\ : InMux
    port map (
            O => \N__27723\,
            I => \quad_counter0.n19681\
        );

    \I__2581\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27716\
        );

    \I__2580\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27713\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__27716\,
            I => \quad_counter0.a_delay_counter_12\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__27713\,
            I => \quad_counter0.a_delay_counter_12\
        );

    \I__2577\ : InMux
    port map (
            O => \N__27708\,
            I => \quad_counter0.n19682\
        );

    \I__2576\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27701\
        );

    \I__2575\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27698\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__27701\,
            I => \quad_counter0.a_delay_counter_13\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__27698\,
            I => \quad_counter0.a_delay_counter_13\
        );

    \I__2572\ : InMux
    port map (
            O => \N__27693\,
            I => \quad_counter0.n19683\
        );

    \I__2571\ : InMux
    port map (
            O => \N__27690\,
            I => \N__27686\
        );

    \I__2570\ : InMux
    port map (
            O => \N__27689\,
            I => \N__27683\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__27686\,
            I => \quad_counter0.a_delay_counter_14\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__27683\,
            I => \quad_counter0.a_delay_counter_14\
        );

    \I__2567\ : InMux
    port map (
            O => \N__27678\,
            I => \quad_counter0.n19684\
        );

    \I__2566\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27671\
        );

    \I__2565\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27668\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__27671\,
            I => \quad_counter0.b_delay_counter_10\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__27668\,
            I => \quad_counter0.b_delay_counter_10\
        );

    \I__2562\ : InMux
    port map (
            O => \N__27663\,
            I => \N__27659\
        );

    \I__2561\ : InMux
    port map (
            O => \N__27662\,
            I => \N__27656\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__27659\,
            I => \quad_counter0.b_delay_counter_11\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__27656\,
            I => \quad_counter0.b_delay_counter_11\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__27651\,
            I => \quad_counter0.n24_adj_4758_cascade_\
        );

    \I__2557\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27645\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__27645\,
            I => \quad_counter0.n18\
        );

    \I__2555\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27639\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__27639\,
            I => \quad_counter0.n26_adj_4759\
        );

    \I__2553\ : InMux
    port map (
            O => \N__27636\,
            I => \N__27631\
        );

    \I__2552\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27626\
        );

    \I__2551\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27626\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__27631\,
            I => a_delay_counter_0
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__27626\,
            I => a_delay_counter_0
        );

    \I__2548\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__27618\,
            I => \N__27615\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__27615\,
            I => n39
        );

    \I__2545\ : InMux
    port map (
            O => \N__27612\,
            I => \bfn_6_13_0_\
        );

    \I__2544\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27605\
        );

    \I__2543\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27602\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__27605\,
            I => \quad_counter0.a_delay_counter_1\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__27602\,
            I => \quad_counter0.a_delay_counter_1\
        );

    \I__2540\ : InMux
    port map (
            O => \N__27597\,
            I => \quad_counter0.n19671\
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__27594\,
            I => \N__27590\
        );

    \I__2538\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27587\
        );

    \I__2537\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27584\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__27587\,
            I => \quad_counter0.a_delay_counter_2\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__27584\,
            I => \quad_counter0.a_delay_counter_2\
        );

    \I__2534\ : InMux
    port map (
            O => \N__27579\,
            I => \quad_counter0.n19672\
        );

    \I__2533\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27572\
        );

    \I__2532\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27569\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__27572\,
            I => \quad_counter0.a_delay_counter_3\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__27569\,
            I => \quad_counter0.a_delay_counter_3\
        );

    \I__2529\ : InMux
    port map (
            O => \N__27564\,
            I => \quad_counter0.n19673\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__27561\,
            I => \N__27557\
        );

    \I__2527\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27554\
        );

    \I__2526\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27551\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__27554\,
            I => \quad_counter0.a_delay_counter_4\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__27551\,
            I => \quad_counter0.a_delay_counter_4\
        );

    \I__2523\ : InMux
    port map (
            O => \N__27546\,
            I => \quad_counter0.n19674\
        );

    \I__2522\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27539\
        );

    \I__2521\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27536\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__27539\,
            I => \quad_counter0.a_delay_counter_5\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__27536\,
            I => \quad_counter0.a_delay_counter_5\
        );

    \I__2518\ : InMux
    port map (
            O => \N__27531\,
            I => \quad_counter0.n19675\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__27528\,
            I => \N__27524\
        );

    \I__2516\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27521\
        );

    \I__2515\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27518\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__27521\,
            I => \quad_counter0.a_delay_counter_6\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__27518\,
            I => \quad_counter0.a_delay_counter_6\
        );

    \I__2512\ : InMux
    port map (
            O => \N__27513\,
            I => \quad_counter0.n19676\
        );

    \I__2511\ : InMux
    port map (
            O => \N__27510\,
            I => \quad_counter0.n19666\
        );

    \I__2510\ : InMux
    port map (
            O => \N__27507\,
            I => \quad_counter0.n19667\
        );

    \I__2509\ : InMux
    port map (
            O => \N__27504\,
            I => \N__27500\
        );

    \I__2508\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27497\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__27500\,
            I => \quad_counter0.b_delay_counter_13\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__27497\,
            I => \quad_counter0.b_delay_counter_13\
        );

    \I__2505\ : InMux
    port map (
            O => \N__27492\,
            I => \quad_counter0.n19668\
        );

    \I__2504\ : InMux
    port map (
            O => \N__27489\,
            I => \quad_counter0.n19669\
        );

    \I__2503\ : InMux
    port map (
            O => \N__27486\,
            I => \quad_counter0.n19670\
        );

    \I__2502\ : CEMux
    port map (
            O => \N__27483\,
            I => \N__27479\
        );

    \I__2501\ : CEMux
    port map (
            O => \N__27482\,
            I => \N__27476\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__27479\,
            I => \N__27473\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__27476\,
            I => \N__27470\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__27473\,
            I => \N__27466\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__27470\,
            I => \N__27463\
        );

    \I__2496\ : InMux
    port map (
            O => \N__27469\,
            I => \N__27460\
        );

    \I__2495\ : Odrv4
    port map (
            O => \N__27466\,
            I => n14315
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__27463\,
            I => n14315
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__27460\,
            I => n14315
        );

    \I__2492\ : SRMux
    port map (
            O => \N__27453\,
            I => \N__27449\
        );

    \I__2491\ : SRMux
    port map (
            O => \N__27452\,
            I => \N__27445\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__27449\,
            I => \N__27442\
        );

    \I__2489\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27439\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27435\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__27442\,
            I => \N__27432\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__27439\,
            I => \N__27429\
        );

    \I__2485\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27426\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__27435\,
            I => \b_delay_counter_15__N_4140\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__27432\,
            I => \b_delay_counter_15__N_4140\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__27429\,
            I => \b_delay_counter_15__N_4140\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__27426\,
            I => \b_delay_counter_15__N_4140\
        );

    \I__2480\ : InMux
    port map (
            O => \N__27417\,
            I => \N__27413\
        );

    \I__2479\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27408\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__27413\,
            I => \N__27405\
        );

    \I__2477\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27402\
        );

    \I__2476\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27399\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__27408\,
            I => \N__27392\
        );

    \I__2474\ : Span4Mux_h
    port map (
            O => \N__27405\,
            I => \N__27392\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__27402\,
            I => \N__27392\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__27399\,
            I => \N__27389\
        );

    \I__2471\ : Sp12to4
    port map (
            O => \N__27392\,
            I => \N__27386\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__27389\,
            I => \N__27383\
        );

    \I__2469\ : Span12Mux_v
    port map (
            O => \N__27386\,
            I => \N__27380\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__27383\,
            I => \N__27377\
        );

    \I__2467\ : Odrv12
    port map (
            O => \N__27380\,
            I => \PIN_8_c\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__27377\,
            I => \PIN_8_c\
        );

    \I__2465\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27369\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__27369\,
            I => \N__27365\
        );

    \I__2463\ : InMux
    port map (
            O => \N__27368\,
            I => \N__27362\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__27365\,
            I => \N__27358\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27355\
        );

    \I__2460\ : InMux
    port map (
            O => \N__27361\,
            I => \N__27352\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__27358\,
            I => \quadB_delayed\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__27355\,
            I => \quadB_delayed\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__27352\,
            I => \quadB_delayed\
        );

    \I__2456\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27342\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__27342\,
            I => n12942
        );

    \I__2454\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27335\
        );

    \I__2453\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27332\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__27335\,
            I => \quad_counter0.b_delay_counter_15\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__27332\,
            I => \quad_counter0.b_delay_counter_15\
        );

    \I__2450\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27323\
        );

    \I__2449\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27320\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__27323\,
            I => \quad_counter0.b_delay_counter_8\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__27320\,
            I => \quad_counter0.b_delay_counter_8\
        );

    \I__2446\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27312\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__27312\,
            I => \quad_counter0.A_delayed\
        );

    \I__2444\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27305\
        );

    \I__2443\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27302\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__27305\,
            I => \N__27299\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__27302\,
            I => \quad_counter0.b_delay_counter_7\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__27299\,
            I => \quad_counter0.b_delay_counter_7\
        );

    \I__2439\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27290\
        );

    \I__2438\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27287\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__27290\,
            I => \quad_counter0.b_delay_counter_12\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__27287\,
            I => \quad_counter0.b_delay_counter_12\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__2434\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27275\
        );

    \I__2433\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27272\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__27275\,
            I => \N__27269\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__27272\,
            I => \quad_counter0.b_delay_counter_5\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__27269\,
            I => \quad_counter0.b_delay_counter_5\
        );

    \I__2429\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27260\
        );

    \I__2428\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27257\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__27260\,
            I => \quad_counter0.b_delay_counter_14\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__27257\,
            I => \quad_counter0.b_delay_counter_14\
        );

    \I__2425\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27248\
        );

    \I__2424\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27245\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__27248\,
            I => \quad_counter0.b_delay_counter_2\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__27245\,
            I => \quad_counter0.b_delay_counter_2\
        );

    \I__2421\ : InMux
    port map (
            O => \N__27240\,
            I => \quad_counter0.n19657\
        );

    \I__2420\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27233\
        );

    \I__2419\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27230\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__27233\,
            I => \quad_counter0.b_delay_counter_3\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__27230\,
            I => \quad_counter0.b_delay_counter_3\
        );

    \I__2416\ : InMux
    port map (
            O => \N__27225\,
            I => \quad_counter0.n19658\
        );

    \I__2415\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27218\
        );

    \I__2414\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27215\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__27218\,
            I => \quad_counter0.b_delay_counter_4\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__27215\,
            I => \quad_counter0.b_delay_counter_4\
        );

    \I__2411\ : InMux
    port map (
            O => \N__27210\,
            I => \quad_counter0.n19659\
        );

    \I__2410\ : InMux
    port map (
            O => \N__27207\,
            I => \quad_counter0.n19660\
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__27204\,
            I => \N__27200\
        );

    \I__2408\ : InMux
    port map (
            O => \N__27203\,
            I => \N__27197\
        );

    \I__2407\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27194\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__27197\,
            I => \quad_counter0.b_delay_counter_6\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__27194\,
            I => \quad_counter0.b_delay_counter_6\
        );

    \I__2404\ : InMux
    port map (
            O => \N__27189\,
            I => \quad_counter0.n19661\
        );

    \I__2403\ : InMux
    port map (
            O => \N__27186\,
            I => \quad_counter0.n19662\
        );

    \I__2402\ : InMux
    port map (
            O => \N__27183\,
            I => \bfn_6_11_0_\
        );

    \I__2401\ : InMux
    port map (
            O => \N__27180\,
            I => \N__27176\
        );

    \I__2400\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27173\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__27176\,
            I => \quad_counter0.b_delay_counter_9\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__27173\,
            I => \quad_counter0.b_delay_counter_9\
        );

    \I__2397\ : InMux
    port map (
            O => \N__27168\,
            I => \quad_counter0.n19664\
        );

    \I__2396\ : InMux
    port map (
            O => \N__27165\,
            I => \quad_counter0.n19665\
        );

    \I__2395\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27158\
        );

    \I__2394\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27155\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__27158\,
            I => \N__27152\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__27155\,
            I => \quad_counter1.b_delay_counter_10\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__27152\,
            I => \quad_counter1.b_delay_counter_10\
        );

    \I__2390\ : InMux
    port map (
            O => \N__27147\,
            I => \quad_counter1.n19695\
        );

    \I__2389\ : InMux
    port map (
            O => \N__27144\,
            I => \N__27140\
        );

    \I__2388\ : InMux
    port map (
            O => \N__27143\,
            I => \N__27137\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__27140\,
            I => \N__27134\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__27137\,
            I => \quad_counter1.b_delay_counter_11\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__27134\,
            I => \quad_counter1.b_delay_counter_11\
        );

    \I__2384\ : InMux
    port map (
            O => \N__27129\,
            I => \quad_counter1.n19696\
        );

    \I__2383\ : InMux
    port map (
            O => \N__27126\,
            I => \quad_counter1.n19697\
        );

    \I__2382\ : InMux
    port map (
            O => \N__27123\,
            I => \quad_counter1.n19698\
        );

    \I__2381\ : InMux
    port map (
            O => \N__27120\,
            I => \quad_counter1.n19699\
        );

    \I__2380\ : InMux
    port map (
            O => \N__27117\,
            I => \quad_counter1.n19700\
        );

    \I__2379\ : CEMux
    port map (
            O => \N__27114\,
            I => \N__27110\
        );

    \I__2378\ : CEMux
    port map (
            O => \N__27113\,
            I => \N__27107\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__27110\,
            I => \N__27104\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27101\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__27104\,
            I => n14425
        );

    \I__2374\ : Odrv12
    port map (
            O => \N__27101\,
            I => n14425
        );

    \I__2373\ : SRMux
    port map (
            O => \N__27096\,
            I => \N__27092\
        );

    \I__2372\ : SRMux
    port map (
            O => \N__27095\,
            I => \N__27089\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__27092\,
            I => \N__27086\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__27089\,
            I => \N__27083\
        );

    \I__2369\ : Span4Mux_v
    port map (
            O => \N__27086\,
            I => \N__27077\
        );

    \I__2368\ : Span4Mux_h
    port map (
            O => \N__27083\,
            I => \N__27077\
        );

    \I__2367\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27074\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__27077\,
            I => \b_delay_counter_15__N_4140_adj_4773\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__27074\,
            I => \b_delay_counter_15__N_4140_adj_4773\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__27069\,
            I => \N__27065\
        );

    \I__2363\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27062\
        );

    \I__2362\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27058\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__27062\,
            I => \N__27055\
        );

    \I__2360\ : InMux
    port map (
            O => \N__27061\,
            I => \N__27052\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__27058\,
            I => b_delay_counter_0
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__27055\,
            I => b_delay_counter_0
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__27052\,
            I => b_delay_counter_0
        );

    \I__2356\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27042\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__27042\,
            I => n187
        );

    \I__2354\ : InMux
    port map (
            O => \N__27039\,
            I => \bfn_6_10_0_\
        );

    \I__2353\ : InMux
    port map (
            O => \N__27036\,
            I => \N__27032\
        );

    \I__2352\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27029\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__27032\,
            I => \quad_counter0.b_delay_counter_1\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__27029\,
            I => \quad_counter0.b_delay_counter_1\
        );

    \I__2349\ : InMux
    port map (
            O => \N__27024\,
            I => \quad_counter0.n19656\
        );

    \I__2348\ : InMux
    port map (
            O => \N__27021\,
            I => \quad_counter1.n19686\
        );

    \I__2347\ : InMux
    port map (
            O => \N__27018\,
            I => \quad_counter1.n19687\
        );

    \I__2346\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27011\
        );

    \I__2345\ : InMux
    port map (
            O => \N__27014\,
            I => \N__27008\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__27011\,
            I => \quad_counter1.b_delay_counter_3\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__27008\,
            I => \quad_counter1.b_delay_counter_3\
        );

    \I__2342\ : InMux
    port map (
            O => \N__27003\,
            I => \quad_counter1.n19688\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__27000\,
            I => \N__26996\
        );

    \I__2340\ : InMux
    port map (
            O => \N__26999\,
            I => \N__26993\
        );

    \I__2339\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26990\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__26993\,
            I => \quad_counter1.b_delay_counter_4\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__26990\,
            I => \quad_counter1.b_delay_counter_4\
        );

    \I__2336\ : InMux
    port map (
            O => \N__26985\,
            I => \quad_counter1.n19689\
        );

    \I__2335\ : InMux
    port map (
            O => \N__26982\,
            I => \quad_counter1.n19690\
        );

    \I__2334\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26975\
        );

    \I__2333\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26972\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__26975\,
            I => \quad_counter1.b_delay_counter_6\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__26972\,
            I => \quad_counter1.b_delay_counter_6\
        );

    \I__2330\ : InMux
    port map (
            O => \N__26967\,
            I => \quad_counter1.n19691\
        );

    \I__2329\ : InMux
    port map (
            O => \N__26964\,
            I => \quad_counter1.n19692\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__26961\,
            I => \N__26958\
        );

    \I__2327\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26954\
        );

    \I__2326\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26951\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__26954\,
            I => \N__26948\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__26951\,
            I => \quad_counter1.b_delay_counter_8\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__26948\,
            I => \quad_counter1.b_delay_counter_8\
        );

    \I__2322\ : InMux
    port map (
            O => \N__26943\,
            I => \bfn_5_18_0_\
        );

    \I__2321\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26936\
        );

    \I__2320\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26933\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__26936\,
            I => \N__26930\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__26933\,
            I => \quad_counter1.b_delay_counter_9\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__26930\,
            I => \quad_counter1.b_delay_counter_9\
        );

    \I__2316\ : InMux
    port map (
            O => \N__26925\,
            I => \quad_counter1.n19694\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__26922\,
            I => \quad_counter0.n27_adj_4756_cascade_\
        );

    \I__2314\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__26916\,
            I => \quad_counter0.n25_adj_4757\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__26913\,
            I => \n9809_cascade_\
        );

    \I__2311\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26907\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__2309\ : Odrv12
    port map (
            O => \N__26904\,
            I => n9809
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__26901\,
            I => \quad_counter1.n25_adj_4202_cascade_\
        );

    \I__2307\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__2305\ : Odrv12
    port map (
            O => \N__26892\,
            I => n12940
        );

    \I__2304\ : InMux
    port map (
            O => \N__26889\,
            I => \N__26886\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__26886\,
            I => \N__26883\
        );

    \I__2302\ : Span4Mux_v
    port map (
            O => \N__26883\,
            I => \N__26878\
        );

    \I__2301\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26875\
        );

    \I__2300\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26872\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__26878\,
            I => \N__26866\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__26875\,
            I => \N__26866\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__26872\,
            I => \N__26863\
        );

    \I__2296\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26860\
        );

    \I__2295\ : Span4Mux_v
    port map (
            O => \N__26866\,
            I => \N__26857\
        );

    \I__2294\ : Span12Mux_v
    port map (
            O => \N__26863\,
            I => \N__26852\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__26860\,
            I => \N__26852\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__26857\,
            I => \N__26849\
        );

    \I__2291\ : Span12Mux_v
    port map (
            O => \N__26852\,
            I => \N__26844\
        );

    \I__2290\ : Sp12to4
    port map (
            O => \N__26849\,
            I => \N__26844\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__26844\,
            I => \PIN_13_c\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__26841\,
            I => \n12940_cascade_\
        );

    \I__2287\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26834\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__26837\,
            I => \N__26830\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__26834\,
            I => \N__26827\
        );

    \I__2284\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26824\
        );

    \I__2283\ : InMux
    port map (
            O => \N__26830\,
            I => \N__26821\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__26827\,
            I => \N__26818\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__26824\,
            I => \N__26815\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__26821\,
            I => \quadB_delayed_adj_4768\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__26818\,
            I => \quadB_delayed_adj_4768\
        );

    \I__2278\ : Odrv12
    port map (
            O => \N__26815\,
            I => \quadB_delayed_adj_4768\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__26808\,
            I => \n14425_cascade_\
        );

    \I__2276\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26802\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__26802\,
            I => \quad_counter1.n26_adj_4200\
        );

    \I__2274\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26794\
        );

    \I__2273\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26789\
        );

    \I__2272\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26789\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__26794\,
            I => b_delay_counter_0_adj_4766
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__26789\,
            I => b_delay_counter_0_adj_4766
        );

    \I__2269\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26781\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__26781\,
            I => n187_adj_4771
        );

    \I__2267\ : InMux
    port map (
            O => \N__26778\,
            I => \bfn_5_17_0_\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__26775\,
            I => \quad_counter0.n25_adj_4760_cascade_\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__26772\,
            I => \n12942_cascade_\
        );

    \I__2264\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26766\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__26766\,
            I => \quad_counter0.n28_adj_4754\
        );

    \I__2262\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26760\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__26760\,
            I => \quad_counter0.n26_adj_4755\
        );

    \I__2260\ : IoInMux
    port map (
            O => \N__26757\,
            I => \N__26754\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__26754\,
            I => tx_enable
        );

    \I__2258\ : IoInMux
    port map (
            O => \N__26751\,
            I => \N__26748\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__26748\,
            I => \N__26745\
        );

    \I__2256\ : IoSpan4Mux
    port map (
            O => \N__26745\,
            I => \N__26742\
        );

    \I__2255\ : Span4Mux_s3_v
    port map (
            O => \N__26742\,
            I => \N__26739\
        );

    \I__2254\ : Span4Mux_v
    port map (
            O => \N__26739\,
            I => \N__26736\
        );

    \I__2253\ : Sp12to4
    port map (
            O => \N__26736\,
            I => \N__26732\
        );

    \I__2252\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26729\
        );

    \I__2251\ : Span12Mux_v
    port map (
            O => \N__26732\,
            I => \N__26724\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__26729\,
            I => \N__26724\
        );

    \I__2249\ : Span12Mux_v
    port map (
            O => \N__26724\,
            I => \N__26721\
        );

    \I__2248\ : Odrv12
    port map (
            O => \N__26721\,
            I => \LED_c\
        );

    \I__2247\ : InMux
    port map (
            O => \N__26718\,
            I => \N__26715\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__26715\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__26712\,
            I => \quad_counter0.n22_cascade_\
        );

    \I__2244\ : IoInMux
    port map (
            O => \N__26709\,
            I => \N__26706\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__26706\,
            I => \N__26703\
        );

    \I__2242\ : IoSpan4Mux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__2241\ : IoSpan4Mux
    port map (
            O => \N__26700\,
            I => \N__26697\
        );

    \I__2240\ : IoSpan4Mux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__26694\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19738\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19746\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19754\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19762\,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19770\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19778\,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19786\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19794\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_5_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_17_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19693\,
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19708\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19663\,
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19678\,
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n19730\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_11_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_26_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_19_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_1_0_\
        );

    \IN_MUX_bfv_19_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19625_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_2_0_\
        );

    \IN_MUX_bfv_19_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19626_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_3_0_\
        );

    \IN_MUX_bfv_19_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19627_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_4_0_\
        );

    \IN_MUX_bfv_19_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19628_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_5_0_\
        );

    \IN_MUX_bfv_19_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19629_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_6_0_\
        );

    \IN_MUX_bfv_19_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19630_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_7_0_\
        );

    \IN_MUX_bfv_19_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19631_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_8_0_\
        );

    \IN_MUX_bfv_19_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19632_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_9_0_\
        );

    \IN_MUX_bfv_19_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19633_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_10_0_\
        );

    \IN_MUX_bfv_19_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19634_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_11_0_\
        );

    \IN_MUX_bfv_19_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19635_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_12_0_\
        );

    \IN_MUX_bfv_19_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19636_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_13_0_\
        );

    \IN_MUX_bfv_19_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19637_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_14_0_\
        );

    \IN_MUX_bfv_19_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19638_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_15_0_\
        );

    \IN_MUX_bfv_19_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19639_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_16_0_\
        );

    \IN_MUX_bfv_19_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19640_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_17_0_\
        );

    \IN_MUX_bfv_19_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19641_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_18_0_\
        );

    \IN_MUX_bfv_19_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19642_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_19_0_\
        );

    \IN_MUX_bfv_19_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19643_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_20_0_\
        );

    \IN_MUX_bfv_19_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19644_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_21_0_\
        );

    \IN_MUX_bfv_19_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19645_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_22_0_\
        );

    \IN_MUX_bfv_19_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19646_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_23_0_\
        );

    \IN_MUX_bfv_19_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19647_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_24_0_\
        );

    \IN_MUX_bfv_19_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19648_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_25_0_\
        );

    \IN_MUX_bfv_19_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19649_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_26_0_\
        );

    \IN_MUX_bfv_19_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19650_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_27_0_\
        );

    \IN_MUX_bfv_19_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19651_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_28_0_\
        );

    \IN_MUX_bfv_19_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19652_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_29_0_\
        );

    \IN_MUX_bfv_19_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19653_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_30_0_\
        );

    \IN_MUX_bfv_19_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19654_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_31_0_\
        );

    \IN_MUX_bfv_19_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19655_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_32_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26709\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28592\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_R_49_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26735\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.r_Rx_Data_R\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.quadB_delayed_62_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26871\,
            lcout => \quadB_delayed_adj_4768\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadB_delayed_62_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27411\,
            lcout => \quadB_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.quadB_I_0_79_2_lut_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26833\,
            lcout => \b_delay_counter_15__N_4140_adj_4773\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26718\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__27448\,
            in1 => \N__27045\,
            in2 => \N__27069\,
            in3 => \N__27469\,
            lcout => b_delay_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.B_65_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101000"
        )
    port map (
            in0 => \N__29891\,
            in1 => \N__26882\,
            in2 => \N__26837\,
            in3 => \N__26898\,
            lcout => \B_filtered_adj_4764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i8_4_lut_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27236\,
            in1 => \N__27221\,
            in2 => \N__27204\,
            in3 => \N__27179\,
            lcout => OPEN,
            ltout => \quad_counter0.n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i11_3_lut_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27035\,
            in2 => \N__26712\,
            in3 => \N__27503\,
            lcout => OPEN,
            ltout => \quad_counter0.n25_adj_4760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i2_4_lut_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__27068\,
            in1 => \N__27251\,
            in2 => \N__26775\,
            in3 => \N__27642\,
            lcout => n12942,
            ltout => \n12942_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011011100"
        )
    port map (
            in0 => \N__27417\,
            in1 => \N__27438\,
            in2 => \N__26772\,
            in3 => \N__27368\,
            lcout => n14315,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadB_I_0_79_2_lut_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27412\,
            in2 => \_gnd_net_\,
            in3 => \N__27361\,
            lcout => \b_delay_counter_15__N_4140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i9_4_lut_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__27542\,
            in1 => \N__27734\,
            in2 => \N__27561\,
            in3 => \N__27634\,
            lcout => \quad_counter0.n25_adj_4757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i12_4_lut_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__27575\,
            in1 => \N__27782\,
            in2 => \N__27594\,
            in3 => \N__27608\,
            lcout => \quad_counter0.n28_adj_4754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_delayed_67_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quad_counter0.A_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_delay_counter__i0_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__28007\,
            in1 => \N__27621\,
            in2 => \N__28029\,
            in3 => \N__27635\,
            lcout => a_delay_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i10_4_lut_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27719\,
            in1 => \N__27704\,
            in2 => \N__27528\,
            in3 => \N__27767\,
            lcout => \quad_counter0.n26_adj_4755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i11_4_lut_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27689\,
            in1 => \N__27797\,
            in2 => \N__27753\,
            in3 => \N__28040\,
            lcout => OPEN,
            ltout => \quad_counter0.n27_adj_4756_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i15_4_lut_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26769\,
            in1 => \N__26763\,
            in2 => \N__26922\,
            in3 => \N__26919\,
            lcout => n9809,
            ltout => \n9809_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_2055_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111010"
        )
    port map (
            in0 => \N__27920\,
            in1 => \_gnd_net_\,
            in2 => \N__26913\,
            in3 => \N__27882\,
            lcout => n14469,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_63_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001000000"
        )
    port map (
            in0 => \N__26910\,
            in1 => \N__27909\,
            in2 => \N__27881\,
            in3 => \N__28134\,
            lcout => \A_filtered\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i9_4_lut_adj_1164_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__26940\,
            in1 => \N__27014\,
            in2 => \N__27000\,
            in3 => \N__26797\,
            lcout => OPEN,
            ltout => \quad_counter1.n25_adj_4202_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i15_4_lut_adj_1165_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27930\,
            in1 => \N__26805\,
            in2 => \N__26901\,
            in3 => \N__27804\,
            lcout => n12940,
            ltout => \n12940_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_2054_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26889\,
            in2 => \N__26841\,
            in3 => \N__26838\,
            lcout => n14425,
            ltout => \n14425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.b_delay_counter__i0_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__26798\,
            in1 => \N__26784\,
            in2 => \N__26808\,
            in3 => \N__27082\,
            lcout => b_delay_counter_0_adj_4766,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i10_4_lut_adj_1162_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27144\,
            in1 => \N__27162\,
            in2 => \N__26961\,
            in3 => \N__26978\,
            lcout => \quad_counter1.n26_adj_4200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_86_2_lut_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26799\,
            in2 => \_gnd_net_\,
            in3 => \N__26778\,
            lcout => n187_adj_4771,
            ltout => OPEN,
            carryin => \bfn_5_17_0_\,
            carryout => \quad_counter1.n19686\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.b_delay_counter__i1_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27969\,
            in2 => \_gnd_net_\,
            in3 => \N__27021\,
            lcout => \quad_counter1.b_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter1.n19686\,
            carryout => \quad_counter1.n19687\,
            clk => \N__78563\,
            ce => \N__27114\,
            sr => \N__27095\
        );

    \quad_counter1.b_delay_counter__i2_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27956\,
            in2 => \_gnd_net_\,
            in3 => \N__27018\,
            lcout => \quad_counter1.b_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter1.n19687\,
            carryout => \quad_counter1.n19688\,
            clk => \N__78563\,
            ce => \N__27114\,
            sr => \N__27095\
        );

    \quad_counter1.b_delay_counter__i3_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27015\,
            in2 => \_gnd_net_\,
            in3 => \N__27003\,
            lcout => \quad_counter1.b_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter1.n19688\,
            carryout => \quad_counter1.n19689\,
            clk => \N__78563\,
            ce => \N__27114\,
            sr => \N__27095\
        );

    \quad_counter1.b_delay_counter__i4_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26999\,
            in2 => \_gnd_net_\,
            in3 => \N__26985\,
            lcout => \quad_counter1.b_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter1.n19689\,
            carryout => \quad_counter1.n19690\,
            clk => \N__78563\,
            ce => \N__27114\,
            sr => \N__27095\
        );

    \quad_counter1.b_delay_counter__i5_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27942\,
            in2 => \_gnd_net_\,
            in3 => \N__26982\,
            lcout => \quad_counter1.b_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter1.n19690\,
            carryout => \quad_counter1.n19691\,
            clk => \N__78563\,
            ce => \N__27114\,
            sr => \N__27095\
        );

    \quad_counter1.b_delay_counter__i6_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26979\,
            in2 => \_gnd_net_\,
            in3 => \N__26967\,
            lcout => \quad_counter1.b_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter1.n19691\,
            carryout => \quad_counter1.n19692\,
            clk => \N__78563\,
            ce => \N__27114\,
            sr => \N__27095\
        );

    \quad_counter1.b_delay_counter__i7_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27843\,
            in2 => \_gnd_net_\,
            in3 => \N__26964\,
            lcout => \quad_counter1.b_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter1.n19692\,
            carryout => \quad_counter1.n19693\,
            clk => \N__78563\,
            ce => \N__27114\,
            sr => \N__27095\
        );

    \quad_counter1.b_delay_counter__i8_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26957\,
            in2 => \_gnd_net_\,
            in3 => \N__26943\,
            lcout => \quad_counter1.b_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_5_18_0_\,
            carryout => \quad_counter1.n19694\,
            clk => \N__78566\,
            ce => \N__27113\,
            sr => \N__27096\
        );

    \quad_counter1.b_delay_counter__i9_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26939\,
            in2 => \_gnd_net_\,
            in3 => \N__26925\,
            lcout => \quad_counter1.b_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter1.n19694\,
            carryout => \quad_counter1.n19695\,
            clk => \N__78566\,
            ce => \N__27113\,
            sr => \N__27096\
        );

    \quad_counter1.b_delay_counter__i10_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27161\,
            in2 => \_gnd_net_\,
            in3 => \N__27147\,
            lcout => \quad_counter1.b_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter1.n19695\,
            carryout => \quad_counter1.n19696\,
            clk => \N__78566\,
            ce => \N__27113\,
            sr => \N__27096\
        );

    \quad_counter1.b_delay_counter__i11_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27143\,
            in2 => \_gnd_net_\,
            in3 => \N__27129\,
            lcout => \quad_counter1.b_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter1.n19696\,
            carryout => \quad_counter1.n19697\,
            clk => \N__78566\,
            ce => \N__27113\,
            sr => \N__27096\
        );

    \quad_counter1.b_delay_counter__i12_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27830\,
            in2 => \_gnd_net_\,
            in3 => \N__27126\,
            lcout => \quad_counter1.b_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter1.n19697\,
            carryout => \quad_counter1.n19698\,
            clk => \N__78566\,
            ce => \N__27113\,
            sr => \N__27096\
        );

    \quad_counter1.b_delay_counter__i13_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27983\,
            in2 => \_gnd_net_\,
            in3 => \N__27123\,
            lcout => \quad_counter1.b_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter1.n19698\,
            carryout => \quad_counter1.n19699\,
            clk => \N__78566\,
            ce => \N__27113\,
            sr => \N__27096\
        );

    \quad_counter1.b_delay_counter__i14_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27855\,
            in2 => \_gnd_net_\,
            in3 => \N__27120\,
            lcout => \quad_counter1.b_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter1.n19699\,
            carryout => \quad_counter1.n19700\,
            clk => \N__78566\,
            ce => \N__27113\,
            sr => \N__27096\
        );

    \quad_counter1.b_delay_counter__i15_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27816\,
            in2 => \_gnd_net_\,
            in3 => \N__27117\,
            lcout => \quad_counter1.b_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78566\,
            ce => \N__27113\,
            sr => \N__27096\
        );

    \quad_counter0.add_86_2_lut_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27061\,
            in2 => \_gnd_net_\,
            in3 => \N__27039\,
            lcout => n187,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \quad_counter0.n19656\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27036\,
            in2 => \_gnd_net_\,
            in3 => \N__27024\,
            lcout => \quad_counter0.b_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter0.n19656\,
            carryout => \quad_counter0.n19657\,
            clk => \N__78602\,
            ce => \N__27483\,
            sr => \N__27452\
        );

    \quad_counter0.b_delay_counter__i2_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27252\,
            in2 => \_gnd_net_\,
            in3 => \N__27240\,
            lcout => \quad_counter0.b_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter0.n19657\,
            carryout => \quad_counter0.n19658\,
            clk => \N__78602\,
            ce => \N__27483\,
            sr => \N__27452\
        );

    \quad_counter0.b_delay_counter__i3_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27237\,
            in2 => \_gnd_net_\,
            in3 => \N__27225\,
            lcout => \quad_counter0.b_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter0.n19658\,
            carryout => \quad_counter0.n19659\,
            clk => \N__78602\,
            ce => \N__27483\,
            sr => \N__27452\
        );

    \quad_counter0.b_delay_counter__i4_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27222\,
            in2 => \_gnd_net_\,
            in3 => \N__27210\,
            lcout => \quad_counter0.b_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter0.n19659\,
            carryout => \quad_counter0.n19660\,
            clk => \N__78602\,
            ce => \N__27483\,
            sr => \N__27452\
        );

    \quad_counter0.b_delay_counter__i5_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27278\,
            in2 => \_gnd_net_\,
            in3 => \N__27207\,
            lcout => \quad_counter0.b_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter0.n19660\,
            carryout => \quad_counter0.n19661\,
            clk => \N__78602\,
            ce => \N__27483\,
            sr => \N__27452\
        );

    \quad_counter0.b_delay_counter__i6_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27203\,
            in2 => \_gnd_net_\,
            in3 => \N__27189\,
            lcout => \quad_counter0.b_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter0.n19661\,
            carryout => \quad_counter0.n19662\,
            clk => \N__78602\,
            ce => \N__27483\,
            sr => \N__27452\
        );

    \quad_counter0.b_delay_counter__i7_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27308\,
            in2 => \_gnd_net_\,
            in3 => \N__27186\,
            lcout => \quad_counter0.b_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter0.n19662\,
            carryout => \quad_counter0.n19663\,
            clk => \N__78602\,
            ce => \N__27483\,
            sr => \N__27452\
        );

    \quad_counter0.b_delay_counter__i8_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27327\,
            in2 => \_gnd_net_\,
            in3 => \N__27183\,
            lcout => \quad_counter0.b_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \quad_counter0.n19664\,
            clk => \N__78593\,
            ce => \N__27482\,
            sr => \N__27453\
        );

    \quad_counter0.b_delay_counter__i9_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27180\,
            in2 => \_gnd_net_\,
            in3 => \N__27168\,
            lcout => \quad_counter0.b_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter0.n19664\,
            carryout => \quad_counter0.n19665\,
            clk => \N__78593\,
            ce => \N__27482\,
            sr => \N__27453\
        );

    \quad_counter0.b_delay_counter__i10_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27675\,
            in2 => \_gnd_net_\,
            in3 => \N__27165\,
            lcout => \quad_counter0.b_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter0.n19665\,
            carryout => \quad_counter0.n19666\,
            clk => \N__78593\,
            ce => \N__27482\,
            sr => \N__27453\
        );

    \quad_counter0.b_delay_counter__i11_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27663\,
            in2 => \_gnd_net_\,
            in3 => \N__27510\,
            lcout => \quad_counter0.b_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter0.n19666\,
            carryout => \quad_counter0.n19667\,
            clk => \N__78593\,
            ce => \N__27482\,
            sr => \N__27453\
        );

    \quad_counter0.b_delay_counter__i12_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27294\,
            in2 => \_gnd_net_\,
            in3 => \N__27507\,
            lcout => \quad_counter0.b_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter0.n19667\,
            carryout => \quad_counter0.n19668\,
            clk => \N__78593\,
            ce => \N__27482\,
            sr => \N__27453\
        );

    \quad_counter0.b_delay_counter__i13_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27504\,
            in2 => \_gnd_net_\,
            in3 => \N__27492\,
            lcout => \quad_counter0.b_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter0.n19668\,
            carryout => \quad_counter0.n19669\,
            clk => \N__78593\,
            ce => \N__27482\,
            sr => \N__27453\
        );

    \quad_counter0.b_delay_counter__i14_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27264\,
            in2 => \_gnd_net_\,
            in3 => \N__27489\,
            lcout => \quad_counter0.b_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter0.n19669\,
            carryout => \quad_counter0.n19670\,
            clk => \N__78593\,
            ce => \N__27482\,
            sr => \N__27453\
        );

    \quad_counter0.b_delay_counter__i15_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27339\,
            in2 => \_gnd_net_\,
            in3 => \N__27486\,
            lcout => \quad_counter0.b_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78593\,
            ce => \N__27482\,
            sr => \N__27453\
        );

    \quad_counter0.B_65_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101000"
        )
    port map (
            in0 => \N__27416\,
            in1 => \N__27372\,
            in2 => \N__28092\,
            in3 => \N__27345\,
            lcout => \B_filtered\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i4_2_lut_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27338\,
            in2 => \_gnd_net_\,
            in3 => \N__27326\,
            lcout => \quad_counter0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i3_4_lut_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28064\,
            in1 => \N__28137\,
            in2 => \N__28090\,
            in3 => \N__27315\,
            lcout => count_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i10_4_lut_adj_2052_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27309\,
            in1 => \N__27293\,
            in2 => \N__27282\,
            in3 => \N__27263\,
            lcout => OPEN,
            ltout => \quad_counter0.n24_adj_4758_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i12_4_lut_adj_2053_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27674\,
            in1 => \N__27662\,
            in2 => \N__27651\,
            in3 => \N__27648\,
            lcout => \quad_counter0.n26_adj_4759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_85_2_lut_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27636\,
            in2 => \_gnd_net_\,
            in3 => \N__27612\,
            lcout => n39,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => \quad_counter0.n19671\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_delay_counter__i1_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27609\,
            in2 => \_gnd_net_\,
            in3 => \N__27597\,
            lcout => \quad_counter0.a_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter0.n19671\,
            carryout => \quad_counter0.n19672\,
            clk => \N__78576\,
            ce => \N__28025\,
            sr => \N__28008\
        );

    \quad_counter0.a_delay_counter__i2_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27593\,
            in2 => \_gnd_net_\,
            in3 => \N__27579\,
            lcout => \quad_counter0.a_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter0.n19672\,
            carryout => \quad_counter0.n19673\,
            clk => \N__78576\,
            ce => \N__28025\,
            sr => \N__28008\
        );

    \quad_counter0.a_delay_counter__i3_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27576\,
            in2 => \_gnd_net_\,
            in3 => \N__27564\,
            lcout => \quad_counter0.a_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter0.n19673\,
            carryout => \quad_counter0.n19674\,
            clk => \N__78576\,
            ce => \N__28025\,
            sr => \N__28008\
        );

    \quad_counter0.a_delay_counter__i4_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27560\,
            in2 => \_gnd_net_\,
            in3 => \N__27546\,
            lcout => \quad_counter0.a_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter0.n19674\,
            carryout => \quad_counter0.n19675\,
            clk => \N__78576\,
            ce => \N__28025\,
            sr => \N__28008\
        );

    \quad_counter0.a_delay_counter__i5_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27543\,
            in2 => \_gnd_net_\,
            in3 => \N__27531\,
            lcout => \quad_counter0.a_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter0.n19675\,
            carryout => \quad_counter0.n19676\,
            clk => \N__78576\,
            ce => \N__28025\,
            sr => \N__28008\
        );

    \quad_counter0.a_delay_counter__i6_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27527\,
            in2 => \_gnd_net_\,
            in3 => \N__27513\,
            lcout => \quad_counter0.a_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter0.n19676\,
            carryout => \quad_counter0.n19677\,
            clk => \N__78576\,
            ce => \N__28025\,
            sr => \N__28008\
        );

    \quad_counter0.a_delay_counter__i7_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27798\,
            in2 => \_gnd_net_\,
            in3 => \N__27786\,
            lcout => \quad_counter0.a_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter0.n19677\,
            carryout => \quad_counter0.n19678\,
            clk => \N__78576\,
            ce => \N__28025\,
            sr => \N__28008\
        );

    \quad_counter0.a_delay_counter__i8_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27783\,
            in2 => \_gnd_net_\,
            in3 => \N__27771\,
            lcout => \quad_counter0.a_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => \quad_counter0.n19679\,
            clk => \N__78573\,
            ce => \N__28024\,
            sr => \N__28003\
        );

    \quad_counter0.a_delay_counter__i9_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27768\,
            in2 => \_gnd_net_\,
            in3 => \N__27756\,
            lcout => \quad_counter0.a_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter0.n19679\,
            carryout => \quad_counter0.n19680\,
            clk => \N__78573\,
            ce => \N__28024\,
            sr => \N__28003\
        );

    \quad_counter0.a_delay_counter__i10_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27752\,
            in2 => \_gnd_net_\,
            in3 => \N__27738\,
            lcout => \quad_counter0.a_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter0.n19680\,
            carryout => \quad_counter0.n19681\,
            clk => \N__78573\,
            ce => \N__28024\,
            sr => \N__28003\
        );

    \quad_counter0.a_delay_counter__i11_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27735\,
            in2 => \_gnd_net_\,
            in3 => \N__27723\,
            lcout => \quad_counter0.a_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter0.n19681\,
            carryout => \quad_counter0.n19682\,
            clk => \N__78573\,
            ce => \N__28024\,
            sr => \N__28003\
        );

    \quad_counter0.a_delay_counter__i12_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27720\,
            in2 => \_gnd_net_\,
            in3 => \N__27708\,
            lcout => \quad_counter0.a_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter0.n19682\,
            carryout => \quad_counter0.n19683\,
            clk => \N__78573\,
            ce => \N__28024\,
            sr => \N__28003\
        );

    \quad_counter0.a_delay_counter__i13_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27705\,
            in2 => \_gnd_net_\,
            in3 => \N__27693\,
            lcout => \quad_counter0.a_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter0.n19683\,
            carryout => \quad_counter0.n19684\,
            clk => \N__78573\,
            ce => \N__28024\,
            sr => \N__28003\
        );

    \quad_counter0.a_delay_counter__i14_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27690\,
            in2 => \_gnd_net_\,
            in3 => \N__27678\,
            lcout => \quad_counter0.a_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter0.n19684\,
            carryout => \quad_counter0.n19685\,
            clk => \N__78573\,
            ce => \N__28024\,
            sr => \N__28003\
        );

    \quad_counter0.a_delay_counter__i15_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28041\,
            in2 => \_gnd_net_\,
            in3 => \N__28044\,
            lcout => \quad_counter0.a_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78573\,
            ce => \N__28024\,
            sr => \N__28003\
        );

    \quad_counter0.quadA_I_0_73_2_lut_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27921\,
            in2 => \_gnd_net_\,
            in3 => \N__27871\,
            lcout => \a_delay_counter_15__N_4123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i21282_1_lut_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28951\,
            lcout => \c0.tx.n25051\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i12_4_lut_adj_1161_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__27984\,
            in1 => \N__27968\,
            in2 => \N__27957\,
            in3 => \N__27941\,
            lcout => \quad_counter1.n28_adj_4199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadA_delayed_61_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quadA_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i11_4_lut_adj_1163_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27854\,
            in1 => \N__27842\,
            in2 => \N__27831\,
            in3 => \N__27815\,
            lcout => \quad_counter1.n27_adj_4201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i13_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29494\,
            in2 => \_gnd_net_\,
            in3 => \N__48978\,
            lcout => \c0.FRAME_MATCHER_state_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78568\,
            ce => 'H',
            sr => \N__29472\
        );

    \c0.rx.n25068_bdd_4_lut_4_lut_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000101"
        )
    port map (
            in0 => \N__50825\,
            in1 => \N__39315\,
            in2 => \N__50177\,
            in3 => \N__28284\,
            lcout => n25071,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100011001000"
        )
    port map (
            in0 => \N__28101\,
            in1 => \N__38463\,
            in2 => \N__28686\,
            in3 => \N__28374\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i1074_1_lut_2_lut_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28060\,
            in2 => \_gnd_net_\,
            in3 => \N__28135\,
            lcout => \quad_counter0.n2313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_filtered_I_0_2_lut_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__28136\,
            in1 => \_gnd_net_\,
            in2 => \N__28065\,
            in3 => \_gnd_net_\,
            lcout => \quad_counter0.count_direction\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5179_4_lut_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__29246\,
            in1 => \N__30577\,
            in2 => \N__28449\,
            in3 => \N__28372\,
            lcout => n8628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000100010"
        )
    port map (
            in0 => \N__29247\,
            in1 => \N__28757\,
            in2 => \_gnd_net_\,
            in3 => \N__28539\,
            lcout => \c0.tx.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_4_lut_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28418\,
            in1 => \N__29245\,
            in2 => \N__30582\,
            in3 => \N__28666\,
            lcout => n9603,
            ltout => \n9603_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__28559\,
            in1 => \N__30131\,
            in2 => \N__28095\,
            in3 => \N__28173\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__3__5450_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__47994\,
            in1 => \N__46098\,
            in2 => \N__44781\,
            in3 => \N__28161\,
            lcout => data_out_frame_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5_1_lut_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28410\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n14374,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.B_delayed_68_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28091\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quad_counter0.B_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_2062_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__31197\,
            in1 => \N__28215\,
            in2 => \N__31329\,
            in3 => \N__28611\,
            lcout => n10_adj_4777,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_21318_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__30966\,
            in1 => \N__40816\,
            in2 => \N__30711\,
            in3 => \N__43219\,
            lcout => OPEN,
            ltout => \c0.n25086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n25086_bdd_4_lut_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__40817\,
            in1 => \N__30003\,
            in2 => \N__28164\,
            in3 => \N__28160\,
            lcout => \c0.n25089\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21035_4_lut_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__32151\,
            in1 => \N__31323\,
            in2 => \N__31417\,
            in3 => \N__28197\,
            lcout => OPEN,
            ltout => \n24802_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_2064_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__31324\,
            in1 => \N__31198\,
            in2 => \N__28149\,
            in3 => \N__28143\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29241\,
            in1 => \N__28414\,
            in2 => \N__28683\,
            in3 => \N__28357\,
            lcout => \c0.tx.r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__28508\,
            in1 => \N__28890\,
            in2 => \N__30146\,
            in3 => \N__30213\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30258\,
            in1 => \N__34935\,
            in2 => \_gnd_net_\,
            in3 => \N__43239\,
            lcout => OPEN,
            ltout => \c0.n11_adj_4715_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21242_4_lut_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__40820\,
            in1 => \N__28260\,
            in2 => \N__28146\,
            in3 => \N__41046\,
            lcout => n25010,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_3_lut_3_lut_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__28405\,
            in1 => \N__29240\,
            in2 => \_gnd_net_\,
            in3 => \N__28876\,
            lcout => OPEN,
            ltout => \c0.tx.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i21285_4_lut_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__28406\,
            in1 => \N__28188\,
            in2 => \N__28227\,
            in3 => \N__28206\,
            lcout => \c0.tx.n17199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21249_4_lut_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__28224\,
            in1 => \N__40819\,
            in2 => \N__29154\,
            in3 => \N__41045\,
            lcout => n25018,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__28669\,
            in1 => \N__29239\,
            in2 => \N__29004\,
            in3 => \N__28875\,
            lcout => \c0.tx.n23980\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__28877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29003\,
            lcout => \r_SM_Main_2_N_3751_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30339\,
            in1 => \N__28920\,
            in2 => \_gnd_net_\,
            in3 => \N__43181\,
            lcout => OPEN,
            ltout => \c0.n5_adj_4712_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21033_4_lut_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__28179\,
            in1 => \N__40818\,
            in2 => \N__28200\,
            in3 => \N__41034\,
            lcout => \c0.n24800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13_4_lut_4_lut_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000101"
        )
    port map (
            in0 => \N__50035\,
            in1 => \N__49941\,
            in2 => \N__50178\,
            in3 => \N__42027\,
            lcout => \c0.rx.n14277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_3_lut_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__28998\,
            in1 => \N__29220\,
            in2 => \_gnd_net_\,
            in3 => \N__28667\,
            lcout => \c0.tx.n5_adj_4207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21182_3_lut_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__28251\,
            in1 => \N__41026\,
            in2 => \_gnd_net_\,
            in3 => \N__43171\,
            lcout => \c0.n24949\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i21204_2_lut_4_lut_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__49685\,
            in1 => \N__49656\,
            in2 => \N__47232\,
            in3 => \N__42018\,
            lcout => \c0.rx.n24875\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i14334_2_lut_3_lut_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__28668\,
            in1 => \N__28999\,
            in2 => \_gnd_net_\,
            in3 => \N__28878\,
            lcout => n17951,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1859_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__40780\,
            in1 => \N__31177\,
            in2 => \_gnd_net_\,
            in3 => \N__41025\,
            lcout => n24682,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_21333_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__30240\,
            in1 => \N__40779\,
            in2 => \N__35166\,
            in3 => \N__43180\,
            lcout => OPEN,
            ltout => \c0.n25104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n25104_bdd_4_lut_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__40781\,
            in1 => \N__29109\,
            in2 => \N__28263\,
            in3 => \N__28308\,
            lcout => \c0.n25107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__7__5478_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48067\,
            in1 => \N__46084\,
            in2 => \N__42618\,
            in3 => \N__28250\,
            lcout => data_out_frame_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__28236\,
            in1 => \N__49956\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1940_2_lut_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49658\,
            lcout => OPEN,
            ltout => \n3821_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__49684\,
            in1 => \N__47103\,
            in2 => \N__28230\,
            in3 => \N__47150\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__7__5446_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48068\,
            in1 => \N__45945\,
            in2 => \N__36711\,
            in3 => \N__28307\,
            lcout => data_out_frame_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101000101010"
        )
    port map (
            in0 => \N__50000\,
            in1 => \N__42022\,
            in2 => \N__50162\,
            in3 => \N__28293\,
            lcout => \c0.rx.n25068\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i26_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31585\,
            in2 => \_gnd_net_\,
            in3 => \N__48960\,
            lcout => \c0.FRAME_MATCHER_state_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78595\,
            ce => 'H',
            sr => \N__30495\
        );

    \c0.FRAME_MATCHER_state_i8_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33466\,
            in2 => \_gnd_net_\,
            in3 => \N__48961\,
            lcout => \c0.FRAME_MATCHER_state_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78614\,
            ce => 'H',
            sr => \N__33444\
        );

    \c0.FRAME_MATCHER_state_i14_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29419\,
            in2 => \_gnd_net_\,
            in3 => \N__48962\,
            lcout => \c0.FRAME_MATCHER_state_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78628\,
            ce => 'H',
            sr => \N__29400\
        );

    \quad_counter1.add_85_2_lut_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29700\,
            in2 => \_gnd_net_\,
            in3 => \N__28278\,
            lcout => n39_adj_4770,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \quad_counter1.n19701\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.a_delay_counter__i1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29607\,
            in2 => \_gnd_net_\,
            in3 => \N__28275\,
            lcout => \quad_counter1.a_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter1.n19701\,
            carryout => \quad_counter1.n19702\,
            clk => \N__78686\,
            ce => \N__29789\,
            sr => \N__29777\
        );

    \quad_counter1.a_delay_counter__i2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29594\,
            in2 => \_gnd_net_\,
            in3 => \N__28272\,
            lcout => \quad_counter1.a_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter1.n19702\,
            carryout => \quad_counter1.n19703\,
            clk => \N__78686\,
            ce => \N__29789\,
            sr => \N__29777\
        );

    \quad_counter1.a_delay_counter__i3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29580\,
            in2 => \_gnd_net_\,
            in3 => \N__28269\,
            lcout => \quad_counter1.a_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter1.n19703\,
            carryout => \quad_counter1.n19704\,
            clk => \N__78686\,
            ce => \N__29789\,
            sr => \N__29777\
        );

    \quad_counter1.a_delay_counter__i4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29714\,
            in2 => \_gnd_net_\,
            in3 => \N__28266\,
            lcout => \quad_counter1.a_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter1.n19704\,
            carryout => \quad_counter1.n19705\,
            clk => \N__78686\,
            ce => \N__29789\,
            sr => \N__29777\
        );

    \quad_counter1.a_delay_counter__i5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29739\,
            in2 => \_gnd_net_\,
            in3 => \N__28335\,
            lcout => \quad_counter1.a_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter1.n19705\,
            carryout => \quad_counter1.n19706\,
            clk => \N__78686\,
            ce => \N__29789\,
            sr => \N__29777\
        );

    \quad_counter1.a_delay_counter__i6_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29664\,
            in2 => \_gnd_net_\,
            in3 => \N__28332\,
            lcout => \quad_counter1.a_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter1.n19706\,
            carryout => \quad_counter1.n19707\,
            clk => \N__78686\,
            ce => \N__29789\,
            sr => \N__29777\
        );

    \quad_counter1.a_delay_counter__i7_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29550\,
            in2 => \_gnd_net_\,
            in3 => \N__28329\,
            lcout => \quad_counter1.a_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter1.n19707\,
            carryout => \quad_counter1.n19708\,
            clk => \N__78686\,
            ce => \N__29789\,
            sr => \N__29777\
        );

    \quad_counter1.a_delay_counter__i8_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29619\,
            in2 => \_gnd_net_\,
            in3 => \N__28326\,
            lcout => \quad_counter1.a_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \quad_counter1.n19709\,
            clk => \N__78669\,
            ce => \N__29796\,
            sr => \N__29778\
        );

    \quad_counter1.a_delay_counter__i9_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29676\,
            in2 => \_gnd_net_\,
            in3 => \N__28323\,
            lcout => \quad_counter1.a_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter1.n19709\,
            carryout => \quad_counter1.n19710\,
            clk => \N__78669\,
            ce => \N__29796\,
            sr => \N__29778\
        );

    \quad_counter1.a_delay_counter__i10_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29537\,
            in2 => \_gnd_net_\,
            in3 => \N__28320\,
            lcout => \quad_counter1.a_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter1.n19710\,
            carryout => \quad_counter1.n19711\,
            clk => \N__78669\,
            ce => \N__29796\,
            sr => \N__29778\
        );

    \quad_counter1.a_delay_counter__i11_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29727\,
            in2 => \_gnd_net_\,
            in3 => \N__28317\,
            lcout => \quad_counter1.a_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter1.n19711\,
            carryout => \quad_counter1.n19712\,
            clk => \N__78669\,
            ce => \N__29796\,
            sr => \N__29778\
        );

    \quad_counter1.a_delay_counter__i12_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29651\,
            in2 => \_gnd_net_\,
            in3 => \N__28314\,
            lcout => \quad_counter1.a_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter1.n19712\,
            carryout => \quad_counter1.n19713\,
            clk => \N__78669\,
            ce => \N__29796\,
            sr => \N__29778\
        );

    \quad_counter1.a_delay_counter__i13_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29637\,
            in2 => \_gnd_net_\,
            in3 => \N__28311\,
            lcout => \quad_counter1.a_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter1.n19713\,
            carryout => \quad_counter1.n19714\,
            clk => \N__78669\,
            ce => \N__29796\,
            sr => \N__29778\
        );

    \quad_counter1.a_delay_counter__i14_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29562\,
            in2 => \_gnd_net_\,
            in3 => \N__28428\,
            lcout => \quad_counter1.a_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter1.n19714\,
            carryout => \quad_counter1.n19715\,
            clk => \N__78669\,
            ce => \N__29796\,
            sr => \N__29778\
        );

    \quad_counter1.a_delay_counter__i15_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29523\,
            in2 => \_gnd_net_\,
            in3 => \N__28425\,
            lcout => \quad_counter1.a_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78669\,
            ce => \N__29796\,
            sr => \N__29778\
        );

    \quad_counter1.count_i0_i1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40411\,
            in1 => \N__32367\,
            in2 => \_gnd_net_\,
            in3 => \N__34737\,
            lcout => encoder1_position_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.B_delayed_68_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29906\,
            lcout => \quad_counter1.B_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i5_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40412\,
            in1 => \N__32568\,
            in2 => \_gnd_net_\,
            in3 => \N__41139\,
            lcout => encoder1_position_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78629\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1962_2_lut_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28726\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28774\,
            lcout => \c0.tx.n3843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_adj_1171_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__29242\,
            in1 => \N__28679\,
            in2 => \N__28422\,
            in3 => \N__28373\,
            lcout => \c0.tx.n22949\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000001001000"
        )
    port map (
            in0 => \N__28341\,
            in1 => \N__28545\,
            in2 => \N__28467\,
            in3 => \N__28532\,
            lcout => \c0.tx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011101"
        )
    port map (
            in0 => \N__29244\,
            in1 => \N__28485\,
            in2 => \_gnd_net_\,
            in3 => \N__28685\,
            lcout => OPEN,
            ltout => \n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28574\,
            in1 => \_gnd_net_\,
            in2 => \N__28602\,
            in3 => \N__38471\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__28563\,
            in1 => \N__29970\,
            in2 => \N__28728\,
            in3 => \N__28766\,
            lcout => \c0.tx.n25080\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_3_lut_adj_1172_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__28439\,
            in1 => \N__29243\,
            in2 => \_gnd_net_\,
            in3 => \N__28530\,
            lcout => \c0.tx.n19492\,
            ltout => \c0.tx.n19492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000011000000"
        )
    port map (
            in0 => \N__28531\,
            in1 => \N__28727\,
            in2 => \N__28515\,
            in3 => \N__28767\,
            lcout => \c0.tx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n25080_bdd_4_lut_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__28720\,
            in1 => \N__28512\,
            in2 => \N__30039\,
            in3 => \N__28494\,
            lcout => OPEN,
            ltout => \c0.tx.n25083_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1436221_i1_3_lut_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__28463\,
            in1 => \_gnd_net_\,
            in2 => \N__28488\,
            in3 => \N__28794\,
            lcout => \c0.tx.o_Tx_Serial_N_3782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__30202\,
            in1 => \N__28788\,
            in2 => \N__30138\,
            in3 => \N__28479\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28462\,
            in1 => \N__28722\,
            in2 => \_gnd_net_\,
            in3 => \N__28778\,
            lcout => \c0.tx.n17832\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_2065_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__31328\,
            in1 => \N__31200\,
            in2 => \N__30288\,
            in3 => \N__30351\,
            lcout => OPEN,
            ltout => \n10_adj_4776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__28803\,
            in1 => \N__30203\,
            in2 => \N__28806\,
            in3 => \N__30125\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n25074_bdd_4_lut_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__28721\,
            in1 => \N__28802\,
            in2 => \N__29871\,
            in3 => \N__28692\,
            lcout => \c0.tx.n25077\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0__bdd_4_lut_21308_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011110000"
        )
    port map (
            in0 => \N__28787\,
            in1 => \N__29292\,
            in2 => \N__28779\,
            in3 => \N__28719\,
            lcout => \c0.tx.n25074\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_1174_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28684\,
            in2 => \_gnd_net_\,
            in3 => \N__30581\,
            lcout => \c0.tx.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__2__5483_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48379\,
            in1 => \N__46091\,
            in2 => \N__47316\,
            in3 => \N__29273\,
            lcout => data_out_frame_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21192_3_lut_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__29139\,
            in1 => \N__41009\,
            in2 => \_gnd_net_\,
            in3 => \N__43061\,
            lcout => OPEN,
            ltout => \c0.n24960_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21039_4_lut_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__41010\,
            in1 => \N__32436\,
            in2 => \N__28617\,
            in3 => \N__40811\,
            lcout => OPEN,
            ltout => \c0.n24806_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21041_4_lut_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31271\,
            in1 => \N__31415\,
            in2 => \N__28614\,
            in3 => \N__28902\,
            lcout => n24808,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20990_4_lut_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__29307\,
            in1 => \N__31270\,
            in2 => \N__31419\,
            in3 => \N__34275\,
            lcout => n24757,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__43060\,
            in1 => \_gnd_net_\,
            in2 => \N__37506\,
            in3 => \N__37698\,
            lcout => \c0.n26_adj_4645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_3_lut_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38174\,
            in2 => \_gnd_net_\,
            in3 => \N__38083\,
            lcout => \c0.data_out_frame_29__7__N_1143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_2060_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__28896\,
            in1 => \N__31176\,
            in2 => \N__31304\,
            in3 => \N__29163\,
            lcout => n10_adj_4779,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i2_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40526\,
            in1 => \N__32607\,
            in2 => \_gnd_net_\,
            in3 => \N__46314\,
            lcout => encoder1_position_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__28835\,
            in1 => \N__29066\,
            in2 => \N__29088\,
            in3 => \N__28820\,
            lcout => OPEN,
            ltout => \c0.tx.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i14291_4_lut_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__29051\,
            in1 => \N__29036\,
            in2 => \N__28881\,
            in3 => \N__29021\,
            lcout => \c0.tx.n17904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__28848\,
            in1 => \N__38400\,
            in2 => \_gnd_net_\,
            in3 => \N__28839\,
            lcout => \c0.tx.n24889\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \c0.tx.n19723\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28836\,
            in2 => \_gnd_net_\,
            in3 => \N__28824\,
            lcout => \c0.tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.tx.n19723\,
            carryout => \c0.tx.n19724\,
            clk => \N__78579\,
            ce => \N__38483\,
            sr => \N__28964\
        );

    \c0.tx.r_Clock_Count__i2_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28821\,
            in2 => \_gnd_net_\,
            in3 => \N__28809\,
            lcout => \c0.tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.tx.n19724\,
            carryout => \c0.tx.n19725\,
            clk => \N__78579\,
            ce => \N__38483\,
            sr => \N__28964\
        );

    \c0.tx.r_Clock_Count__i3_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29084\,
            in2 => \_gnd_net_\,
            in3 => \N__29070\,
            lcout => \c0.tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.tx.n19725\,
            carryout => \c0.tx.n19726\,
            clk => \N__78579\,
            ce => \N__38483\,
            sr => \N__28964\
        );

    \c0.tx.r_Clock_Count__i4_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29067\,
            in2 => \_gnd_net_\,
            in3 => \N__29055\,
            lcout => \c0.tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.tx.n19726\,
            carryout => \c0.tx.n19727\,
            clk => \N__78579\,
            ce => \N__38483\,
            sr => \N__28964\
        );

    \c0.tx.r_Clock_Count__i5_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29052\,
            in2 => \_gnd_net_\,
            in3 => \N__29040\,
            lcout => \c0.tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.tx.n19727\,
            carryout => \c0.tx.n19728\,
            clk => \N__78579\,
            ce => \N__38483\,
            sr => \N__28964\
        );

    \c0.tx.r_Clock_Count__i6_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29037\,
            in2 => \_gnd_net_\,
            in3 => \N__29025\,
            lcout => \c0.tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.tx.n19728\,
            carryout => \c0.tx.n19729\,
            clk => \N__78579\,
            ce => \N__38483\,
            sr => \N__28964\
        );

    \c0.tx.r_Clock_Count__i7_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29022\,
            in2 => \_gnd_net_\,
            in3 => \N__29010\,
            lcout => \c0.tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \c0.tx.n19729\,
            carryout => \c0.tx.n19730\,
            clk => \N__78579\,
            ce => \N__38483\,
            sr => \N__28964\
        );

    \c0.tx.r_Clock_Count__i8_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28987\,
            in2 => \_gnd_net_\,
            in3 => \N__29007\,
            lcout => \c0.tx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78570\,
            ce => \N__38484\,
            sr => \N__28965\
        );

    \c0.tx.i2_4_lut_adj_1169_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__28935\,
            in1 => \N__29258\,
            in2 => \N__38478\,
            in3 => \N__29212\,
            lcout => OPEN,
            ltout => \c0.tx.n14290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__29213\,
            in1 => \_gnd_net_\,
            in2 => \N__28923\,
            in3 => \N__30520\,
            lcout => \c0.tx_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__7__5470_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48185\,
            in1 => \N__46089\,
            in2 => \N__44715\,
            in3 => \N__28916\,
            lcout => data_out_frame_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__31095\,
            in1 => \N__29291\,
            in2 => \N__30130\,
            in3 => \N__30217\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001000100"
        )
    port map (
            in0 => \N__41038\,
            in1 => \N__30414\,
            in2 => \N__29277\,
            in3 => \N__43125\,
            lcout => \c0.n6_adj_4649\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__38467\,
            in1 => \N__29259\,
            in2 => \_gnd_net_\,
            in3 => \N__29214\,
            lcout => \r_SM_Main_1_adj_4774\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21238_4_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__38274\,
            in1 => \N__40810\,
            in2 => \N__32454\,
            in3 => \N__41008\,
            lcout => n25006,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29117\,
            in1 => \N__35085\,
            in2 => \_gnd_net_\,
            in3 => \N__43175\,
            lcout => \c0.n11_adj_4663\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__1__5484_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__46085\,
            in1 => \N__48376\,
            in2 => \N__47027\,
            in3 => \N__29135\,
            lcout => data_out_frame_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__3__5418_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__48374\,
            in1 => \N__45505\,
            in2 => \N__29121\,
            in3 => \N__46088\,
            lcout => data_out_frame_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14240_4_lut_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__31157\,
            in1 => \N__29313\,
            in2 => \N__31303\,
            in3 => \N__29319\,
            lcout => \c0.n17846\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__7__5454_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48375\,
            in1 => \N__46087\,
            in2 => \N__29108\,
            in3 => \N__39558\,
            lcout => data_out_frame_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__6__5423_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48373\,
            in1 => \N__46086\,
            in2 => \N__29334\,
            in3 => \N__33702\,
            lcout => data_out_frame_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1472_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33471\,
            in1 => \N__29501\,
            in2 => \N__29433\,
            in3 => \N__49200\,
            lcout => \c0.n14_adj_4520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30018\,
            in1 => \N__43034\,
            in2 => \_gnd_net_\,
            in3 => \N__29330\,
            lcout => \c0.n11_adj_4703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21265_2_lut_3_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__30565\,
            in1 => \N__30526\,
            in2 => \_gnd_net_\,
            in3 => \N__39441\,
            lcout => \c0.tx_transmit_N_3650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__40648\,
            in1 => \N__43032\,
            in2 => \_gnd_net_\,
            in3 => \N__40929\,
            lcout => \c0.n5_adj_4334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1345_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__30072\,
            in1 => \N__29357\,
            in2 => \_gnd_net_\,
            in3 => \N__29375\,
            lcout => \c0.n4_adj_4332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41805\,
            in1 => \N__43033\,
            in2 => \_gnd_net_\,
            in3 => \N__31004\,
            lcout => \c0.n26_adj_4662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1413__i0_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43054\,
            in2 => \N__33215\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \c0.n19795\,
            clk => \N__78605\,
            ce => \N__30471\,
            sr => \N__30462\
        );

    \c0.byte_transmit_counter_1413__i1_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40684\,
            in2 => \_gnd_net_\,
            in3 => \N__29295\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \c0.n19795\,
            carryout => \c0.n19796\,
            clk => \N__78605\,
            ce => \N__30471\,
            sr => \N__30462\
        );

    \c0.byte_transmit_counter_1413__i2_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40995\,
            in2 => \_gnd_net_\,
            in3 => \N__29388\,
            lcout => \c0.byte_transmit_counter_2\,
            ltout => OPEN,
            carryin => \c0.n19796\,
            carryout => \c0.n19797\,
            clk => \N__78605\,
            ce => \N__30471\,
            sr => \N__30462\
        );

    \c0.byte_transmit_counter_1413__i3_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31156\,
            in2 => \_gnd_net_\,
            in3 => \N__29385\,
            lcout => byte_transmit_counter_3,
            ltout => OPEN,
            carryin => \c0.n19797\,
            carryout => \c0.n19798\,
            clk => \N__78605\,
            ce => \N__30471\,
            sr => \N__30462\
        );

    \c0.byte_transmit_counter_1413__i4_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31266\,
            in2 => \_gnd_net_\,
            in3 => \N__29382\,
            lcout => byte_transmit_counter_4,
            ltout => OPEN,
            carryin => \c0.n19798\,
            carryout => \c0.n19799\,
            clk => \N__78605\,
            ce => \N__30471\,
            sr => \N__30462\
        );

    \c0.byte_transmit_counter_1413__i5_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30090\,
            in2 => \_gnd_net_\,
            in3 => \N__29379\,
            lcout => byte_transmit_counter_5,
            ltout => OPEN,
            carryin => \c0.n19799\,
            carryout => \c0.n19800\,
            clk => \N__78605\,
            ce => \N__30471\,
            sr => \N__30462\
        );

    \c0.byte_transmit_counter_1413__i6_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29376\,
            in2 => \_gnd_net_\,
            in3 => \N__29364\,
            lcout => \c0.byte_transmit_counter_6\,
            ltout => OPEN,
            carryin => \c0.n19800\,
            carryout => \c0.n19801\,
            clk => \N__78605\,
            ce => \N__30471\,
            sr => \N__30462\
        );

    \c0.byte_transmit_counter_1413__i7_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29358\,
            in2 => \_gnd_net_\,
            in3 => \N__29361\,
            lcout => \c0.byte_transmit_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78605\,
            ce => \N__30471\,
            sr => \N__30462\
        );

    \c0.FRAME_MATCHER_state_i17_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31559\,
            in2 => \_gnd_net_\,
            in3 => \N__48837\,
            lcout => \c0.FRAME_MATCHER_state_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78616\,
            ce => 'H',
            sr => \N__29457\
        );

    \c0.i1_2_lut_4_lut_adj_1812_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__35784\,
            in1 => \N__44219\,
            in2 => \N__35463\,
            in3 => \N__38951\,
            lcout => \c0.n21611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i3_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35453\,
            in2 => \_gnd_net_\,
            in3 => \N__48825\,
            lcout => \c0.FRAME_MATCHER_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78630\,
            ce => 'H',
            sr => \N__29346\
        );

    \c0.i1_2_lut_4_lut_adj_1845_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__35785\,
            in1 => \N__44220\,
            in2 => \N__33525\,
            in3 => \N__38952\,
            lcout => \c0.n21575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1846_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__35786\,
            in1 => \N__44221\,
            in2 => \N__29505\,
            in3 => \N__38953\,
            lcout => \c0.n21573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1909_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__38954\,
            in1 => \N__31558\,
            in2 => \N__44226\,
            in3 => \N__35787\,
            lcout => \c0.n21581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i9_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33523\,
            in2 => \_gnd_net_\,
            in3 => \N__48838\,
            lcout => \c0.FRAME_MATCHER_state_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78643\,
            ce => 'H',
            sr => \N__29445\
        );

    \c0.i1_2_lut_4_lut_adj_1858_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__35757\,
            in1 => \N__44225\,
            in2 => \N__29429\,
            in3 => \N__38955\,
            lcout => \c0.n21577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i14287_2_lut_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31899\,
            in2 => \_gnd_net_\,
            in3 => \N__31658\,
            lcout => \c0.rx.r_SM_Main_2_N_3680_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i25_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36249\,
            in2 => \_gnd_net_\,
            in3 => \N__48991\,
            lcout => \c0.FRAME_MATCHER_state_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78685\,
            ce => 'H',
            sr => \N__36225\
        );

    \quad_counter1.quadA_delayed_61_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29853\,
            lcout => \quadA_delayed_adj_4767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.quadA_I_0_73_2_lut_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__29852\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29815\,
            lcout => \a_delay_counter_15__N_4123_adj_4772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i15_4_lut_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29625\,
            in1 => \N__29511\,
            in2 => \N__29685\,
            in3 => \N__29568\,
            lcout => n9806,
            ltout => \n9806_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.A_63_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001000"
        )
    port map (
            in0 => \N__29846\,
            in1 => \N__29817\,
            in2 => \N__29856\,
            in3 => \N__30656\,
            lcout => \A_filtered_adj_4763\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__29845\,
            in1 => \N__29816\,
            in2 => \_gnd_net_\,
            in3 => \N__29802\,
            lcout => n14345,
            ltout => \n14345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.a_delay_counter__i0_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__29770\,
            in1 => \N__29699\,
            in2 => \N__29748\,
            in3 => \N__29745\,
            lcout => a_delay_counter_0_adj_4765,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i9_4_lut_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__29738\,
            in1 => \N__29726\,
            in2 => \N__29715\,
            in3 => \N__29698\,
            lcout => \quad_counter1.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i10_4_lut_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29675\,
            in1 => \N__29663\,
            in2 => \N__29652\,
            in3 => \N__29636\,
            lcout => \quad_counter1.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i12_4_lut_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__29618\,
            in1 => \N__29606\,
            in2 => \N__29595\,
            in3 => \N__29579\,
            lcout => \quad_counter1.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i11_4_lut_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29561\,
            in1 => \N__29549\,
            in2 => \N__29538\,
            in3 => \N__29522\,
            lcout => \quad_counter1.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31662\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31917\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78656\,
            ce => 'H',
            sr => \N__49881\
        );

    \CONSTANT_ONE_LUT4_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i3_4_lut_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29877\,
            in1 => \N__30623\,
            in2 => \N__29907\,
            in3 => \N__30658\,
            lcout => count_enable_adj_4769,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.A_delayed_67_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30659\,
            lcout => \quad_counter1.A_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78644\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i1075_1_lut_2_lut_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30622\,
            in2 => \_gnd_net_\,
            in3 => \N__30657\,
            lcout => \quad_counter1.n2226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30732\,
            in1 => \N__45540\,
            in2 => \_gnd_net_\,
            in3 => \N__43222\,
            lcout => \c0.n5_adj_4660\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_2017_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35112\,
            in1 => \N__32140\,
            in2 => \N__41779\,
            in3 => \N__34154\,
            lcout => \c0.data_out_frame_29__7__N_1148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33693\,
            in1 => \N__32201\,
            in2 => \N__33995\,
            in3 => \N__33855\,
            lcout => \c0.n12464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__29870\,
            in1 => \N__29925\,
            in2 => \N__30147\,
            in3 => \N__30201\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1699_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32706\,
            in1 => \N__33854\,
            in2 => \N__33700\,
            in3 => \N__32141\,
            lcout => \c0.n22291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38165\,
            in1 => \N__34609\,
            in2 => \_gnd_net_\,
            in3 => \N__38031\,
            lcout => \c0.n6_adj_4456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1680_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32707\,
            in1 => \N__32200\,
            in2 => \N__33994\,
            in3 => \N__32142\,
            lcout => \c0.n21391\,
            ltout => \c0.n21391_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1529_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38164\,
            in1 => \N__38226\,
            in2 => \N__29916\,
            in3 => \N__38059\,
            lcout => \c0.n12539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1885_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34433\,
            in1 => \N__37287\,
            in2 => \N__35297\,
            in3 => \N__30941\,
            lcout => \c0.n28_adj_4698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i21252_3_lut_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32928\,
            in1 => \N__31199\,
            in2 => \_gnd_net_\,
            in3 => \N__32088\,
            lcout => n25021,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1205_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__38177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38228\,
            lcout => \c0.n21362\,
            ltout => \c0.n21362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1967_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34765\,
            in1 => \N__41364\,
            in2 => \N__29913\,
            in3 => \N__37265\,
            lcout => \c0.n21244\,
            ltout => \c0.n21244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_2006_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37115\,
            in2 => \N__29910\,
            in3 => \N__41413\,
            lcout => \c0.n21309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i25_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40467\,
            in1 => \N__32769\,
            in2 => \_gnd_net_\,
            in3 => \N__35344\,
            lcout => encoder1_position_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1841_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38176\,
            in1 => \N__38227\,
            in2 => \_gnd_net_\,
            in3 => \N__46590\,
            lcout => \c0.n21475\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__4__5297_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38090\,
            in1 => \N__32232\,
            in2 => \N__30810\,
            in3 => \N__46606\,
            lcout => \c0.data_out_frame_28_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78598\,
            ce => \N__45036\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1308_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37939\,
            lcout => \c0.n22163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1272_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35040\,
            in2 => \_gnd_net_\,
            in3 => \N__32345\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1274_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29952\,
            in1 => \N__42147\,
            in2 => \N__29946\,
            in3 => \N__34155\,
            lcout => \c0.n12604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29943\,
            in1 => \N__45075\,
            in2 => \_gnd_net_\,
            in3 => \N__43220\,
            lcout => OPEN,
            ltout => \n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i21253_4_lut_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__31319\,
            in1 => \N__31418\,
            in2 => \N__29937\,
            in3 => \N__29934\,
            lcout => n25022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1765_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37938\,
            in1 => \N__34650\,
            in2 => \_gnd_net_\,
            in3 => \N__36706\,
            lcout => \c0.n22593\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1177_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41430\,
            in2 => \_gnd_net_\,
            in3 => \N__38089\,
            lcout => \c0.n22757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1683_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__38254\,
            in1 => \N__46221\,
            in2 => \N__38189\,
            in3 => \N__32261\,
            lcout => \c0.n22544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1684_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30844\,
            in1 => \N__38178\,
            in2 => \N__38265\,
            in3 => \N__46213\,
            lcout => \c0.n22478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1835_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38179\,
            in1 => \N__50574\,
            in2 => \N__38263\,
            in3 => \N__41495\,
            lcout => \c0.n24033\,
            ltout => \c0.n24033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1476_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38180\,
            in2 => \N__29985\,
            in3 => \N__38025\,
            lcout => n21307,
            ltout => \n21307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32260\,
            in1 => \N__37721\,
            in2 => \N__29982\,
            in3 => \N__50651\,
            lcout => OPEN,
            ltout => \c0.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1184_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32233\,
            in1 => \N__30825\,
            in2 => \N__29979\,
            in3 => \N__29976\,
            lcout => \c0.n22475\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1992_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32259\,
            in1 => \N__46132\,
            in2 => \N__37138\,
            in3 => \N__30772\,
            lcout => \c0.n23918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i13_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50436\,
            in1 => \N__37812\,
            in2 => \_gnd_net_\,
            in3 => \N__37872\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i22_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40485\,
            in1 => \N__32790\,
            in2 => \_gnd_net_\,
            in3 => \N__34649\,
            lcout => encoder1_position_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__2__5475_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__30902\,
            in1 => \N__46083\,
            in2 => \N__37056\,
            in3 => \N__48362\,
            lcout => data_out_frame_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__29966\,
            in1 => \N__30139\,
            in2 => \N__30221\,
            in3 => \N__31038\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1734_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38184\,
            in1 => \N__38010\,
            in2 => \N__40032\,
            in3 => \N__37209\,
            lcout => \c0.n20341\,
            ltout => \c0.n20341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_2031_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__38011\,
            in1 => \N__38262\,
            in2 => \N__30261\,
            in3 => \N__46607\,
            lcout => \c0.n12514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__5__5432_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48348\,
            in1 => \N__46062\,
            in2 => \N__40278\,
            in3 => \N__30308\,
            lcout => data_out_frame_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__7__5414_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__46060\,
            in1 => \N__34595\,
            in2 => \N__48378\,
            in3 => \N__30254\,
            lcout => data_out_frame_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__7__5438_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48347\,
            in1 => \N__46061\,
            in2 => \N__40335\,
            in3 => \N__30236\,
            lcout => data_out_frame_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__30318\,
            in1 => \N__30032\,
            in2 => \N__30222\,
            in3 => \N__30129\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__1__5420_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__48349\,
            in1 => \N__32468\,
            in2 => \N__34785\,
            in3 => \N__46063\,
            lcout => data_out_frame_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__6__5415_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__46059\,
            in1 => \N__34437\,
            in2 => \N__48377\,
            in3 => \N__30017\,
            lcout => data_out_frame_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__3__5458_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48345\,
            in1 => \N__46022\,
            in2 => \N__36564\,
            in3 => \N__29999\,
            lcout => data_out_frame_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21029_4_lut_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__31313\,
            in1 => \N__30786\,
            in2 => \N__31416\,
            in3 => \N__31473\,
            lcout => n24796,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__7__5462_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__46021\,
            in1 => \N__48346\,
            in2 => \N__42720\,
            in3 => \N__30335\,
            lcout => data_out_frame_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101000100"
        )
    port map (
            in0 => \N__40996\,
            in1 => \N__30372\,
            in2 => \N__34860\,
            in3 => \N__43164\,
            lcout => \c0.n6_adj_4659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21038_4_lut_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__31071\,
            in1 => \N__34512\,
            in2 => \N__31318\,
            in3 => \N__31401\,
            lcout => OPEN,
            ltout => \n24805_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__31314\,
            in1 => \N__31158\,
            in2 => \N__30321\,
            in3 => \N__30426\,
            lcout => n10_adj_4780,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_21323_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__38648\,
            in1 => \N__40806\,
            in2 => \N__30312\,
            in3 => \N__43179\,
            lcout => OPEN,
            ltout => \c0.n25092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n25092_bdd_4_lut_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__40807\,
            in1 => \N__35403\,
            in2 => \N__30294\,
            in3 => \N__30269\,
            lcout => OPEN,
            ltout => \c0.n25095_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21246_4_lut_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__41000\,
            in1 => \N__30420\,
            in2 => \N__30291\,
            in3 => \N__40809\,
            lcout => n25014,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__5__5448_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48372\,
            in1 => \N__46026\,
            in2 => \N__30273\,
            in3 => \N__45399\,
            lcout => data_out_frame_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21240_4_lut_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__40808\,
            in1 => \N__30978\,
            in2 => \N__30927\,
            in3 => \N__41001\,
            lcout => n25008,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43178\,
            in1 => \N__35148\,
            in2 => \_gnd_net_\,
            in3 => \N__30387\,
            lcout => \c0.n11_adj_4681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21185_4_lut_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110100000000"
        )
    port map (
            in0 => \N__40949\,
            in1 => \N__30404\,
            in2 => \N__40685\,
            in3 => \N__43053\,
            lcout => \c0.n24953\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21222_2_lut_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40650\,
            in2 => \_gnd_net_\,
            in3 => \N__30395\,
            lcout => \c0.n24897\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__0__5485_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48294\,
            in1 => \N__46025\,
            in2 => \N__45189\,
            in3 => \N__30405\,
            lcout => data_out_frame_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__2__5523_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__33380\,
            in1 => \N__30396\,
            in2 => \N__43838\,
            in3 => \N__43925\,
            lcout => data_out_frame_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__5__5424_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48293\,
            in1 => \N__46024\,
            in2 => \N__32715\,
            in3 => \N__30386\,
            lcout => data_out_frame_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21161_2_lut_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__30359\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40649\,
            lcout => \c0.n24900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1579_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30437\,
            in1 => \N__30456\,
            in2 => \_gnd_net_\,
            in3 => \N__39038\,
            lcout => n14247,
            ltout => \n14247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__3__5522_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011111010"
        )
    port map (
            in0 => \N__30360\,
            in1 => \N__43829\,
            in2 => \N__30363\,
            in3 => \N__43926\,
            lcout => data_out_frame_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1946_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__33600\,
            in1 => \N__35963\,
            in2 => \N__31614\,
            in3 => \N__39111\,
            lcout => OPEN,
            ltout => \c0.n8_adj_4740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19189_4_lut_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__39112\,
            in1 => \N__35826\,
            in2 => \N__30477\,
            in3 => \N__35470\,
            lcout => \c0.n22952\,
            ltout => \c0.n22952_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1960_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30447\,
            in2 => \N__30474\,
            in3 => \N__43533\,
            lcout => \c0.n14380\,
            ltout => \c0.n14380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11327_2_lut_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30465\,
            in3 => \N__44004\,
            lcout => \c0.n14942\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2553_3_lut_4_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__39488\,
            in1 => \N__43830\,
            in2 => \N__48323\,
            in3 => \N__43923\,
            lcout => \c0.n4728\,
            ltout => \c0.n4728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i75_3_lut_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35719\,
            in2 => \N__30450\,
            in3 => \N__44003\,
            lcout => \c0.n58_adj_4742\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_5282_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__35720\,
            in1 => \N__33198\,
            in2 => \N__48324\,
            in3 => \N__39039\,
            lcout => \c0.r_SM_Main_2_N_3754_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78608\,
            ce => 'H',
            sr => \N__30441\
        );

    \c0.rx.i2_4_lut_adj_1167_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__50025\,
            in1 => \N__42007\,
            in2 => \N__50157\,
            in3 => \N__49944\,
            lcout => n14484,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__30555\,
            in1 => \N__30528\,
            in2 => \N__39458\,
            in3 => \N__39144\,
            lcout => \c0.n9_adj_4549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__4__5441_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48271\,
            in1 => \N__46030\,
            in2 => \N__39990\,
            in3 => \N__33254\,
            lcout => data_out_frame_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13932_2_lut_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30554\,
            in2 => \_gnd_net_\,
            in3 => \N__30527\,
            lcout => \c0.n17533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1197_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__39114\,
            in1 => \N__48511\,
            in2 => \N__35691\,
            in3 => \N__30483\,
            lcout => \c0.n5\,
            ltout => \c0.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i22_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30498\,
            in3 => \N__35901\,
            lcout => \c0.FRAME_MATCHER_state_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78632\,
            ce => 'H',
            sr => \N__31605\
        );

    \c0.i1_2_lut_4_lut_adj_1942_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__35780\,
            in1 => \N__44197\,
            in2 => \N__36171\,
            in3 => \N__38944\,
            lcout => \c0.n21595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1943_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__38945\,
            in1 => \N__31593\,
            in2 => \N__44217\,
            in3 => \N__35781\,
            lcout => \c0.n21585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1947_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__35782\,
            in1 => \N__44201\,
            in2 => \N__33610\,
            in3 => \N__38946\,
            lcout => \c0.n21587\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1958_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__38947\,
            in1 => \N__31692\,
            in2 => \N__44218\,
            in3 => \N__35783\,
            lcout => \c0.n21597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_2037_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100000000"
        )
    port map (
            in0 => \N__39451\,
            in1 => \N__39143\,
            in2 => \N__39392\,
            in3 => \N__39113\,
            lcout => \c0.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i30_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31691\,
            in2 => \_gnd_net_\,
            in3 => \N__48824\,
            lcout => \c0.FRAME_MATCHER_state_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78645\,
            ce => 'H',
            sr => \N__30600\
        );

    \c0.FRAME_MATCHER_state_i16_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35545\,
            in2 => \_gnd_net_\,
            in3 => \N__48870\,
            lcout => \c0.FRAME_MATCHER_state_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78655\,
            ce => 'H',
            sr => \N__33633\
        );

    \c0.FRAME_MATCHER_state_i28_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33592\,
            in2 => \_gnd_net_\,
            in3 => \N__48882\,
            lcout => \c0.FRAME_MATCHER_state_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78671\,
            ce => 'H',
            sr => \N__30594\
        );

    \c0.FRAME_MATCHER_state_i23_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49103\,
            in2 => \_gnd_net_\,
            in3 => \N__48984\,
            lcout => \c0.FRAME_MATCHER_state_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78703\,
            ce => 'H',
            sr => \N__31845\
        );

    \c0.i6_4_lut_adj_1385_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32099\,
            in1 => \N__30681\,
            in2 => \N__45613\,
            in3 => \N__39797\,
            lcout => \c0.n14_adj_4368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i4_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47648\,
            in1 => \N__36282\,
            in2 => \_gnd_net_\,
            in3 => \N__45228\,
            lcout => encoder0_position_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78690\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1600_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46357\,
            in1 => \N__45506\,
            in2 => \N__34780\,
            in3 => \N__34610\,
            lcout => \c0.n22218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47647\,
            in1 => \N__36315\,
            in2 => \_gnd_net_\,
            in3 => \N__36349\,
            lcout => encoder0_position_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78690\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1282_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34091\,
            in1 => \N__38809\,
            in2 => \N__33911\,
            in3 => \N__33884\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_2002_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45612\,
            in1 => \N__39549\,
            in2 => \N__30585\,
            in3 => \N__39626\,
            lcout => \c0.n21399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1367_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36788\,
            in2 => \_gnd_net_\,
            in3 => \N__36870\,
            lcout => \c0.n22531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i29_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36843\,
            in1 => \N__47598\,
            in2 => \_gnd_net_\,
            in3 => \N__36871\,
            lcout => encoder0_position_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i13_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40440\,
            in1 => \N__32661\,
            in2 => \_gnd_net_\,
            in3 => \N__32694\,
            lcout => encoder1_position_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i14_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40409\,
            in1 => \N__32643\,
            in2 => \_gnd_net_\,
            in3 => \N__33671\,
            lcout => encoder1_position_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1355_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36801\,
            in2 => \_gnd_net_\,
            in3 => \N__30680\,
            lcout => \c0.n22800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1281_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36489\,
            in1 => \N__30609\,
            in2 => \_gnd_net_\,
            in3 => \N__44409\,
            lcout => \c0.n22611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1352_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36951\,
            in1 => \N__39625\,
            in2 => \_gnd_net_\,
            in3 => \N__44707\,
            lcout => \c0.n13741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1307_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32684\,
            in2 => \_gnd_net_\,
            in3 => \N__32139\,
            lcout => \c0.n22294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1349_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30608\,
            in1 => \N__30743\,
            in2 => \N__38685\,
            in3 => \N__36490\,
            lcout => \c0.n13121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.encoder0_position_27__I_0_2_lut_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__37034\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45598\,
            lcout => \c0.data_out_frame_29__7__N_849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i11_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40410\,
            in1 => \N__32745\,
            in2 => \_gnd_net_\,
            in3 => \N__35116\,
            lcout => encoder1_position_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_2005_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36540\,
            in1 => \N__37033\,
            in2 => \N__42611\,
            in3 => \N__41326\,
            lcout => \c0.n22246\,
            ltout => \c0.n22246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1368_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36488\,
            in1 => \N__42658\,
            in2 => \N__30684\,
            in3 => \N__36597\,
            lcout => \c0.n22846\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i9_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40413\,
            in1 => \N__32523\,
            in2 => \_gnd_net_\,
            in3 => \N__40064\,
            lcout => encoder1_position_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i10_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36598\,
            in1 => \N__47597\,
            in2 => \_gnd_net_\,
            in3 => \N__36579\,
            lcout => encoder0_position_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1306_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43292\,
            in1 => \N__30717\,
            in2 => \_gnd_net_\,
            in3 => \N__43416\,
            lcout => \c0.n20379\,
            ltout => \c0.n20379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1578_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41753\,
            in2 => \N__30666\,
            in3 => \N__32138\,
            lcout => \c0.n13938\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.A_filtered_I_0_2_lut_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__30663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30630\,
            lcout => \quad_counter1.count_direction\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1235_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37116\,
            in2 => \_gnd_net_\,
            in3 => \N__41412\,
            lcout => n21484,
            ltout => \n21484_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1816_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41232\,
            in1 => \N__30753\,
            in2 => \N__30747\,
            in3 => \N__41491\,
            lcout => \c0.n22452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1252_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39982\,
            in1 => \N__34320\,
            in2 => \_gnd_net_\,
            in3 => \N__30744\,
            lcout => \c0.n13384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__0__5469_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48189\,
            in1 => \N__46095\,
            in2 => \N__32502\,
            in3 => \N__36802\,
            lcout => data_out_frame_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__3__5466_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48190\,
            in1 => \N__46096\,
            in2 => \N__42408\,
            in3 => \N__30731\,
            lcout => data_out_frame_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1305_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42818\,
            in1 => \N__42497\,
            in2 => \N__38367\,
            in3 => \N__42263\,
            lcout => \c0.n10_adj_4313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1682_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__38185\,
            in1 => \N__46220\,
            in2 => \N__38264\,
            in3 => \N__50621\,
            lcout => \c0.n22617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__3__5434_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__32853\,
            in1 => \N__30704\,
            in2 => \N__48269\,
            in3 => \N__46097\,
            lcout => data_out_frame_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34263\,
            in1 => \N__38029\,
            in2 => \N__38190\,
            in3 => \N__37605\,
            lcout => \c0.n22668\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1187_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30690\,
            in1 => \N__30759\,
            in2 => \N__41952\,
            in3 => \N__50620\,
            lcout => \c0.n10_adj_4214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1186_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__50588\,
            in1 => \N__34344\,
            in2 => \N__32318\,
            in3 => \N__38092\,
            lcout => \c0.n22534\,
            ltout => \c0.n22534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__2__5299_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30824\,
            in1 => \N__41657\,
            in2 => \N__30831\,
            in3 => \N__30855\,
            lcout => \c0.data_out_frame_28_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78609\,
            ce => \N__45042\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1180_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46883\,
            in2 => \_gnd_net_\,
            in3 => \N__41564\,
            lcout => \c0.n20415\,
            ltout => \c0.n20415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__37137\,
            in1 => \N__41370\,
            in2 => \N__30828\,
            in3 => \N__34367\,
            lcout => \c0.n24530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1661_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30823\,
            in1 => \N__32028\,
            in2 => \N__33996\,
            in3 => \N__32349\,
            lcout => \c0.n22414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1188_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38091\,
            in2 => \_gnd_net_\,
            in3 => \N__46599\,
            lcout => \c0.n20384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__5__5296_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30774\,
            in1 => \N__30809\,
            in2 => \N__46140\,
            in3 => \N__41639\,
            lcout => \c0.data_out_frame_28_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78600\,
            ce => \N__45043\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__43233\,
            in1 => \_gnd_net_\,
            in2 => \N__30795\,
            in3 => \N__34467\,
            lcout => \c0.n26_adj_4680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1633_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37139\,
            in1 => \N__41431\,
            in2 => \_gnd_net_\,
            in3 => \N__30845\,
            lcout => \c0.n21496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1226_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46134\,
            in2 => \_gnd_net_\,
            in3 => \N__30773\,
            lcout => n22735,
            ltout => \n22735_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i21229_4_lut_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30861\,
            in1 => \N__37535\,
            in2 => \N__30876\,
            in3 => \N__34345\,
            lcout => n24904,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1825_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30846\,
            in1 => \N__46135\,
            in2 => \N__30873\,
            in3 => \N__32301\,
            lcout => OPEN,
            ltout => \c0.n20_adj_4699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__0__5293_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50505\,
            in2 => \N__30864\,
            in3 => \N__41850\,
            lcout => \c0.data_out_frame_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78600\,
            ce => \N__45043\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1229_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41562\,
            lcout => n22285,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__47179\,
            in1 => \N__47098\,
            in2 => \_gnd_net_\,
            in3 => \N__47149\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1601_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50650\,
            in1 => \N__38093\,
            in2 => \_gnd_net_\,
            in3 => \N__46608\,
            lcout => \c0.n22330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i7_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40567\,
            in1 => \N__32535\,
            in2 => \_gnd_net_\,
            in3 => \N__34594\,
            lcout => encoder1_position_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_2035_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__41563\,
            in1 => \N__41432\,
            in2 => \_gnd_net_\,
            in3 => \N__38094\,
            lcout => \c0.n6_adj_4210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1808_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__46800\,
            in1 => \N__41366\,
            in2 => \_gnd_net_\,
            in3 => \N__46391\,
            lcout => \c0.n13683\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i15_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40535\,
            in1 => \N__32625\,
            in2 => \_gnd_net_\,
            in3 => \N__34963\,
            lcout => encoder1_position_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__3__5442_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48319\,
            in1 => \N__46056\,
            in2 => \N__34899\,
            in3 => \N__30962\,
            lcout => data_out_frame_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1185_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41230\,
            in1 => \N__41429\,
            in2 => \N__30948\,
            in3 => \N__37742\,
            lcout => \c0.n20641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i3_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32595\,
            in1 => \N__40536\,
            in2 => \_gnd_net_\,
            in3 => \N__45479\,
            lcout => encoder1_position_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__6__5431_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__46055\,
            in1 => \N__48322\,
            in2 => \N__34655\,
            in3 => \N__31532\,
            lcout => data_out_frame_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__2__5459_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48321\,
            in1 => \N__46057\,
            in2 => \N__36622\,
            in3 => \N__31058\,
            lcout => data_out_frame_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33185\,
            in1 => \N__30911\,
            in2 => \_gnd_net_\,
            in3 => \N__43234\,
            lcout => \c0.n11_adj_4572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__0__5421_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__48320\,
            in1 => \N__33953\,
            in2 => \N__30915\,
            in3 => \N__46058\,
            lcout => data_out_frame_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34548\,
            in1 => \N__30903\,
            in2 => \_gnd_net_\,
            in3 => \N__43216\,
            lcout => OPEN,
            ltout => \c0.n5_adj_4650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21042_4_lut_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__40773\,
            in1 => \N__41019\,
            in2 => \N__30888\,
            in3 => \N__30885\,
            lcout => \c0.n24809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21036_4_lut_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__41020\,
            in1 => \N__32487\,
            in2 => \N__31083\,
            in3 => \N__40774\,
            lcout => \c0.n24803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n25056_bdd_4_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__40775\,
            in1 => \N__33342\,
            in2 => \N__31059\,
            in3 => \N__30972\,
            lcout => OPEN,
            ltout => \c0.n25059_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21236_4_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__41021\,
            in1 => \N__32427\,
            in2 => \N__31044\,
            in3 => \N__40776\,
            lcout => OPEN,
            ltout => \n25004_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_2061_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__31189\,
            in1 => \N__31023\,
            in2 => \N__31041\,
            in3 => \N__31317\,
            lcout => n10_adj_4778,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21044_4_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__32409\,
            in1 => \N__31029\,
            in2 => \N__31395\,
            in3 => \N__31312\,
            lcout => n24811,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__3__5298_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__46019\,
            in1 => \N__48252\,
            in2 => \N__31005\,
            in3 => \N__31017\,
            lcout => data_out_frame_28_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_21338_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__33269\,
            in1 => \N__40772\,
            in2 => \N__31446\,
            in3 => \N__43176\,
            lcout => OPEN,
            ltout => \c0.n25110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n25110_bdd_4_lut_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__35226\,
            in1 => \N__34695\,
            in2 => \N__30981\,
            in3 => \N__40805\,
            lcout => \c0.n25113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_21313_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__43177\,
            in1 => \N__31457\,
            in2 => \N__32913\,
            in3 => \N__40804\,
            lcout => \c0.n25056\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__2__5443_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__48250\,
            in1 => \N__31458\,
            in2 => \N__38366\,
            in3 => \N__46020\,
            lcout => data_out_frame_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__0__5437_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__46018\,
            in1 => \N__48251\,
            in2 => \N__34073\,
            in3 => \N__31445\,
            lcout => data_out_frame_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i12_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47653\,
            in1 => \N__36453\,
            in2 => \_gnd_net_\,
            in3 => \N__36487\,
            lcout => encoder0_position_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__5__5480_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__47064\,
            in1 => \N__46023\,
            in2 => \N__31497\,
            in3 => \N__48256\,
            lcout => data_out_frame_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21244_4_lut_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__40778\,
            in1 => \N__31515\,
            in2 => \N__31434\,
            in3 => \N__41023\,
            lcout => n25012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21178_3_lut_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__41022\,
            in1 => \N__34995\,
            in2 => \_gnd_net_\,
            in3 => \N__43217\,
            lcout => OPEN,
            ltout => \c0.n24945_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21030_4_lut_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__40777\,
            in1 => \N__31464\,
            in2 => \N__31422\,
            in3 => \N__41024\,
            lcout => OPEN,
            ltout => \c0.n24797_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21032_4_lut_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31405\,
            in1 => \N__41601\,
            in2 => \N__31332\,
            in3 => \N__31315\,
            lcout => OPEN,
            ltout => \n24799_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_2063_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__31316\,
            in1 => \N__31190\,
            in2 => \N__31104\,
            in3 => \N__31101\,
            lcout => n10_adj_4775,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_21328_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__40769\,
            in1 => \N__35319\,
            in2 => \N__31536\,
            in3 => \N__43085\,
            lcout => OPEN,
            ltout => \c0.n25098_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n25098_bdd_4_lut_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__45699\,
            in1 => \N__33413\,
            in2 => \N__31518\,
            in3 => \N__40771\,
            lcout => \c0.n25101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35385\,
            in1 => \N__31505\,
            in2 => \_gnd_net_\,
            in3 => \N__43084\,
            lcout => \c0.n5_adj_4679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__5__5472_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48363\,
            in1 => \N__45936\,
            in2 => \N__31509\,
            in3 => \N__36897\,
            lcout => data_out_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21247_4_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000100"
        )
    port map (
            in0 => \N__40768\,
            in1 => \N__43087\,
            in2 => \N__41033\,
            in3 => \N__31493\,
            lcout => OPEN,
            ltout => \c0.n25016_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21027_4_lut_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__40994\,
            in1 => \N__31482\,
            in2 => \N__31476\,
            in3 => \N__40770\,
            lcout => \c0.n24794\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43086\,
            in1 => \N__35487\,
            in2 => \_gnd_net_\,
            in3 => \N__33398\,
            lcout => \c0.n5_adj_4700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1849_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__39257\,
            in1 => \N__43825\,
            in2 => \N__43708\,
            in3 => \N__43654\,
            lcout => \c0.n4_adj_4678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i23_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50466\,
            in1 => \N__44499\,
            in2 => \_gnd_net_\,
            in3 => \N__38868\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78633\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i21170_3_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__50044\,
            in1 => \N__31907\,
            in2 => \_gnd_net_\,
            in3 => \N__31654\,
            lcout => n24922,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_105_i4_2_lut_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__49722\,
            in1 => \N__49634\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n4_adj_4761,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1944_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39756\,
            in1 => \N__33552\,
            in2 => \N__36099\,
            in3 => \N__49047\,
            lcout => \c0.n24255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1936_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__35779\,
            in1 => \N__44196\,
            in2 => \N__35908\,
            in3 => \N__38934\,
            lcout => \c0.n21583\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1842_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__44056\,
            in1 => \N__44087\,
            in2 => \N__43997\,
            in3 => \N__43526\,
            lcout => \c0.n13056\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1956_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31592\,
            in2 => \_gnd_net_\,
            in3 => \N__31563\,
            lcout => \c0.n14530\,
            ltout => \c0.n14530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_1964_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35897\,
            in1 => \N__36265\,
            in2 => \N__31539\,
            in3 => \N__36003\,
            lcout => \c0.n6_adj_4495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_2004_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33593\,
            in2 => \_gnd_net_\,
            in3 => \N__33543\,
            lcout => \c0.n14784\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_2_lut_3_lut_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__31976\,
            in1 => \_gnd_net_\,
            in2 => \N__32007\,
            in3 => \N__31900\,
            lcout => OPEN,
            ltout => \c0.rx.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5_4_lut_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__31776\,
            in1 => \N__31953\,
            in2 => \N__31695\,
            in3 => \N__31812\,
            lcout => \c0.rx.r_SM_Main_2_N_3686_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1957_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__36212\,
            in1 => \N__48420\,
            in2 => \_gnd_net_\,
            in3 => \N__31687\,
            lcout => \c0.n22131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_2007_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36170\,
            in2 => \_gnd_net_\,
            in3 => \N__35544\,
            lcout => \c0.n14721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13988_2_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__31749\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31775\,
            lcout => \c0.rx.n17590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13930_2_lut_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31975\,
            in2 => \_gnd_net_\,
            in3 => \N__32003\,
            lcout => OPEN,
            ltout => \c0.rx.n17531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__31722\,
            in1 => \N__31948\,
            in2 => \N__31671\,
            in3 => \N__31668\,
            lcout => \c0.rx.n17848\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5_3_lut_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31949\,
            in1 => \N__31977\,
            in2 => \_gnd_net_\,
            in3 => \N__31805\,
            lcout => \c0.rx.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i20933_3_lut_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__39300\,
            in1 => \N__50865\,
            in2 => \_gnd_net_\,
            in3 => \N__31894\,
            lcout => OPEN,
            ltout => \c0.rx.n24697_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i21217_4_lut_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101010101"
        )
    port map (
            in0 => \N__50042\,
            in1 => \N__31626\,
            in2 => \N__31620\,
            in3 => \N__31818\,
            lcout => OPEN,
            ltout => \c0.rx.n24914_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__50106\,
            in1 => \N__49957\,
            in2 => \N__31617\,
            in3 => \N__42017\,
            lcout => n14895,
            ltout => \n14895_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__31804\,
            in1 => \N__31785\,
            in2 => \N__31833\,
            in3 => \N__39275\,
            lcout => \r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i21223_3_lut_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__39301\,
            in1 => \N__50043\,
            in2 => \_gnd_net_\,
            in3 => \N__50866\,
            lcout => OPEN,
            ltout => \n24921_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000101000101"
        )
    port map (
            in0 => \N__49958\,
            in1 => \N__50107\,
            in2 => \N__31830\,
            in3 => \N__31827\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i21234_4_lut_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__31747\,
            in1 => \N__31773\,
            in2 => \N__31721\,
            in3 => \N__32001\,
            lcout => \c0.rx.n24916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__31803\,
            in1 => \N__31713\,
            in2 => \_gnd_net_\,
            in3 => \N__31746\,
            lcout => \c0.rx.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_2_lut_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31806\,
            in2 => \_gnd_net_\,
            in3 => \N__31779\,
            lcout => n226,
            ltout => OPEN,
            carryin => \bfn_11_26_0_\,
            carryout => \c0.rx.n19716\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i1_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31774\,
            in2 => \_gnd_net_\,
            in3 => \N__31752\,
            lcout => \c0.rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.rx.n19716\,
            carryout => \c0.rx.n19717\,
            clk => \N__78689\,
            ce => \N__39279\,
            sr => \N__31857\
        );

    \c0.rx.r_Clock_Count__i2_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31748\,
            in2 => \_gnd_net_\,
            in3 => \N__31725\,
            lcout => \c0.rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.rx.n19717\,
            carryout => \c0.rx.n19718\,
            clk => \N__78689\,
            ce => \N__39279\,
            sr => \N__31857\
        );

    \c0.rx.r_Clock_Count__i3_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31720\,
            in2 => \_gnd_net_\,
            in3 => \N__32010\,
            lcout => \c0.rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.rx.n19718\,
            carryout => \c0.rx.n19719\,
            clk => \N__78689\,
            ce => \N__39279\,
            sr => \N__31857\
        );

    \c0.rx.r_Clock_Count__i4_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32002\,
            in2 => \_gnd_net_\,
            in3 => \N__31980\,
            lcout => \c0.rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.rx.n19719\,
            carryout => \c0.rx.n19720\,
            clk => \N__78689\,
            ce => \N__39279\,
            sr => \N__31857\
        );

    \c0.rx.r_Clock_Count__i5_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31974\,
            in2 => \_gnd_net_\,
            in3 => \N__31956\,
            lcout => \c0.rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.rx.n19720\,
            carryout => \c0.rx.n19721\,
            clk => \N__78689\,
            ce => \N__39279\,
            sr => \N__31857\
        );

    \c0.rx.r_Clock_Count__i6_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31947\,
            in2 => \_gnd_net_\,
            in3 => \N__31923\,
            lcout => \c0.rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.rx.n19721\,
            carryout => \c0.rx.n19722\,
            clk => \N__78689\,
            ce => \N__39279\,
            sr => \N__31857\
        );

    \c0.rx.r_Clock_Count__i7_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31898\,
            in2 => \_gnd_net_\,
            in3 => \N__31920\,
            lcout => \c0.rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78689\,
            ce => \N__39279\,
            sr => \N__31857\
        );

    \c0.FRAME_MATCHER_state_i4_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36031\,
            in2 => \_gnd_net_\,
            in3 => \N__48992\,
            lcout => \c0.FRAME_MATCHER_state_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78702\,
            ce => 'H',
            sr => \N__33480\
        );

    \c0.i1_2_lut_adj_1986_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49102\,
            in2 => \_gnd_net_\,
            in3 => \N__47836\,
            lcout => \c0.n21645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1351_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36421\,
            in2 => \_gnd_net_\,
            in3 => \N__36341\,
            lcout => \c0.n22638\,
            ltout => \c0.n22638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1760_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36964\,
            in1 => \N__39613\,
            in2 => \N__31836\,
            in3 => \N__44708\,
            lcout => \c0.n6_adj_4336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1254_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__33891\,
            in1 => \N__33869\,
            in2 => \_gnd_net_\,
            in3 => \N__34028\,
            lcout => \c0.n20333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.encoder0_position_29__I_0_2_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__36874\,
            in1 => \_gnd_net_\,
            in2 => \N__36975\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_frame_29__7__N_855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1404_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34011\,
            in1 => \N__33852\,
            in2 => \_gnd_net_\,
            in3 => \N__42330\,
            lcout => \c0.n21323\,
            ltout => \c0.n21323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1266_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__34746\,
            in1 => \_gnd_net_\,
            in2 => \N__32052\,
            in3 => \N__38122\,
            lcout => \c0.n21406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1314_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32848\,
            in1 => \N__36342\,
            in2 => \_gnd_net_\,
            in3 => \N__36872\,
            lcout => \c0.n22608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1386_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44382\,
            in1 => \N__37899\,
            in2 => \N__36974\,
            in3 => \N__32049\,
            lcout => \c0.n12488\,
            ltout => \c0.n12488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1750_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__45591\,
            in1 => \_gnd_net_\,
            in2 => \N__32043\,
            in3 => \N__36873\,
            lcout => \c0.n20449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1354_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35188\,
            in2 => \_gnd_net_\,
            in3 => \N__36422\,
            lcout => \c0.n22791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_2015_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35111\,
            in1 => \N__32040\,
            in2 => \_gnd_net_\,
            in3 => \N__34136\,
            lcout => \c0.n13531\,
            ltout => \c0.n13531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1332_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41752\,
            in1 => \N__38551\,
            in2 => \N__32031\,
            in3 => \N__32021\,
            lcout => \c0.n29_adj_4329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1322_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36697\,
            in1 => \N__35353\,
            in2 => \_gnd_net_\,
            in3 => \N__42552\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4317_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1324_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44349\,
            in1 => \N__32073\,
            in2 => \N__32067\,
            in3 => \N__32064\,
            lcout => \c0.n20388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1323_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34181\,
            in1 => \N__39553\,
            in2 => \N__42174\,
            in3 => \N__34027\,
            lcout => \c0.n15_adj_4318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1334_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38552\,
            lcout => \c0.n6_adj_4330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1335_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39915\,
            in1 => \N__32058\,
            in2 => \N__44432\,
            in3 => \N__42400\,
            lcout => \c0.n20348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_2010_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39875\,
            in1 => \N__37035\,
            in2 => \_gnd_net_\,
            in3 => \N__41318\,
            lcout => \c0.n20_adj_4321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i19_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32847\,
            in1 => \N__32820\,
            in2 => \_gnd_net_\,
            in3 => \N__40528\,
            lcout => encoder1_position_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i11_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47654\,
            in1 => \N__36522\,
            in2 => \_gnd_net_\,
            in3 => \N__36547\,
            lcout => encoder0_position_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i28_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36957\,
            in1 => \N__36912\,
            in2 => \_gnd_net_\,
            in3 => \N__47656\,
            lcout => encoder0_position_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i12_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40527\,
            in1 => \N__32730\,
            in2 => \_gnd_net_\,
            in3 => \N__41760\,
            lcout => encoder1_position_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i26_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__37008\,
            in1 => \_gnd_net_\,
            in2 => \N__37045\,
            in3 => \N__47655\,
            lcout => encoder0_position_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i4_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32580\,
            in1 => \N__40543\,
            in2 => \_gnd_net_\,
            in3 => \N__35268\,
            lcout => encoder1_position_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1303_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34895\,
            in1 => \N__34316\,
            in2 => \_gnd_net_\,
            in3 => \N__42498\,
            lcout => \c0.n20367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1353_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32112\,
            in1 => \N__47485\,
            in2 => \N__32889\,
            in3 => \N__32103\,
            lcout => \c0.n13395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n25062_bdd_4_lut_4_lut_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011000"
        )
    port map (
            in0 => \N__41053\,
            in1 => \N__40599\,
            in2 => \N__33369\,
            in3 => \N__43238\,
            lcout => n25065,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i6_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40541\,
            in1 => \N__32550\,
            in2 => \_gnd_net_\,
            in3 => \N__34421\,
            lcout => encoder1_position_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i20_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40542\,
            in1 => \N__32805\,
            in2 => \_gnd_net_\,
            in3 => \N__33798\,
            lcout => encoder1_position_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40540\,
            in1 => \N__32382\,
            in2 => \_gnd_net_\,
            in3 => \N__33942\,
            lcout => encoder1_position_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1524_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44626\,
            in1 => \N__35261\,
            in2 => \N__41172\,
            in3 => \N__34814\,
            lcout => \c0.n10500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_4_lut_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34815\,
            in1 => \N__46877\,
            in2 => \N__35283\,
            in3 => \N__44627\,
            lcout => \c0.n9_adj_4562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1811_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32234\,
            in1 => \N__32344\,
            in2 => \N__32319\,
            in3 => \N__32274\,
            lcout => \c0.n12_adj_4688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1815_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32297\,
            in1 => \N__46696\,
            in2 => \N__46395\,
            in3 => \N__34449\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4690_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1814_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32286\,
            in1 => \N__34352\,
            in2 => \N__32277\,
            in3 => \N__37091\,
            lcout => \c0.n22710\,
            ltout => \c0.n22710_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1793_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32268\,
            in3 => \N__32265\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4683_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__6__5287_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32235\,
            in1 => \N__37779\,
            in2 => \N__32208\,
            in3 => \N__32175\,
            lcout => \c0.data_out_frame_29_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78634\,
            ce => \N__45054\,
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1810_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32168\,
            in1 => \N__46557\,
            in2 => \N__32205\,
            in3 => \N__32181\,
            lcout => \c0.n20360\,
            ltout => \c0.n20360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__7__5286_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32169\,
            in2 => \N__32160\,
            in3 => \N__38030\,
            lcout => \c0.data_out_frame_29_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78622\,
            ce => \N__45035\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43231\,
            in1 => \N__32157\,
            in2 => \_gnd_net_\,
            in3 => \N__41472\,
            lcout => \c0.n26_adj_4713\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33234\,
            in1 => \N__32498\,
            in2 => \_gnd_net_\,
            in3 => \N__43229\,
            lcout => \c0.n5_adj_4567\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43227\,
            in1 => \N__32475\,
            in2 => \_gnd_net_\,
            in3 => \N__33171\,
            lcout => \c0.n11_adj_4646\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34842\,
            in1 => \N__41283\,
            in2 => \_gnd_net_\,
            in3 => \N__43230\,
            lcout => \c0.n5_adj_4644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__43232\,
            in1 => \_gnd_net_\,
            in2 => \N__35064\,
            in3 => \N__33315\,
            lcout => \c0.n11_adj_4652\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41262\,
            in1 => \N__32415\,
            in2 => \_gnd_net_\,
            in3 => \N__43228\,
            lcout => \c0.n26_adj_4651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_1_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32995\,
            in2 => \N__33074\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \quad_counter1.n19731\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_2_lut_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33946\,
            in2 => \N__32394\,
            in3 => \N__32370\,
            lcout => n2291,
            ltout => OPEN,
            carryin => \quad_counter1.n19731\,
            carryout => \quad_counter1.n19732\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_3_lut_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34775\,
            in2 => \N__33075\,
            in3 => \N__32352\,
            lcout => n2290,
            ltout => OPEN,
            carryin => \quad_counter1.n19732\,
            carryout => \quad_counter1.n19733\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_4_lut_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46329\,
            in2 => \N__33071\,
            in3 => \N__32598\,
            lcout => n2289,
            ltout => OPEN,
            carryin => \quad_counter1.n19733\,
            carryout => \quad_counter1.n19734\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_5_lut_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45493\,
            in2 => \N__33076\,
            in3 => \N__32583\,
            lcout => n2288,
            ltout => OPEN,
            carryin => \quad_counter1.n19734\,
            carryout => \quad_counter1.n19735\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_6_lut_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35284\,
            in2 => \N__33072\,
            in3 => \N__32571\,
            lcout => n2287,
            ltout => OPEN,
            carryin => \quad_counter1.n19735\,
            carryout => \quad_counter1.n19736\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_7_lut_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41185\,
            in2 => \N__33077\,
            in3 => \N__32553\,
            lcout => n2286,
            ltout => OPEN,
            carryin => \quad_counter1.n19736\,
            carryout => \quad_counter1.n19737\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_8_lut_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34425\,
            in2 => \N__33073\,
            in3 => \N__32538\,
            lcout => n2285,
            ltout => OPEN,
            carryin => \quad_counter1.n19737\,
            carryout => \quad_counter1.n19738\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_9_lut_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34593\,
            in2 => \N__33129\,
            in3 => \N__32529\,
            lcout => n2284,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \quad_counter1.n19739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_10_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33081\,
            in2 => \N__40174\,
            in3 => \N__32526\,
            lcout => n2283,
            ltout => OPEN,
            carryin => \quad_counter1.n19739\,
            carryout => \quad_counter1.n19740\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_11_lut_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40084\,
            in2 => \N__33130\,
            in3 => \N__32508\,
            lcout => n2282,
            ltout => OPEN,
            carryin => \quad_counter1.n19740\,
            carryout => \quad_counter1.n19741\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_12_lut_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33085\,
            in2 => \N__35038\,
            in3 => \N__32505\,
            lcout => n2281,
            ltout => OPEN,
            carryin => \quad_counter1.n19741\,
            carryout => \quad_counter1.n19742\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_13_lut_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35132\,
            in2 => \N__33131\,
            in3 => \N__32733\,
            lcout => n2280,
            ltout => OPEN,
            carryin => \quad_counter1.n19742\,
            carryout => \quad_counter1.n19743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_14_lut_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33089\,
            in2 => \N__41780\,
            in3 => \N__32718\,
            lcout => n2279,
            ltout => OPEN,
            carryin => \quad_counter1.n19743\,
            carryout => \quad_counter1.n19744\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_15_lut_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32711\,
            in2 => \N__33132\,
            in3 => \N__32646\,
            lcout => n2278,
            ltout => OPEN,
            carryin => \quad_counter1.n19744\,
            carryout => \quad_counter1.n19745\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_16_lut_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33093\,
            in2 => \N__33701\,
            in3 => \N__32628\,
            lcout => n2277,
            ltout => OPEN,
            carryin => \quad_counter1.n19745\,
            carryout => \quad_counter1.n19746\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_17_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34959\,
            in2 => \N__33133\,
            in3 => \N__32619\,
            lcout => n2276,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \quad_counter1.n19747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_18_lut_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33097\,
            in2 => \N__34083\,
            in3 => \N__32616\,
            lcout => n2275,
            ltout => OPEN,
            carryin => \quad_counter1.n19747\,
            carryout => \quad_counter1.n19748\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_19_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35207\,
            in2 => \N__33134\,
            in3 => \N__32613\,
            lcout => n2274,
            ltout => OPEN,
            carryin => \quad_counter1.n19748\,
            carryout => \quad_counter1.n19749\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_20_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33101\,
            in2 => \N__32888\,
            in3 => \N__32610\,
            lcout => n2273,
            ltout => OPEN,
            carryin => \quad_counter1.n19749\,
            carryout => \quad_counter1.n19750\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_21_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32849\,
            in2 => \N__33135\,
            in3 => \N__32808\,
            lcout => n2272,
            ltout => OPEN,
            carryin => \quad_counter1.n19750\,
            carryout => \quad_counter1.n19751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_22_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33105\,
            in2 => \N__33806\,
            in3 => \N__32796\,
            lcout => n2271,
            ltout => OPEN,
            carryin => \quad_counter1.n19751\,
            carryout => \quad_counter1.n19752\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_23_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40264\,
            in2 => \N__33136\,
            in3 => \N__32793\,
            lcout => n2270,
            ltout => OPEN,
            carryin => \quad_counter1.n19752\,
            carryout => \quad_counter1.n19753\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_24_lut_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33109\,
            in2 => \N__34659\,
            in3 => \N__32778\,
            lcout => n2269,
            ltout => OPEN,
            carryin => \quad_counter1.n19753\,
            carryout => \quad_counter1.n19754\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_25_lut_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38542\,
            in2 => \N__33137\,
            in3 => \N__32775\,
            lcout => n2268,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \quad_counter1.n19755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_26_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33113\,
            in2 => \N__37946\,
            in3 => \N__32772\,
            lcout => n2267,
            ltout => OPEN,
            carryin => \quad_counter1.n19755\,
            carryout => \quad_counter1.n19756\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_27_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35360\,
            in2 => \N__33138\,
            in3 => \N__32754\,
            lcout => n2266,
            ltout => OPEN,
            carryin => \quad_counter1.n19756\,
            carryout => \quad_counter1.n19757\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_28_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33117\,
            in2 => \N__38365\,
            in3 => \N__32751\,
            lcout => n2265,
            ltout => OPEN,
            carryin => \quad_counter1.n19757\,
            carryout => \quad_counter1.n19758\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_29_lut_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34884\,
            in2 => \N__33139\,
            in3 => \N__32748\,
            lcout => n2264,
            ltout => OPEN,
            carryin => \quad_counter1.n19758\,
            carryout => \quad_counter1.n19759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_30_lut_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33121\,
            in2 => \N__39972\,
            in3 => \N__33150\,
            lcout => n2263,
            ltout => OPEN,
            carryin => \quad_counter1.n19759\,
            carryout => \quad_counter1.n19760\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_31_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38673\,
            in2 => \N__33140\,
            in3 => \N__33147\,
            lcout => n2262,
            ltout => OPEN,
            carryin => \quad_counter1.n19760\,
            carryout => \quad_counter1.n19761\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_32_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33125\,
            in2 => \N__38811\,
            in3 => \N__33144\,
            lcout => n2261,
            ltout => OPEN,
            carryin => \quad_counter1.n19761\,
            carryout => \quad_counter1.n19762\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_613_33_lut_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40331\,
            in1 => \N__33141\,
            in2 => \_gnd_net_\,
            in3 => \N__32934\,
            lcout => n2260,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__1__5452_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__38288\,
            in1 => \N__48249\,
            in2 => \N__36363\,
            in3 => \N__45991\,
            lcout => data_out_frame_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21017_4_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__41017\,
            in1 => \N__35409\,
            in2 => \N__40815\,
            in3 => \N__33240\,
            lcout => OPEN,
            ltout => \c0.n24784_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21250_4_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__42891\,
            in1 => \N__40767\,
            in2 => \N__32931\,
            in3 => \N__41018\,
            lcout => n25019,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__2__5435_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__45989\,
            in1 => \N__32912\,
            in2 => \N__32884\,
            in3 => \N__48248\,
            lcout => data_out_frame_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i18_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32898\,
            in1 => \N__32877\,
            in2 => \_gnd_net_\,
            in3 => \N__40545\,
            lcout => encoder1_position_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i16_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40544\,
            in1 => \N__33282\,
            in2 => \_gnd_net_\,
            in3 => \N__34074\,
            lcout => encoder1_position_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__0__5445_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48247\,
            in1 => \N__45990\,
            in2 => \N__37950\,
            in3 => \N__33270\,
            lcout => data_out_frame_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14062_2_lut_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43796\,
            in2 => \_gnd_net_\,
            in3 => \N__43901\,
            lcout => \c0.data_out_frame_29_7_N_1482_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21016_3_lut_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43206\,
            in1 => \N__33326\,
            in2 => \_gnd_net_\,
            in3 => \N__33258\,
            lcout => \c0.n24783\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__0__5477_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45882\,
            in1 => \N__48255\,
            in2 => \N__42567\,
            in3 => \N__33233\,
            lcout => data_out_frame_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21165_4_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010100010"
        )
    port map (
            in0 => \N__43516\,
            in1 => \N__43998\,
            in2 => \N__33219\,
            in3 => \N__39495\,
            lcout => \c0.n24888\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__0__5429_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45880\,
            in1 => \N__48253\,
            in2 => \N__40179\,
            in3 => \N__33186\,
            lcout => data_out_frame_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i19_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50391\,
            in1 => \N__38718\,
            in2 => \_gnd_net_\,
            in3 => \N__43329\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__1__5428_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45881\,
            in1 => \N__48254\,
            in2 => \N__40098\,
            in3 => \N__33164\,
            lcout => data_out_frame_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__6__5447_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45873\,
            in1 => \N__48246\,
            in2 => \N__42789\,
            in3 => \N__33414\,
            lcout => data_out_frame_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__6__5471_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48243\,
            in1 => \N__45875\,
            in2 => \N__39645\,
            in3 => \N__33399\,
            lcout => data_out_frame_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__4__5521_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011111010"
        )
    port map (
            in0 => \N__33387\,
            in1 => \N__43824\,
            in2 => \N__33362\,
            in3 => \N__43911\,
            lcout => data_out_frame_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__2__5451_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45872\,
            in1 => \N__48245\,
            in2 => \N__39861\,
            in3 => \N__33341\,
            lcout => data_out_frame_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__4__5433_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48242\,
            in1 => \N__45874\,
            in2 => \N__33810\,
            in3 => \N__33327\,
            lcout => data_out_frame_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__2__5419_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__45871\,
            in1 => \N__48244\,
            in2 => \N__33311\,
            in3 => \N__46356\,
            lcout => data_out_frame_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1985_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__35964\,
            in1 => \N__33291\,
            in2 => \N__43431\,
            in3 => \N__39110\,
            lcout => \c0.n4_adj_4212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1687_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43491\,
            in2 => \_gnd_net_\,
            in3 => \N__39412\,
            lcout => \c0.n12976\,
            ltout => \c0.n12976_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1237_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__35982\,
            in1 => \N__39089\,
            in2 => \N__33285\,
            in3 => \N__48443\,
            lcout => \c0.n63_adj_4249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1175_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36213\,
            in2 => \_gnd_net_\,
            in3 => \N__47787\,
            lcout => \c0.n21649\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1972_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__43968\,
            in1 => \N__44086\,
            in2 => \_gnd_net_\,
            in3 => \N__44262\,
            lcout => \c0.n58_adj_4706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14178_2_lut_3_lut_4_lut_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__35616\,
            in1 => \N__43816\,
            in2 => \N__44142\,
            in3 => \N__35664\,
            lcout => \c0.data_out_frame_29_7_N_1482_0\,
            ltout => \c0.data_out_frame_29_7_N_1482_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1725_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__33612\,
            in1 => \N__39088\,
            in2 => \N__33435\,
            in3 => \N__33551\,
            lcout => \c0.n13052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i15_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44548\,
            in1 => \N__50453\,
            in2 => \_gnd_net_\,
            in3 => \N__38875\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1670_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__35614\,
            in1 => \_gnd_net_\,
            in2 => \N__43834\,
            in3 => \N__35662\,
            lcout => \c0.n9706\,
            ltout => \c0.n9706_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14180_4_lut_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__33432\,
            in1 => \N__33426\,
            in2 => \N__33420\,
            in3 => \N__49043\,
            lcout => \c0.n9248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1545_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__35615\,
            in1 => \N__43698\,
            in2 => \N__43835\,
            in3 => \N__35663\,
            lcout => \c0.n9587\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1771_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__49793\,
            in1 => \N__33620\,
            in2 => \N__35814\,
            in3 => \N__38913\,
            lcout => \c0.n6\,
            ltout => \c0.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1916_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33501\,
            in2 => \N__33417\,
            in3 => \_gnd_net_\,
            lcout => \c0.n21625\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1868_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__35756\,
            in1 => \N__44195\,
            in2 => \N__35562\,
            in3 => \N__38914\,
            lcout => \c0.n21579\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1772_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__33621\,
            in1 => \N__35813\,
            in2 => \_gnd_net_\,
            in3 => \N__49794\,
            lcout => \c0.n17682\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19210_3_lut_4_lut_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__35975\,
            in1 => \N__39071\,
            in2 => \N__33611\,
            in3 => \N__33544\,
            lcout => \c0.n22907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1474_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33524\,
            in1 => \N__39202\,
            in2 => \N__39705\,
            in3 => \N__33499\,
            lcout => \c0.n9_adj_4522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i5_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33500\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48941\,
            lcout => \c0.FRAME_MATCHER_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78674\,
            ce => 'H',
            sr => \N__33486\
        );

    \c0.i1_2_lut_adj_1912_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36041\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47788\,
            lcout => \c0.n8_adj_4561\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1922_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47789\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36080\,
            lcout => \c0.n21637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1934_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47790\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33470\,
            lcout => \c0.n8_adj_4558\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i10_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39206\,
            in2 => \_gnd_net_\,
            in3 => \N__48928\,
            lcout => \c0.FRAME_MATCHER_state_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78691\,
            ce => 'H',
            sr => \N__39186\
        );

    \c0.FRAME_MATCHER_state_i6_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36076\,
            in2 => \_gnd_net_\,
            in3 => \N__48969\,
            lcout => \c0.FRAME_MATCHER_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78704\,
            ce => 'H',
            sr => \N__33759\
        );

    \c0.i2_3_lut_adj_1387_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36976\,
            in1 => \N__45602\,
            in2 => \_gnd_net_\,
            in3 => \N__33717\,
            lcout => OPEN,
            ltout => \c0.n22831_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1325_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33747\,
            in1 => \N__42307\,
            in2 => \N__33741\,
            in3 => \N__36688\,
            lcout => \c0.n14_adj_4319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1326_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45229\,
            in1 => \N__39835\,
            in2 => \N__44762\,
            in3 => \N__39914\,
            lcout => OPEN,
            ltout => \c0.n13_adj_4320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1327_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33738\,
            in1 => \N__42822\,
            in2 => \N__33729\,
            in3 => \N__33726\,
            lcout => OPEN,
            ltout => \c0.n28_adj_4322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1331_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34090\,
            in1 => \N__40266\,
            in2 => \N__33720\,
            in3 => \N__39927\,
            lcout => \c0.n34_adj_4328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1751_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40324\,
            in1 => \N__47497\,
            in2 => \_gnd_net_\,
            in3 => \N__33715\,
            lcout => \c0.n22656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1359_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__33716\,
            in1 => \_gnd_net_\,
            in2 => \N__47502\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n20318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1309_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33686\,
            in1 => \N__34976\,
            in2 => \N__33636\,
            in3 => \N__38810\,
            lcout => \c0.n22466\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1392_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34977\,
            in1 => \N__34205\,
            in2 => \N__34098\,
            in3 => \N__34029\,
            lcout => \c0.n10_adj_4374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21196_2_lut_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34677\,
            in2 => \_gnd_net_\,
            in3 => \N__43182\,
            lcout => \c0.n24901\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1253_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34002\,
            in1 => \N__33993\,
            in2 => \N__33954\,
            in3 => \N__33915\,
            lcout => \c0.n10_adj_4274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i16_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__36753\,
            in1 => \N__47726\,
            in2 => \N__36803\,
            in3 => \_gnd_net_\,
            lcout => encoder0_position_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78705\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_1758_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47312\,
            in1 => \N__44862\,
            in2 => \N__33885\,
            in3 => \N__47028\,
            lcout => \c0.n10_adj_4339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1329_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40127\,
            in1 => \N__33870\,
            in2 => \N__33771\,
            in3 => \N__45437\,
            lcout => OPEN,
            ltout => \c0.n30_adj_4326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1333_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33853\,
            in1 => \N__33828\,
            in2 => \N__33819\,
            in3 => \N__33816\,
            lcout => \c0.n22408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1310_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__33799\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39623\,
            lcout => \c0.n22788\,
            ltout => \c0.n22788_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1297_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44861\,
            in1 => \N__39841\,
            in2 => \N__33762\,
            in3 => \N__36784\,
            lcout => \c0.n22149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i17_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40479\,
            in1 => \N__34233\,
            in2 => \_gnd_net_\,
            in3 => \N__35194\,
            lcout => encoder1_position_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i8_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40144\,
            in1 => \N__40565\,
            in2 => \_gnd_net_\,
            in3 => \N__34218\,
            lcout => encoder1_position_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1356_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45336\,
            in1 => \N__34206\,
            in2 => \N__34191\,
            in3 => \N__39780\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1358_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34170\,
            in1 => \N__34805\,
            in2 => \N__34161\,
            in3 => \N__42351\,
            lcout => \c0.n20455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1295_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40143\,
            in2 => \_gnd_net_\,
            in3 => \N__34109\,
            lcout => \c0.n20461\,
            ltout => \c0.n20461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1778_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40267\,
            in1 => \N__44773\,
            in2 => \N__34158\,
            in3 => \N__44370\,
            lcout => \c0.n22327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i25_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41325\,
            in1 => \N__37065\,
            in2 => \_gnd_net_\,
            in3 => \N__47657\,
            lcout => encoder0_position_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i27_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47658\,
            in1 => \N__36993\,
            in2 => \_gnd_net_\,
            in3 => \N__45587\,
            lcout => encoder0_position_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1339_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37188\,
            in1 => \N__34150\,
            in2 => \N__34614\,
            in3 => \N__34113\,
            lcout => \c0.n21364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i6_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42770\,
            in1 => \N__36723\,
            in2 => \_gnd_net_\,
            in3 => \N__47610\,
            lcout => encoder0_position_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78659\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1770_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41317\,
            in1 => \N__43415\,
            in2 => \N__36623\,
            in3 => \N__42535\,
            lcout => \c0.n22268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1761_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45519\,
            in1 => \N__46440\,
            in2 => \N__46361\,
            in3 => \N__45436\,
            lcout => \c0.n10497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20988_4_lut_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__40835\,
            in1 => \N__41054\,
            in2 => \N__34305\,
            in3 => \N__34287\,
            lcout => \c0.n24755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i24_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__37074\,
            in1 => \_gnd_net_\,
            in2 => \N__47652\,
            in3 => \N__42537\,
            lcout => encoder0_position_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78659\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1821_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41365\,
            in1 => \N__34262\,
            in2 => \N__44631\,
            in3 => \N__34448\,
            lcout => OPEN,
            ltout => \c0.n19_adj_4693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1819_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46179\,
            in1 => \N__37218\,
            in2 => \N__34245\,
            in3 => \N__34239\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4691_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1818_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41229\,
            in1 => \N__41943\,
            in2 => \N__34242\,
            in3 => \N__34455\,
            lcout => \c0.n20404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1820_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50584\,
            in1 => \N__41535\,
            in2 => \N__46448\,
            in3 => \N__45440\,
            lcout => \c0.n21_adj_4692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1312_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35033\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40079\,
            lcout => \c0.n22372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1420_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40080\,
            in1 => \N__35034\,
            in2 => \_gnd_net_\,
            in3 => \N__37201\,
            lcout => \c0.n20766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1791_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__41536\,
            in1 => \_gnd_net_\,
            in2 => \N__37170\,
            in3 => \N__41104\,
            lcout => \c0.n21457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1817_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__41179\,
            in1 => \N__37164\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n21489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1341_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44901\,
            in1 => \N__34377\,
            in2 => \N__34432\,
            in3 => \N__34389\,
            lcout => \c0.n21330\,
            ltout => \c0.n21330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1342_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__41107\,
            in1 => \_gnd_net_\,
            in2 => \N__34380\,
            in3 => \_gnd_net_\,
            lcout => \c0.n20511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1340_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__37577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45123\,
            lcout => \c0.n6_adj_4331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1990_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41108\,
            in1 => \N__34371\,
            in2 => \_gnd_net_\,
            in3 => \N__37169\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__0__5301_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__38021\,
            in1 => \N__34356\,
            in2 => \N__34323\,
            in3 => \N__37601\,
            lcout => \c0.data_out_frame_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78636\,
            ce => \N__45050\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34530\,
            in1 => \N__34518\,
            in2 => \_gnd_net_\,
            in3 => \N__43218\,
            lcout => \c0.n26_adj_4570\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45439\,
            in1 => \N__34781\,
            in2 => \N__45517\,
            in3 => \N__37258\,
            lcout => \c0.n10529\,
            ltout => \c0.n10529_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1293_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46789\,
            in2 => \N__34500\,
            in3 => \N__46247\,
            lcout => \c0.n21437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46790\,
            in1 => \N__34476\,
            in2 => \_gnd_net_\,
            in3 => \N__46752\,
            lcout => \c0.n21393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1285_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35285\,
            in2 => \_gnd_net_\,
            in3 => \N__45438\,
            lcout => \c0.n22489\,
            ltout => \c0.n22489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1289_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45507\,
            in1 => \N__41911\,
            in2 => \N__34497\,
            in3 => \N__34816\,
            lcout => \c0.n21416\,
            ltout => \c0.n21416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_2051_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101101001"
        )
    port map (
            in0 => \N__46522\,
            in1 => \N__41912\,
            in2 => \N__34494\,
            in3 => \_gnd_net_\,
            lcout => \c0.n22671\,
            ltout => \c0.n22671_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_2044_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35286\,
            in1 => \N__34491\,
            in2 => \N__34479\,
            in3 => \N__34817\,
            lcout => \c0.n20230\,
            ltout => \c0.n20230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__5__5288_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46884\,
            in1 => \N__46791\,
            in2 => \N__34470\,
            in3 => \N__45105\,
            lcout => \c0.data_out_frame_29_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78624\,
            ce => \N__45060\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__1__5468_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45994\,
            in1 => \N__48132\,
            in2 => \N__40227\,
            in3 => \N__34841\,
            lcout => data_out_frame_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i21_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34827\,
            in1 => \_gnd_net_\,
            in2 => \N__40575\,
            in3 => \N__40265\,
            lcout => encoder1_position_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1291_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35287\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34821\,
            lcout => \c0.n22722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1823_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34776\,
            in2 => \_gnd_net_\,
            in3 => \N__46348\,
            lcout => \c0.n22797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__0__5453_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45995\,
            in1 => \N__48133\,
            in2 => \N__36432\,
            in3 => \N__34691\,
            lcout => data_out_frame_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__4__5481_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48131\,
            in1 => \N__45996\,
            in2 => \N__43296\,
            in3 => \N__34673\,
            lcout => data_out_frame_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1337_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34654\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34602\,
            lcout => \c0.n22366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_8_i3_2_lut_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52695\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__71543\,
            lcout => \c0.n3_adj_4420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__2__5467_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__34544\,
            in1 => \N__46050\,
            in2 => \N__44871\,
            in3 => \N__48142\,
            lcout => data_out_frame_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__3__5426_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__46047\,
            in1 => \N__35078\,
            in2 => \N__48240\,
            in3 => \N__35133\,
            lcout => data_out_frame_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__2__5427_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__35060\,
            in1 => \N__48134\,
            in2 => \N__35039\,
            in3 => \N__46051\,
            lcout => data_out_frame_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i10_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40568\,
            in1 => \N__35046\,
            in2 => \_gnd_net_\,
            in3 => \N__35032\,
            lcout => encoder1_position_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__6__5479_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__46048\,
            in1 => \N__34991\,
            in2 => \N__48241\,
            in3 => \N__43408\,
            lcout => data_out_frame_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__7__5422_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__34928\,
            in1 => \N__46049\,
            in2 => \N__34975\,
            in3 => \N__48141\,
            lcout => data_out_frame_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1214_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__37833\,
            in1 => \N__41682\,
            in2 => \N__37827\,
            in3 => \N__38734\,
            lcout => \c0.n63_adj_4238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i28_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40563\,
            in1 => \N__34914\,
            in2 => \_gnd_net_\,
            in3 => \N__39962\,
            lcout => encoder1_position_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i27_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40562\,
            in2 => \N__34908\,
            in3 => \N__34888\,
            lcout => encoder1_position_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__3__5482_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48239\,
            in1 => \N__45993\,
            in2 => \N__46962\,
            in3 => \N__34856\,
            lcout => data_out_frame_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i29_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38674\,
            in1 => \N__35325\,
            in2 => \_gnd_net_\,
            in3 => \N__40564\,
            lcout => encoder1_position_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__6__5439_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48238\,
            in1 => \N__45992\,
            in2 => \N__35318\,
            in3 => \N__38808\,
            lcout => data_out_frame_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1209_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__38612\,
            in1 => \N__48632\,
            in2 => \N__44492\,
            in3 => \N__49242\,
            lcout => \c0.n16_adj_4233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__4__5417_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45983\,
            in1 => \N__48205\,
            in2 => \N__35298\,
            in3 => \N__35418\,
            lcout => data_out_frame_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__0__5461_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48204\,
            in1 => \N__45988\,
            in2 => \N__42882\,
            in3 => \N__35225\,
            lcout => data_out_frame_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__4__5465_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__45985\,
            in1 => \N__45348\,
            in2 => \N__48381\,
            in3 => \N__35507\,
            lcout => data_out_frame_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__1__5436_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48202\,
            in1 => \N__45986\,
            in2 => \N__35211\,
            in3 => \N__38306\,
            lcout => data_out_frame_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1211_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__39171\,
            in1 => \N__38568\,
            in2 => \N__41838\,
            in3 => \N__35172\,
            lcout => \c0.n63_adj_4235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__7__5430_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48203\,
            in1 => \N__45987\,
            in2 => \N__38553\,
            in3 => \N__35162\,
            lcout => data_out_frame_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__5__5416_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__45984\,
            in1 => \N__41190\,
            in2 => \N__48380\,
            in3 => \N__35147\,
            lcout => data_out_frame_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35417\,
            in1 => \N__43160\,
            in2 => \_gnd_net_\,
            in3 => \N__41718\,
            lcout => \c0.n11_adj_4669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__4__5457_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48207\,
            in1 => \N__45878\,
            in2 => \N__36500\,
            in3 => \N__42905\,
            lcout => data_out_frame_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i32_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__76384\,
            in1 => \N__50482\,
            in2 => \_gnd_net_\,
            in3 => \N__38761\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i6_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50481\,
            in1 => \N__42436\,
            in2 => \_gnd_net_\,
            in3 => \N__38847\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14067_3_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__35637\,
            in1 => \N__43623\,
            in2 => \_gnd_net_\,
            in3 => \N__35603\,
            lcout => \data_out_frame_29_7_N_2878_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__5__5456_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__48208\,
            in1 => \N__35399\,
            in2 => \N__42329\,
            in3 => \N__45879\,
            lcout => data_out_frame_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__5__5464_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__45876\,
            in1 => \N__48209\,
            in2 => \N__45672\,
            in3 => \N__35381\,
            lcout => data_out_frame_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__1__5444_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48206\,
            in1 => \N__45877\,
            in2 => \N__35367\,
            in3 => \N__38319\,
            lcout => data_out_frame_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1950_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39704\,
            in2 => \_gnd_net_\,
            in3 => \N__47814\,
            lcout => \c0.n8_adj_4555\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__4__5473_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__48364\,
            in1 => \N__35520\,
            in2 => \N__45997\,
            in3 => \N__36984\,
            lcout => data_out_frame_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1688_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35602\,
            in2 => \_gnd_net_\,
            in3 => \N__35651\,
            lcout => \c0.n7570\,
            ltout => \c0.n7570_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1671_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001111111111"
        )
    port map (
            in0 => \N__35471\,
            in1 => \N__43752\,
            in2 => \N__35523\,
            in3 => \N__43899\,
            lcout => \c0.n4_adj_4654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35519\,
            in1 => \N__43062\,
            in2 => \_gnd_net_\,
            in3 => \N__35511\,
            lcout => \c0.n5_adj_4217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1437_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__39240\,
            in1 => \N__43753\,
            in2 => \N__35430\,
            in3 => \N__43900\,
            lcout => \c0.n13055\,
            ltout => \c0.n13055_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1781_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__43967\,
            in1 => \N__44104\,
            in2 => \N__35493\,
            in3 => \N__43515\,
            lcout => n13058,
            ltout => \n13058_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__6__5463_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__48365\,
            in1 => \N__42267\,
            in2 => \N__35490\,
            in3 => \N__35486\,
            lcout => data_out_frame_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1531_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__44045\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43513\,
            lcout => \c0.n12992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1539_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35472\,
            in1 => \N__43611\,
            in2 => \N__47895\,
            in3 => \N__35953\,
            lcout => \c0.n5_adj_4477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__47235\,
            in1 => \N__47102\,
            in2 => \N__49638\,
            in3 => \N__47142\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1905_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43655\,
            in2 => \_gnd_net_\,
            in3 => \N__39333\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4727_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1907_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101110"
        )
    port map (
            in0 => \N__48510\,
            in1 => \N__35721\,
            in2 => \N__35694\,
            in3 => \N__35690\,
            lcout => \c0.n6_adj_4728\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1894_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101011"
        )
    port map (
            in0 => \N__39334\,
            in1 => \N__35689\,
            in2 => \N__48515\,
            in3 => \N__43865\,
            lcout => \c0.n24386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100110011"
        )
    port map (
            in0 => \N__35604\,
            in1 => \N__43809\,
            in2 => \N__43452\,
            in3 => \N__35652\,
            lcout => \c0.data_out_frame_29_7_N_1482_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1245_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39120\,
            in1 => \N__47366\,
            in2 => \N__45998\,
            in3 => \N__53807\,
            lcout => \c0.n2004\,
            ltout => \c0.n2004_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1572_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35653\,
            in1 => \N__35605\,
            in2 => \N__35574\,
            in3 => \N__43820\,
            lcout => \c0.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20970_4_lut_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__44327\,
            in1 => \N__36009\,
            in2 => \N__35571\,
            in3 => \N__39090\,
            lcout => \c0.n24736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1530_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__39755\,
            in1 => \_gnd_net_\,
            in2 => \N__35561\,
            in3 => \N__36159\,
            lcout => \c0.n28_adj_4565\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1658_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44325\,
            in1 => \N__35554\,
            in2 => \N__36166\,
            in3 => \N__39754\,
            lcout => \c0.n16919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1557_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__47894\,
            in1 => \N__43610\,
            in2 => \_gnd_net_\,
            in3 => \N__44326\,
            lcout => \c0.n6_adj_4583\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1475_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36081\,
            in1 => \N__36054\,
            in2 => \N__36042\,
            in3 => \N__36015\,
            lcout => \c0.n22145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1533_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36259\,
            in1 => \N__49036\,
            in2 => \N__35915\,
            in3 => \N__35849\,
            lcout => \c0.n20_adj_4265\,
            ltout => \c0.n20_adj_4265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1248_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47893\,
            in1 => \N__35999\,
            in2 => \N__35985\,
            in3 => \N__35922\,
            lcout => \c0.n22148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1247_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43609\,
            in2 => \_gnd_net_\,
            in3 => \N__35943\,
            lcout => \c0.n6_adj_4264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_1963_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35916\,
            in1 => \N__36266\,
            in2 => \N__35871\,
            in3 => \N__35853\,
            lcout => \c0.n7_adj_4741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_2003_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__49829\,
            in1 => \N__39250\,
            in2 => \N__53916\,
            in3 => \N__43836\,
            lcout => \c0.n9683\,
            ltout => \c0.n9683_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__35799\,
            in1 => \N__48475\,
            in2 => \N__35790\,
            in3 => \N__44276\,
            lcout => \c0.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1981_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49073\,
            lcout => \c0.n21643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_2008_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36267\,
            in2 => \_gnd_net_\,
            in3 => \N__47818\,
            lcout => \c0.n21653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1971_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39744\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47815\,
            lcout => \c0.n21639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1976_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__47816\,
            in1 => \_gnd_net_\,
            in2 => \N__49139\,
            in3 => \_gnd_net_\,
            lcout => \c0.n21641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i29_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36205\,
            in2 => \_gnd_net_\,
            in3 => \N__48985\,
            lcout => \c0.FRAME_MATCHER_state_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78716\,
            ce => 'H',
            sr => \N__36183\
        );

    \c0.FRAME_MATCHER_state_i24_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48987\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36155\,
            lcout => \c0.FRAME_MATCHER_state_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78728\,
            ce => 'H',
            sr => \N__36126\
        );

    \c0.FRAME_MATCHER_state_i21_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49069\,
            in2 => \_gnd_net_\,
            in3 => \N__48989\,
            lcout => \c0.FRAME_MATCHER_state_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78741\,
            ce => 'H',
            sr => \N__36111\
        );

    \quad_counter0.count_i0_i2_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47728\,
            in1 => \N__36300\,
            in2 => \_gnd_net_\,
            in3 => \N__39840\,
            lcout => encoder0_position_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i3_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44755\,
            in1 => \N__36291\,
            in2 => \_gnd_net_\,
            in3 => \N__47730\,
            lcout => encoder0_position_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i7_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36689\,
            in1 => \N__36645\,
            in2 => \_gnd_net_\,
            in3 => \N__47731\,
            lcout => encoder0_position_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i30_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39612\,
            in1 => \N__36825\,
            in2 => \_gnd_net_\,
            in3 => \N__47729\,
            lcout => encoder0_position_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i0_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47727\,
            in1 => \N__36372\,
            in2 => \_gnd_net_\,
            in3 => \N__36414\,
            lcout => encoder0_position_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_1_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37384\,
            in2 => \N__37447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \quad_counter0.n19763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_2_lut_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36413\,
            in2 => \N__36387\,
            in3 => \N__36366\,
            lcout => n2357,
            ltout => OPEN,
            carryin => \quad_counter0.n19763\,
            carryout => \quad_counter0.n19764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_3_lut_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36356\,
            in2 => \N__37448\,
            in3 => \N__36303\,
            lcout => n2356,
            ltout => OPEN,
            carryin => \quad_counter0.n19764\,
            carryout => \quad_counter0.n19765\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_4_lut_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39836\,
            in2 => \N__37444\,
            in3 => \N__36294\,
            lcout => n2355,
            ltout => OPEN,
            carryin => \quad_counter0.n19765\,
            carryout => \quad_counter0.n19766\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_5_lut_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44774\,
            in2 => \N__37449\,
            in3 => \N__36285\,
            lcout => n2354,
            ltout => OPEN,
            carryin => \quad_counter0.n19766\,
            carryout => \quad_counter0.n19767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_6_lut_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45263\,
            in2 => \N__37445\,
            in3 => \N__36270\,
            lcout => n2353,
            ltout => OPEN,
            carryin => \quad_counter0.n19767\,
            carryout => \quad_counter0.n19768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_7_lut_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45380\,
            in2 => \N__37450\,
            in3 => \N__36726\,
            lcout => n2352,
            ltout => OPEN,
            carryin => \quad_counter0.n19768\,
            carryout => \quad_counter0.n19769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_8_lut_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42771\,
            in2 => \N__37446\,
            in3 => \N__36714\,
            lcout => n2351,
            ltout => OPEN,
            carryin => \quad_counter0.n19769\,
            carryout => \quad_counter0.n19770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_9_lut_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36693\,
            in2 => \N__37484\,
            in3 => \N__36636\,
            lcout => n2350,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \quad_counter0.n19771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_10_lut_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37454\,
            in2 => \N__42881\,
            in3 => \N__36633\,
            lcout => n2349,
            ltout => OPEN,
            carryin => \quad_counter0.n19771\,
            carryout => \quad_counter0.n19772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_11_lut_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42656\,
            in2 => \N__37485\,
            in3 => \N__36630\,
            lcout => n2348,
            ltout => OPEN,
            carryin => \quad_counter0.n19772\,
            carryout => \quad_counter0.n19773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_12_lut_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37458\,
            in2 => \N__36627\,
            in3 => \N__36567\,
            lcout => n2347,
            ltout => OPEN,
            carryin => \quad_counter0.n19773\,
            carryout => \quad_counter0.n19774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_13_lut_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36554\,
            in2 => \N__37486\,
            in3 => \N__36507\,
            lcout => n2346,
            ltout => OPEN,
            carryin => \quad_counter0.n19774\,
            carryout => \quad_counter0.n19775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_14_lut_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37462\,
            in2 => \N__36504\,
            in3 => \N__36435\,
            lcout => n2345,
            ltout => OPEN,
            carryin => \quad_counter0.n19775\,
            carryout => \quad_counter0.n19776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_15_lut_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42328\,
            in2 => \N__37487\,
            in3 => \N__36813\,
            lcout => n2344,
            ltout => OPEN,
            carryin => \quad_counter0.n19776\,
            carryout => \quad_counter0.n19777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_16_lut_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37466\,
            in2 => \N__47501\,
            in3 => \N__36810\,
            lcout => n2343,
            ltout => OPEN,
            carryin => \quad_counter0.n19777\,
            carryout => \quad_counter0.n19778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_17_lut_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39554\,
            in2 => \N__37488\,
            in3 => \N__36807\,
            lcout => n2342,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \quad_counter0.n19779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_18_lut_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37470\,
            in2 => \N__36804\,
            in3 => \N__36744\,
            lcout => n2341,
            ltout => OPEN,
            carryin => \quad_counter0.n19779\,
            carryout => \quad_counter0.n19780\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_19_lut_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40213\,
            in2 => \N__37489\,
            in3 => \N__36741\,
            lcout => n2340,
            ltout => OPEN,
            carryin => \quad_counter0.n19780\,
            carryout => \quad_counter0.n19781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_20_lut_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37474\,
            in2 => \N__44863\,
            in3 => \N__36738\,
            lcout => n2339,
            ltout => OPEN,
            carryin => \quad_counter0.n19781\,
            carryout => \quad_counter0.n19782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_21_lut_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42401\,
            in2 => \N__37490\,
            in3 => \N__36735\,
            lcout => n2338,
            ltout => OPEN,
            carryin => \quad_counter0.n19782\,
            carryout => \quad_counter0.n19783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_22_lut_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37478\,
            in2 => \N__45344\,
            in3 => \N__36732\,
            lcout => n2337,
            ltout => OPEN,
            carryin => \quad_counter0.n19783\,
            carryout => \quad_counter0.n19784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_23_lut_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37479\,
            in2 => \N__45656\,
            in3 => \N__36729\,
            lcout => n2336,
            ltout => OPEN,
            carryin => \quad_counter0.n19784\,
            carryout => \quad_counter0.n19785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_24_lut_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42257\,
            in2 => \N__37491\,
            in3 => \N__37080\,
            lcout => n2335,
            ltout => OPEN,
            carryin => \quad_counter0.n19785\,
            carryout => \quad_counter0.n19786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_25_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37337\,
            in2 => \N__42716\,
            in3 => \N__37077\,
            lcout => n2334,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \quad_counter0.n19787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_26_lut_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42536\,
            in2 => \N__37380\,
            in3 => \N__37068\,
            lcout => n2333,
            ltout => OPEN,
            carryin => \quad_counter0.n19787\,
            carryout => \quad_counter0.n19788\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_27_lut_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37341\,
            in2 => \N__41327\,
            in3 => \N__37059\,
            lcout => n2332,
            ltout => OPEN,
            carryin => \quad_counter0.n19788\,
            carryout => \quad_counter0.n19789\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_28_lut_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37052\,
            in2 => \N__37381\,
            in3 => \N__36996\,
            lcout => n2331,
            ltout => OPEN,
            carryin => \quad_counter0.n19789\,
            carryout => \quad_counter0.n19790\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_29_lut_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37345\,
            in2 => \N__45614\,
            in3 => \N__36987\,
            lcout => n2330,
            ltout => OPEN,
            carryin => \quad_counter0.n19790\,
            carryout => \quad_counter0.n19791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_30_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36977\,
            in2 => \N__37382\,
            in3 => \N__36900\,
            lcout => n2329,
            ltout => OPEN,
            carryin => \quad_counter0.n19791\,
            carryout => \quad_counter0.n19792\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_31_lut_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37349\,
            in2 => \N__36893\,
            in3 => \N__36828\,
            lcout => n2328,
            ltout => OPEN,
            carryin => \quad_counter0.n19792\,
            carryout => \quad_counter0.n19793\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_32_lut_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39624\,
            in2 => \N__37383\,
            in3 => \N__36816\,
            lcout => n2327,
            ltout => OPEN,
            carryin => \quad_counter0.n19793\,
            carryout => \quad_counter0.n19794\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_647_33_lut_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44684\,
            in1 => \N__37483\,
            in2 => \_gnd_net_\,
            in3 => \N__37293\,
            lcout => OPEN,
            ltout => \n2326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i31_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44685\,
            in2 => \N__37290\,
            in3 => \N__47696\,
            lcout => encoder0_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1364_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44683\,
            in2 => \_gnd_net_\,
            in3 => \N__45174\,
            lcout => \c0.n10427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1822_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__37637\,
            in1 => \N__37283\,
            in2 => \N__37266\,
            in3 => \N__37227\,
            lcout => \c0.n20_adj_4694\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1782_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37208\,
            in1 => \N__50528\,
            in2 => \N__40022\,
            in3 => \N__41102\,
            lcout => \c0.n21355\,
            ltout => \c0.n21355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1790_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41103\,
            in1 => \N__37168\,
            in2 => \N__37146\,
            in3 => \N__41537\,
            lcout => \c0.n21327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_1799_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37143\,
            in2 => \_gnd_net_\,
            in3 => \N__37092\,
            lcout => \c0.n15_adj_4686\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1219_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__38493\,
            in1 => \N__41820\,
            in2 => \N__44485\,
            in3 => \N__48606\,
            lcout => \c0.n13046\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i18_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41821\,
            in1 => \_gnd_net_\,
            in2 => \N__49314\,
            in3 => \N__50438\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1784_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37638\,
            in1 => \N__46610\,
            in2 => \N__46873\,
            in3 => \N__37597\,
            lcout => \c0.n24028\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1792_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41106\,
            in1 => \N__46854\,
            in2 => \_gnd_net_\,
            in3 => \N__50526\,
            lcout => \c0.n13268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i22_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47711\,
            in1 => \N__37626\,
            in2 => \_gnd_net_\,
            in3 => \N__42247\,
            lcout => encoder0_position_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1301_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44433\,
            in1 => \N__45261\,
            in2 => \N__37617\,
            in3 => \N__37556\,
            lcout => \c0.n21360\,
            ltout => \c0.n21360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1296_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41105\,
            in2 => \N__37608\,
            in3 => \_gnd_net_\,
            lcout => \c0.n10504\,
            ltout => \c0.n10504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1299_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37581\,
            in1 => \N__44699\,
            in2 => \N__37560\,
            in3 => \N__37557\,
            lcout => \c0.n12_adj_4312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1880_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37545\,
            in1 => \N__41589\,
            in2 => \N__41189\,
            in3 => \N__46671\,
            lcout => OPEN,
            ltout => \c0.n25_adj_4695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__1__5292_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__37521\,
            in1 => \N__37671\,
            in2 => \N__37509\,
            in3 => \N__37752\,
            lcout => \c0.data_out_frame_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78638\,
            ce => \N__45059\,
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1884_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37785\,
            in1 => \N__37778\,
            in2 => \N__37761\,
            in3 => \N__41448\,
            lcout => \c0.n26_adj_4697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__1__5300_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37743\,
            in1 => \N__37725\,
            in2 => \_gnd_net_\,
            in3 => \N__37710\,
            lcout => \c0.data_out_frame_28_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78638\,
            ce => \N__45059\,
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1834_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38006\,
            in1 => \N__41067\,
            in2 => \N__37683\,
            in3 => \N__46155\,
            lcout => \c0.n27_adj_4696\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i8_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48628\,
            in1 => \N__50429\,
            in2 => \_gnd_net_\,
            in3 => \N__38988\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78626\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i5_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37652\,
            in1 => \N__50428\,
            in2 => \_gnd_net_\,
            in3 => \N__37826\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78626\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i1_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__42063\,
            in1 => \_gnd_net_\,
            in2 => \N__50465\,
            in3 => \N__37665\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78626\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1215_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__43363\,
            in1 => \N__37664\,
            in2 => \N__37653\,
            in3 => \N__38987\,
            lcout => \c0.n10_adj_4239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1221_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__37860\,
            in1 => \N__44525\,
            in2 => \N__42066\,
            in3 => \N__37878\,
            lcout => OPEN,
            ltout => \c0.n15_adj_4242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1222_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__41698\,
            in1 => \N__38736\,
            in2 => \N__37641\,
            in3 => \N__37791\,
            lcout => \c0.n12898\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1806_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__38258\,
            in1 => \N__38175\,
            in2 => \_gnd_net_\,
            in3 => \N__38082\,
            lcout => \c0.n21464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i24_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37962\,
            in1 => \N__40573\,
            in2 => \_gnd_net_\,
            in3 => \N__37926\,
            lcout => encoder1_position_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i21_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37865\,
            in1 => \N__50426\,
            in2 => \_gnd_net_\,
            in3 => \N__42092\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i174_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__75909\,
            in1 => \N__79786\,
            in2 => \_gnd_net_\,
            in3 => \N__67648\,
            lcout => data_in_frame_21_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1384_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47014\,
            in2 => \_gnd_net_\,
            in3 => \N__42341\,
            lcout => \c0.n10_adj_4367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1216_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__42091\,
            in1 => \N__39009\,
            in2 => \_gnd_net_\,
            in3 => \N__37884\,
            lcout => \c0.n13049\,
            ltout => \c0.n13049_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1212_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__42438\,
            in1 => \N__37861\,
            in2 => \N__37839\,
            in3 => \N__38630\,
            lcout => OPEN,
            ltout => \c0.n18_adj_4236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1213_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__44526\,
            in1 => \N__49424\,
            in2 => \N__37836\,
            in3 => \N__38585\,
            lcout => \c0.n20_adj_4237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1220_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__42437\,
            in1 => \N__37822\,
            in2 => \_gnd_net_\,
            in3 => \N__49423\,
            lcout => \c0.n14_adj_4241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1210_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__46919\,
            in1 => \N__49310\,
            in2 => \N__38586\,
            in3 => \N__48679\,
            lcout => \c0.n17_adj_4234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i23_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38562\,
            in1 => \N__40558\,
            in2 => \_gnd_net_\,
            in3 => \N__38535\,
            lcout => encoder1_position_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78627\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i13_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47732\,
            in1 => \N__38508\,
            in2 => \_gnd_net_\,
            in3 => \N__42297\,
            lcout => encoder0_position_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78627\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1217_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39170\,
            in2 => \_gnd_net_\,
            in3 => \N__46918\,
            lcout => \c0.n10_adj_4240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__38393\,
            in1 => \N__38482\,
            in2 => \_gnd_net_\,
            in3 => \N__38415\,
            lcout => \c0.tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78627\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i26_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40569\,
            in1 => \N__38379\,
            in2 => \_gnd_net_\,
            in3 => \N__38343\,
            lcout => encoder1_position_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__38318\,
            in1 => \N__40821\,
            in2 => \N__38307\,
            in3 => \N__43221\,
            lcout => OPEN,
            ltout => \c0.n25116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n25116_bdd_4_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__40822\,
            in1 => \N__38693\,
            in2 => \N__38292\,
            in3 => \N__38289\,
            lcout => \c0.n25119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_1168_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__47227\,
            in1 => \N__46656\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n12981,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i11_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50472\,
            in1 => \N__38735\,
            in2 => \_gnd_net_\,
            in3 => \N__49264\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__1__5460_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48200\,
            in1 => \N__46011\,
            in2 => \N__38697\,
            in3 => \N__42663\,
            lcout => data_out_frame_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__5__5440_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__46010\,
            in1 => \N__48201\,
            in2 => \N__38649\,
            in3 => \N__38675\,
            lcout => data_out_frame_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1690_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__38846\,
            in1 => \N__38631\,
            in2 => \N__42122\,
            in3 => \N__38616\,
            lcout => OPEN,
            ltout => \c0.n20_adj_4308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_1290_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38595\,
            in2 => \N__38598\,
            in3 => \N__38886\,
            lcout => n63,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1691_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__44558\,
            in1 => \N__42466\,
            in2 => \N__38762\,
            in3 => \N__38879\,
            lcout => \c0.n19_adj_4307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1206_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__42200\,
            in1 => \N__44557\,
            in2 => \N__42470\,
            in3 => \N__49260\,
            lcout => OPEN,
            ltout => \c0.n16_adj_4231_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1208_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__38754\,
            in1 => \N__42114\,
            in2 => \N__38589\,
            in3 => \N__38829\,
            lcout => \c0.n12986\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20978_4_lut_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43318\,
            in1 => \N__42201\,
            in2 => \N__49268\,
            in3 => \N__43346\,
            lcout => \c0.n24745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1207_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__43345\,
            in1 => \N__43317\,
            in2 => \N__38880\,
            in3 => \N__38845\,
            lcout => \c0.n17_adj_4232\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i192_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__80988\,
            in1 => \N__63965\,
            in2 => \N__76382\,
            in3 => \N__80429\,
            lcout => \c0.data_in_frame_23_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i30_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38823\,
            in1 => \N__40574\,
            in2 => \_gnd_net_\,
            in3 => \N__38787\,
            lcout => encoder1_position_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1742_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__44141\,
            in1 => \N__39109\,
            in2 => \_gnd_net_\,
            in3 => \N__44103\,
            lcout => \c0.n13001\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i88_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__61719\,
            in1 => \N__73707\,
            in2 => \N__76383\,
            in3 => \N__69236\,
            lcout => \c0.data_in_frame_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i24_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38763\,
            in1 => \N__50462\,
            in2 => \_gnd_net_\,
            in3 => \N__39007\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i213_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__79442\,
            in1 => \N__69237\,
            in2 => \N__77332\,
            in3 => \N__71887\,
            lcout => \c0.data_in_frame_26_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i212_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__69235\,
            in1 => \N__68349\,
            in2 => \N__76916\,
            in3 => \N__79443\,
            lcout => \c0.data_in_frame_26_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i30_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50460\,
            in1 => \N__79648\,
            in2 => \_gnd_net_\,
            in3 => \N__39168\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i22_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39169\,
            in1 => \N__50461\,
            in2 => \_gnd_net_\,
            in3 => \N__42462\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__47429\,
            in1 => \N__76883\,
            in2 => \N__50908\,
            in3 => \N__50726\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i237_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__56481\,
            in1 => \N__52013\,
            in2 => \N__71938\,
            in3 => \N__75397\,
            lcout => \c0.data_in_frame_29_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_2046_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__43493\,
            in1 => \N__39370\,
            in2 => \N__44011\,
            in3 => \N__39421\,
            lcout => \c0.n13063\,
            ltout => \c0.n13063_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_2047_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__39422\,
            in1 => \N__39371\,
            in2 => \N__39123\,
            in3 => \N__39020\,
            lcout => \c0.n6_adj_4263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1979_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__39108\,
            in1 => \N__38967\,
            in2 => \N__44331\,
            in3 => \N__39336\,
            lcout => \c0.n8_adj_4553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1265_2_lut_3_lut_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__44131\,
            in1 => \N__39097\,
            in2 => \_gnd_net_\,
            in3 => \N__43492\,
            lcout => \c0.n3325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i16_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50463\,
            in1 => \N__39008\,
            in2 => \_gnd_net_\,
            in3 => \N__38981\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1961_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__43605\,
            in1 => \N__38966\,
            in2 => \_gnd_net_\,
            in3 => \N__38933\,
            lcout => \c0.n21659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1779_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__44002\,
            in1 => \N__44058\,
            in2 => \N__48519\,
            in3 => \N__44108\,
            lcout => \c0.n24422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_2041_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__39465\,
            in1 => \N__39423\,
            in2 => \N__39399\,
            in3 => \N__39375\,
            lcout => OPEN,
            ltout => \c0.n24596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1287_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000100"
        )
    port map (
            in0 => \N__39348\,
            in1 => \N__43514\,
            in2 => \N__39339\,
            in3 => \N__39335\,
            lcout => \c0.n4_adj_4306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4626_2_lut_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48270\,
            in2 => \_gnd_net_\,
            in3 => \N__45889\,
            lcout => \c0.n8162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50048\,
            in2 => \_gnd_net_\,
            in3 => \N__39314\,
            lcout => OPEN,
            ltout => \c0.rx.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i21269_4_lut_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__50161\,
            in1 => \N__49962\,
            in2 => \N__39282\,
            in3 => \N__50867\,
            lcout => n14439,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1840_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__43709\,
            in1 => \N__39258\,
            in2 => \N__43842\,
            in3 => \N__43445\,
            lcout => OPEN,
            ltout => \c0.n24302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1896_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__43667\,
            in1 => \N__39219\,
            in2 => \N__39210\,
            in3 => \N__43531\,
            lcout => \c0.n4_adj_4721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1939_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39207\,
            in2 => \_gnd_net_\,
            in3 => \N__47827\,
            lcout => \c0.n8_adj_4556\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i18_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39745\,
            in2 => \_gnd_net_\,
            in3 => \N__48986\,
            lcout => \c0.FRAME_MATCHER_state_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78729\,
            ce => 'H',
            sr => \N__39717\
        );

    \c0.FRAME_MATCHER_state_i12_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48988\,
            in2 => \_gnd_net_\,
            in3 => \N__39694\,
            lcout => \c0.FRAME_MATCHER_state_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78742\,
            ce => 'H',
            sr => \N__39672\
        );

    \c0.FRAME_MATCHER_state_i19_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49129\,
            in2 => \_gnd_net_\,
            in3 => \N__48990\,
            lcout => \c0.FRAME_MATCHER_state_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78755\,
            ce => 'H',
            sr => \N__39657\
        );

    \c0.i1_2_lut_3_lut_adj_1999_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39529\,
            in1 => \N__39595\,
            in2 => \_gnd_net_\,
            in3 => \N__39779\,
            lcout => \c0.n22785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i15_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39567\,
            in1 => \N__47724\,
            in2 => \_gnd_net_\,
            in3 => \N__39542\,
            lcout => encoder0_position_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i5_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45381\,
            in1 => \N__39504\,
            in2 => \_gnd_net_\,
            in3 => \N__47725\,
            lcout => encoder0_position_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14227_2_lut_3_lut_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__74279\,
            in1 => \N__74643\,
            in2 => \_gnd_net_\,
            in3 => \N__74441\,
            lcout => \c0.n17830\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1915_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__49155\,
            in1 => \N__51627\,
            in2 => \N__57159\,
            in3 => \N__61335\,
            lcout => OPEN,
            ltout => \c0.n30_adj_4730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1931_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48570\,
            in1 => \N__44439\,
            in2 => \N__39498\,
            in3 => \N__51252\,
            lcout => \c0.n17539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40021\,
            in1 => \N__44345\,
            in2 => \N__39989\,
            in3 => \N__42655\,
            lcout => \c0.n31_adj_4325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_1_i3_2_lut_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__74447\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__71538\,
            lcout => \c0.n3_adj_4434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1313_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45382\,
            in1 => \N__45626\,
            in2 => \N__42788\,
            in3 => \N__43285\,
            lcout => \c0.n22775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i9_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__39891\,
            in1 => \_gnd_net_\,
            in2 => \N__47733\,
            in3 => \N__42657\,
            lcout => encoder0_position_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i21_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45655\,
            in1 => \N__39885\,
            in2 => \_gnd_net_\,
            in3 => \N__47716\,
            lcout => encoder0_position_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1294_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39879\,
            in1 => \N__39848\,
            in2 => \_gnd_net_\,
            in3 => \N__39798\,
            lcout => \c0.n13422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1756_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44686\,
            in1 => \N__45173\,
            in2 => \_gnd_net_\,
            in3 => \N__40204\,
            lcout => \c0.n13630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i17_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40205\,
            in1 => \N__47715\,
            in2 => \_gnd_net_\,
            in3 => \N__39762\,
            lcout => encoder0_position_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101011010000"
        )
    port map (
            in0 => \N__41055\,
            in1 => \N__40854\,
            in2 => \N__40836\,
            in3 => \N__40611\,
            lcout => \c0.n25062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1320_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43275\,
            in2 => \_gnd_net_\,
            in3 => \N__42262\,
            lcout => \c0.n22635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1255_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45116\,
            in2 => \_gnd_net_\,
            in3 => \N__42143\,
            lcout => \c0.n6_adj_4276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1317_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42380\,
            in2 => \_gnd_net_\,
            in3 => \N__40206\,
            lcout => \c0.n13558\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i31_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__40314\,
            in1 => \N__40590\,
            in2 => \N__40566\,
            in3 => \_gnd_net_\,
            lcout => encoder1_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i19_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47611\,
            in1 => \N__40284\,
            in2 => \_gnd_net_\,
            in3 => \N__42381\,
            lcout => encoder0_position_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i90_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76613\,
            in1 => \N__73651\,
            in2 => \N__65286\,
            in3 => \N__75195\,
            lcout => \c0.data_in_frame_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1777_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40274\,
            in1 => \N__42389\,
            in2 => \_gnd_net_\,
            in3 => \N__40214\,
            lcout => \c0.n22580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1256_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40178\,
            in1 => \N__40128\,
            in2 => \N__40094\,
            in3 => \N__40038\,
            lcout => \c0.n10467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i28_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50437\,
            in1 => \N__76997\,
            in2 => \_gnd_net_\,
            in3 => \N__48666\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1284_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46349\,
            in2 => \_gnd_net_\,
            in3 => \N__46444\,
            lcout => \c0.n21441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__1__5476_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__48086\,
            in1 => \N__41276\,
            in2 => \N__41334\,
            in3 => \N__46094\,
            lcout => data_out_frame_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__4__5449_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__46092\,
            in1 => \N__48087\,
            in2 => \N__45267\,
            in3 => \N__42923\,
            lcout => data_out_frame_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__2__5291_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48085\,
            in1 => \N__46093\,
            in2 => \N__41261\,
            in3 => \N__41865\,
            lcout => data_out_frame_29_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1300_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41907\,
            in1 => \N__44864\,
            in2 => \N__45285\,
            in3 => \N__41241\,
            lcout => \c0.n24113\,
            ltout => \c0.n24113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_2019_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41181\,
            in1 => \N__44899\,
            in2 => \N__41235\,
            in3 => \N__50527\,
            lcout => \c0.n21349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1436_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41231\,
            in2 => \_gnd_net_\,
            in3 => \N__46484\,
            lcout => \c0.n21358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_2021_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41180\,
            in1 => \N__44900\,
            in2 => \N__41115\,
            in3 => \N__41066\,
            lcout => \c0.n21311\,
            ltout => \c0.n21311_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_2050_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__46270\,
            in1 => \_gnd_net_\,
            in2 => \N__41670\,
            in3 => \N__46815\,
            lcout => OPEN,
            ltout => \c0.n21273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__6__5295_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41667\,
            in1 => \N__41646\,
            in2 => \N__41625\,
            in3 => \N__46461\,
            lcout => \c0.data_out_frame_28_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78663\,
            ce => \N__45041\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43223\,
            in1 => \N__41622\,
            in2 => \_gnd_net_\,
            in3 => \N__41610\,
            lcout => \c0.n26_adj_4702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1797_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41588\,
            in1 => \N__41454\,
            in2 => \N__46264\,
            in3 => \N__41922\,
            lcout => OPEN,
            ltout => \c0.n18_adj_4684_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1798_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41571\,
            in1 => \N__45098\,
            in2 => \N__41541\,
            in3 => \N__41538\,
            lcout => OPEN,
            ltout => \c0.n20_adj_4685_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__7__5294_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41945\,
            in1 => \N__41517\,
            in2 => \N__41505\,
            in3 => \N__41502\,
            lcout => \c0.data_out_frame_28_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78651\,
            ce => \N__45055\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1743_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46139\,
            in1 => \N__46498\,
            in2 => \_gnd_net_\,
            in3 => \N__46151\,
            lcout => \c0.n22461\,
            ltout => \c0.n22461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1440_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41447\,
            in1 => \N__46716\,
            in2 => \N__41436\,
            in3 => \N__41921\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4478_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1470_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41433\,
            in1 => \N__41944\,
            in2 => \N__41925\,
            in3 => \N__46539\,
            lcout => \data_out_frame_29__2__N_1748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1438_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46533\,
            in2 => \_gnd_net_\,
            in3 => \N__46460\,
            lcout => \c0.n22193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1888_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41913\,
            in1 => \N__46632\,
            in2 => \N__41877\,
            in3 => \N__41861\,
            lcout => \c0.n19_adj_4720\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i96_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__73520\,
            in1 => \N__76625\,
            in2 => \N__76398\,
            in3 => \N__55611\,
            lcout => \c0.data_in_frame_11_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i10_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50424\,
            in1 => \N__41837\,
            in2 => \_gnd_net_\,
            in3 => \N__43367\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i4_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41700\,
            in1 => \N__50423\,
            in2 => \_gnd_net_\,
            in3 => \N__42123\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__3__5290_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__46078\,
            in1 => \N__48188\,
            in2 => \N__41801\,
            in3 => \N__46670\,
            lcout => data_out_frame_29_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__4__5425_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48187\,
            in1 => \N__46079\,
            in2 => \N__41781\,
            in3 => \N__41714\,
            lcout => data_out_frame_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41699\,
            in2 => \_gnd_net_\,
            in3 => \N__42064\,
            lcout => \c0.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i29_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__71916\,
            in1 => \N__50427\,
            in2 => \_gnd_net_\,
            in3 => \N__42093\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i93_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76624\,
            in1 => \N__73522\,
            in2 => \N__70774\,
            in3 => \N__71917\,
            lcout => \c0.data_in_frame_11_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i23_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47721\,
            in1 => \N__42078\,
            in2 => \_gnd_net_\,
            in3 => \N__42701\,
            lcout => encoder0_position_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i224_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__79464\,
            in1 => \N__76355\,
            in2 => \N__56560\,
            in3 => \N__76653\,
            lcout => \c0.data_in_frame_27_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i9_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50425\,
            in1 => \N__42065\,
            in2 => \_gnd_net_\,
            in3 => \N__42194\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i217_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__79463\,
            in1 => \N__80616\,
            in2 => \N__75678\,
            in3 => \N__76652\,
            lcout => \c0.data_in_frame_27_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i8_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47722\,
            in1 => \N__42042\,
            in2 => \_gnd_net_\,
            in3 => \N__42855\,
            lcout => encoder0_position_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_4_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__42026\,
            in1 => \N__50034\,
            in2 => \N__50183\,
            in3 => \N__49940\,
            lcout => \c0.rx.n12909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i236_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__77045\,
            in1 => \N__56480\,
            in2 => \N__47408\,
            in3 => \N__75326\,
            lcout => \c0.data_in_frame_29_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1363_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43396\,
            in2 => \_gnd_net_\,
            in3 => \N__42559\,
            lcout => OPEN,
            ltout => \c0.n22199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1383_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42390\,
            in1 => \N__42845\,
            in2 => \N__42354\,
            in3 => \N__42207\,
            lcout => \c0.n22834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1360_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42288\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47456\,
            lcout => \c0.n13665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1752_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__47051\,
            in1 => \N__42688\,
            in2 => \_gnd_net_\,
            in3 => \N__42261\,
            lcout => \c0.n6_adj_4366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i17_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__42193\,
            in1 => \N__50404\,
            in2 => \_gnd_net_\,
            in3 => \N__49425\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14131_2_lut_3_lut_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__50403\,
            in1 => \N__50208\,
            in2 => \_gnd_net_\,
            in3 => \N__53802\,
            lcout => \c0.n17734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i7_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42597\,
            in1 => \N__71133\,
            in2 => \_gnd_net_\,
            in3 => \N__47351\,
            lcout => control_mode_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1336_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46949\,
            in2 => \_gnd_net_\,
            in3 => \N__45340\,
            lcout => OPEN,
            ltout => \c0.n22256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1270_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42170\,
            in1 => \N__42726\,
            in2 => \N__42150\,
            in3 => \N__47276\,
            lcout => \c0.n22772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i12_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50483\,
            in1 => \N__42121\,
            in2 => \_gnd_net_\,
            in3 => \N__46920\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i4_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43274\,
            in1 => \N__60573\,
            in2 => \_gnd_net_\,
            in3 => \N__47350\,
            lcout => control_mode_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21015_3_lut_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43186\,
            in1 => \N__42924\,
            in2 => \_gnd_net_\,
            in3 => \N__42909\,
            lcout => \c0.n24782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i0_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45158\,
            in1 => \N__61068\,
            in2 => \_gnd_net_\,
            in3 => \N__47349\,
            lcout => control_mode_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1321_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42703\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42856\,
            lcout => \c0.n22423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1268_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47053\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42787\,
            lcout => \c0.n6_adj_4293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1382_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__42702\,
            in1 => \N__47052\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n22385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1304_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42659\,
            in1 => \N__42601\,
            in2 => \N__42570\,
            in3 => \N__42560\,
            lcout => \c0.n20325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i14_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__42427\,
            in1 => \N__50464\,
            in2 => \_gnd_net_\,
            in3 => \N__42471\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i225_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__80605\,
            in1 => \N__80094\,
            in2 => \N__51800\,
            in3 => \N__79420\,
            lcout => \c0.data_in_frame_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13969_2_lut_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49730\,
            in3 => \N__49648\,
            lcout => n17571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_107_i4_2_lut_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__49649\,
            in1 => \N__49723\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n4_adj_4762,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i6_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43395\,
            in1 => \N__58056\,
            in2 => \_gnd_net_\,
            in3 => \N__47348\,
            lcout => control_mode_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i195_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__67532\,
            in1 => \N__79084\,
            in2 => \N__72996\,
            in3 => \N__79366\,
            lcout => \c0.data_in_frame_24_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14114_2_lut_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53894\,
            in2 => \_gnd_net_\,
            in3 => \N__49828\,
            lcout => \c0.n937\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i2_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50458\,
            in1 => \N__43347\,
            in2 => \_gnd_net_\,
            in3 => \N__43371\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i27_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__79083\,
            in1 => \N__50459\,
            in2 => \N__43328\,
            in3 => \_gnd_net_\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19184_3_lut_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__44046\,
            in1 => \N__44158\,
            in2 => \_gnd_net_\,
            in3 => \N__44269\,
            lcout => \c0.n17856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i155_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__76675\,
            in1 => \N__80428\,
            in2 => \N__79141\,
            in3 => \N__63328\,
            lcout => \c0.data_in_frame_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i173_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__67640\,
            in1 => \_gnd_net_\,
            in2 => \N__71966\,
            in3 => \N__66746\,
            lcout => data_in_frame_21_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53448\,
            in2 => \_gnd_net_\,
            in3 => \N__52769\,
            lcout => \c0.n39_adj_4295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_7_i3_2_lut_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52632\,
            in2 => \_gnd_net_\,
            in3 => \N__71428\,
            lcout => \c0.n3_adj_4422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1280_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__66662\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56148\,
            lcout => \c0.n5_adj_4302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1374_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63961\,
            in2 => \_gnd_net_\,
            in3 => \N__63507\,
            lcout => \c0.n22577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1484_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47878\,
            in2 => \_gnd_net_\,
            in3 => \N__43604\,
            lcout => \c0.n74_adj_4525\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i11_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47879\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49003\,
            lcout => \c0.FRAME_MATCHER_state_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78695\,
            ce => 'H',
            sr => \N__47850\
        );

    \c0.i1_2_lut_3_lut_adj_1988_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__62253\,
            in1 => \N__74666\,
            in2 => \_gnd_net_\,
            in3 => \N__74470\,
            lcout => \c0.n4_adj_4266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1246_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__74469\,
            in1 => \N__74382\,
            in2 => \N__74674\,
            in3 => \N__49552\,
            lcout => \c0.n23912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14109_2_lut_3_lut_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__53909\,
            in1 => \N__80924\,
            in2 => \_gnd_net_\,
            in3 => \N__49553\,
            lcout => \c0.n3844\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_2030_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001101"
        )
    port map (
            in0 => \N__49554\,
            in1 => \N__53910\,
            in2 => \N__80951\,
            in3 => \N__44277\,
            lcout => OPEN,
            ltout => \c0.n22098_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1286_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__53911\,
            in1 => \N__49827\,
            in2 => \N__44238\,
            in3 => \N__48483\,
            lcout => OPEN,
            ltout => \c0.n63_adj_4305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i0_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__44013\,
            in1 => \N__44235\,
            in2 => \N__44229\,
            in3 => \N__44194\,
            lcout => \c0.FRAME_MATCHER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78707\,
            ce => 'H',
            sr => \N__44995\
        );

    \c0.i1_2_lut_4_lut_adj_1996_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__44109\,
            in1 => \N__44057\,
            in2 => \N__44012\,
            in3 => \N__43530\,
            lcout => \c0.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1906_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__43924\,
            in1 => \N__43869\,
            in2 => \N__49755\,
            in3 => \N__43837\,
            lcout => OPEN,
            ltout => \c0.n24591_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i2_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__43710\,
            in1 => \N__43671\,
            in2 => \N__43638\,
            in3 => \N__43635\,
            lcout => \c0.FRAME_MATCHER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78717\,
            ce => 'H',
            sr => \N__45027\
        );

    \c0.FRAME_MATCHER_state_i15_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43598\,
            in2 => \_gnd_net_\,
            in3 => \N__48979\,
            lcout => \c0.FRAME_MATCHER_state_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78731\,
            ce => 'H',
            sr => \N__43563\
        );

    \c0.FRAME_MATCHER_state_i1_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111011100"
        )
    port map (
            in0 => \N__49786\,
            in1 => \N__43551\,
            in2 => \N__43545\,
            in3 => \N__43532\,
            lcout => \c0.FRAME_MATCHER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78743\,
            ce => 'H',
            sr => \N__45028\
        );

    \c0.FRAME_MATCHER_state_i20_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44314\,
            in2 => \_gnd_net_\,
            in3 => \N__48999\,
            lcout => \c0.FRAME_MATCHER_state_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78756\,
            ce => 'H',
            sr => \N__44292\
        );

    \c0.equal_88_i9_2_lut_3_lut_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__74344\,
            in1 => \N__74480\,
            in2 => \_gnd_net_\,
            in3 => \N__74636\,
            lcout => \c0.n9_adj_4273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i200_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__72860\,
            in1 => \N__76324\,
            in2 => \N__52071\,
            in3 => \N__79483\,
            lcout => \c0.data_in_frame_24_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i65_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__80707\,
            in1 => \N__73596\,
            in2 => \N__61548\,
            in3 => \N__72861\,
            lcout => \c0.data_in_frame_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i215_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69166\,
            in1 => \N__73155\,
            in2 => \N__75989\,
            in3 => \N__79484\,
            lcout => \c0.data_in_frame_26_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i154_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76623\,
            in1 => \N__80398\,
            in2 => \N__63412\,
            in3 => \N__75243\,
            lcout => \c0.data_in_frame_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i82_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__73595\,
            in1 => \N__75244\,
            in2 => \N__69200\,
            in3 => \N__55070\,
            lcout => \c0.data_in_frame_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i9_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__70151\,
            in1 => \N__74069\,
            in2 => \N__80739\,
            in3 => \N__61035\,
            lcout => data_in_frame_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i26_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76622\,
            in1 => \N__70152\,
            in2 => \N__54950\,
            in3 => \N__75242\,
            lcout => \c0.data_in_frame_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1904_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70299\,
            in1 => \N__51336\,
            in2 => \N__61176\,
            in3 => \N__71100\,
            lcout => \c0.n20_adj_4726\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i7_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50401\,
            in1 => \N__44565\,
            in2 => \_gnd_net_\,
            in3 => \N__44513\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i31_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__73153\,
            in1 => \N__50402\,
            in2 => \_gnd_net_\,
            in3 => \N__44466\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__44588\,
            in1 => \N__73154\,
            in2 => \N__50864\,
            in3 => \N__49389\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1929_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111110"
        )
    port map (
            in0 => \N__48594\,
            in1 => \N__61142\,
            in2 => \N__44448\,
            in3 => \N__68217\,
            lcout => \c0.n27_adj_4735\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_2_i3_2_lut_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74659\,
            in2 => \_gnd_net_\,
            in3 => \N__71542\,
            lcout => \c0.n3_adj_4432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_74_i9_2_lut_3_lut_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__74365\,
            in1 => \N__74498\,
            in2 => \_gnd_net_\,
            in3 => \N__74658\,
            lcout => \c0.n9_adj_4601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_2__I_0_2_lut_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47294\,
            in2 => \_gnd_net_\,
            in3 => \N__47012\,
            lcout => \c0.data_out_frame_29__7__N_735\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1362_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47293\,
            in1 => \N__44830\,
            in2 => \N__45323\,
            in3 => \N__44405\,
            lcout => \c0.n22754\,
            ltout => \c0.n22754_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1318_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44363\,
            in1 => \N__45627\,
            in2 => \N__44352\,
            in3 => \N__44808\,
            lcout => \c0.n22243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1298_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47298\,
            in1 => \N__44910\,
            in2 => \N__44802\,
            in3 => \N__45262\,
            lcout => \c0.n10477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i18_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__44880\,
            in1 => \_gnd_net_\,
            in2 => \N__44846\,
            in3 => \N__47720\,
            lcout => encoder0_position_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78718\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1759_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__47013\,
            in1 => \_gnd_net_\,
            in2 => \N__47305\,
            in3 => \N__44831\,
            lcout => \c0.n22641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1316_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47011\,
            in2 => \_gnd_net_\,
            in3 => \N__45184\,
            lcout => \c0.n22583\,
            ltout => \c0.n22583_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1292_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44798\,
            in1 => \N__44769\,
            in2 => \N__44718\,
            in3 => \N__44703\,
            lcout => \c0.n13872\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i20_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__47612\,
            in1 => \_gnd_net_\,
            in2 => \N__44607\,
            in3 => \N__45322\,
            lcout => encoder0_position_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1720_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__61391\,
            in1 => \N__62244\,
            in2 => \_gnd_net_\,
            in3 => \N__75327\,
            lcout => n22101,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__44589\,
            in1 => \N__76154\,
            in2 => \N__50913\,
            in3 => \N__50718\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1315_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45648\,
            in2 => \_gnd_net_\,
            in3 => \N__46954\,
            lcout => \c0.n22252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__3__5474_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__48077\,
            in1 => \N__46031\,
            in2 => \N__45615\,
            in3 => \N__45533\,
            lcout => data_out_frame_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1405_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__45518\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45444\,
            lcout => \c0.n22553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1763_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45392\,
            in1 => \N__46955\,
            in2 => \_gnd_net_\,
            in3 => \N__45321\,
            lcout => \c0.n22689\,
            ltout => \c0.n22689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1338_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45276\,
            in1 => \N__45260\,
            in2 => \N__45192\,
            in3 => \N__45185\,
            lcout => \c0.n10455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46483\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46272\,
            lcout => \c0.n22522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_2048_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46271\,
            in1 => \N__46553\,
            in2 => \N__46827\,
            in3 => \N__46482\,
            lcout => \c0.n20312\,
            ltout => \c0.n20312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1749_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46500\,
            in1 => \N__46879\,
            in2 => \N__45087\,
            in3 => \N__46822\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4674_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__4__5289_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45084\,
            in1 => \N__46704\,
            in2 => \N__45078\,
            in3 => \N__46743\,
            lcout => \c0.data_out_frame_29_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78679\,
            ce => \N__45037\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1275_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46742\,
            in1 => \N__46631\,
            in2 => \_gnd_net_\,
            in3 => \N__46614\,
            lcout => \c0.n20786\,
            ltout => \c0.n20786_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1451_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46542\,
            in3 => \N__46499\,
            lcout => \c0.n9_adj_4494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1344_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46741\,
            in1 => \N__46184\,
            in2 => \N__46485\,
            in3 => \N__46532\,
            lcout => \c0.n21433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_2023_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46183\,
            in1 => \N__46478\,
            in2 => \N__46826\,
            in3 => \N__46740\,
            lcout => \c0.n12590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1655_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46449\,
            in1 => \N__46378\,
            in2 => \N__46362\,
            in3 => \N__46254\,
            lcout => \c0.n10531\,
            ltout => \c0.n10531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_2025_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46823\,
            in1 => \N__46188\,
            in2 => \N__46158\,
            in3 => \N__46744\,
            lcout => \c0.n21451\,
            ltout => \c0.n21451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1346_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46133\,
            in2 => \N__46101\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_frame_29__3__N_1730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__6__5455_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__48186\,
            in1 => \N__46090\,
            in2 => \N__45692\,
            in3 => \N__47484\,
            lcout => data_out_frame_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__6__I_721_2_lut_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46878\,
            in2 => \_gnd_net_\,
            in3 => \N__46825\,
            lcout => \c0.data_out_frame_29__6__N_1538\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1439_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46745\,
            lcout => \c0.n4_adj_4271\,
            ltout => \c0.n4_adj_4271_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1251_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46710\,
            in1 => \N__46703\,
            in2 => \N__46680\,
            in3 => \N__46677\,
            lcout => \data_out_frame_29__3__N_1661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47231\,
            in2 => \_gnd_net_\,
            in3 => \N__46652\,
            lcout => n12904,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_2036_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48768\,
            in2 => \_gnd_net_\,
            in3 => \N__47841\,
            lcout => \c0.n21647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1544_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__61384\,
            in1 => \N__62309\,
            in2 => \_gnd_net_\,
            in3 => \N__61425\,
            lcout => \c0.n22112\,
            ltout => \c0.n22112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i86_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__61582\,
            in1 => \N__69161\,
            in2 => \N__46635\,
            in3 => \N__79791\,
            lcout => \c0.data_in_frame_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i166_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__80417\,
            in1 => \N__79984\,
            in2 => \N__79796\,
            in3 => \N__56143\,
            lcout => \c0.data_in_frame_20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i151_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__73214\,
            in1 => \N__80418\,
            in2 => \N__61897\,
            in3 => \N__69162\,
            lcout => \c0.data_in_frame_18_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i102_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__79787\,
            in1 => \N__73519\,
            in2 => \N__55742\,
            in3 => \N__79985\,
            lcout => \c0.data_in_frame_12_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i124_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__73518\,
            in1 => \N__80867\,
            in2 => \N__65426\,
            in3 => \N__77128\,
            lcout => \c0.data_in_frame_15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i20_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50454\,
            in1 => \N__48680\,
            in2 => \_gnd_net_\,
            in3 => \N__46906\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_2011_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__74673\,
            in1 => \N__74520\,
            in2 => \N__74386\,
            in3 => \N__61424\,
            lcout => \c0.n22099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1783_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__66099\,
            in1 => \N__66569\,
            in2 => \_gnd_net_\,
            in3 => \N__65406\,
            lcout => OPEN,
            ltout => \c0.n82_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i61_4_lut_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56056\,
            in1 => \N__66637\,
            in2 => \N__46887\,
            in3 => \N__72049\,
            lcout => \c0.n142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i146_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__72050\,
            in1 => \N__75110\,
            in2 => \N__69199\,
            in3 => \N__80420\,
            lcout => \c0.data_in_frame_18_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i118_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__62396\,
            in1 => \N__59190\,
            in2 => \_gnd_net_\,
            in3 => \N__79776\,
            lcout => data_in_frame_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i150_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__79777\,
            in1 => \N__80419\,
            in2 => \N__56072\,
            in3 => \N__69157\,
            lcout => \c0.data_in_frame_18_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i122_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__80899\,
            in1 => \N__73521\,
            in2 => \N__62459\,
            in3 => \N__75111\,
            lcout => \c0.data_in_frame_15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1925_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49196\,
            in2 => \_gnd_net_\,
            in3 => \N__47837\,
            lcout => \c0.n21629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_adj_1166_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__47234\,
            in1 => \N__49718\,
            in2 => \_gnd_net_\,
            in3 => \N__49657\,
            lcout => OPEN,
            ltout => \c0.rx.n17834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i11373_3_lut_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__50153\,
            in1 => \_gnd_net_\,
            in2 => \N__47154\,
            in3 => \N__47151\,
            lcout => n14988,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1445_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__67884\,
            in1 => \N__64133\,
            in2 => \_gnd_net_\,
            in3 => \N__56632\,
            lcout => \c0.n17_adj_4483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1867_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__56223\,
            in1 => \N__62296\,
            in2 => \_gnd_net_\,
            in3 => \N__75301\,
            lcout => n22103,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i5_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47057\,
            in1 => \N__60438\,
            in2 => \_gnd_net_\,
            in3 => \N__47347\,
            lcout => control_mode_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1520_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62397\,
            in2 => \_gnd_net_\,
            in3 => \N__62458\,
            lcout => \c0.n4_adj_4352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i1_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47007\,
            in1 => \N__51237\,
            in2 => \_gnd_net_\,
            in3 => \N__47343\,
            lcout => control_mode_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i3_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46953\,
            in2 => \N__47352\,
            in3 => \N__51480\,
            lcout => control_mode_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i134_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__79785\,
            in1 => \N__80421\,
            in2 => \N__62526\,
            in3 => \N__72990\,
            lcout => \c0.data_in_frame_16_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i14_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47723\,
            in1 => \N__47520\,
            in2 => \_gnd_net_\,
            in3 => \N__47468\,
            lcout => encoder0_position_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__47430\,
            in1 => \N__78979\,
            in2 => \N__50912\,
            in3 => \N__49369\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1442_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51944\,
            in1 => \N__63942\,
            in2 => \N__47409\,
            in3 => \N__51887\,
            lcout => OPEN,
            ltout => \c0.n26_adj_4480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_1447_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47739\,
            in1 => \N__47388\,
            in2 => \N__47376\,
            in3 => \N__76710\,
            lcout => \c0.n24539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1507_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__47373\,
            in1 => \N__67680\,
            in2 => \N__56925\,
            in3 => \N__49533\,
            lcout => OPEN,
            ltout => \c0.n34_adj_4546_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1522_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__47241\,
            in1 => \N__56946\,
            in2 => \N__47355\,
            in3 => \N__60000\,
            lcout => n24622,
            ltout => \n24622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i2_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__57270\,
            in1 => \_gnd_net_\,
            in2 => \N__47319\,
            in3 => \N__47277\,
            lcout => control_mode_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20968_4_lut_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100000000"
        )
    port map (
            in0 => \N__51888\,
            in1 => \N__49431\,
            in2 => \N__59670\,
            in3 => \N__47247\,
            lcout => \c0.n24733\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i157_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__80422\,
            in1 => \N__76682\,
            in2 => \N__71967\,
            in3 => \N__56185\,
            lcout => \c0.data_in_frame_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i238_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__49446\,
            in1 => \N__56487\,
            in2 => \N__79800\,
            in3 => \N__75337\,
            lcout => \c0.data_in_frame_29_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1739_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__75611\,
            in1 => \N__76749\,
            in2 => \N__75576\,
            in3 => \N__63609\,
            lcout => \c0.n18_adj_4485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i199_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__73207\,
            in1 => \N__72981\,
            in2 => \N__67150\,
            in3 => \N__79361\,
            lcout => \c0.data_in_frame_24_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i207_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__79359\,
            in1 => \N__74220\,
            in2 => \N__59629\,
            in3 => \N__73209\,
            lcout => \c0.data_in_frame_25_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i193_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__80738\,
            in1 => \N__72980\,
            in2 => \N__78017\,
            in3 => \N__79360\,
            lcout => \c0.data_in_frame_24_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i135_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__72979\,
            in1 => \N__80423\,
            in2 => \N__58930\,
            in3 => \N__73208\,
            lcout => \c0.data_in_frame_16_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1443_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56814\,
            in1 => \N__59578\,
            in2 => \N__63877\,
            in3 => \N__67248\,
            lcout => \c0.n24384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i196_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__76912\,
            in1 => \N__72942\,
            in2 => \N__59587\,
            in3 => \N__79356\,
            lcout => \c0.data_in_frame_24_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1660_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__56241\,
            in1 => \N__62319\,
            in2 => \_gnd_net_\,
            in3 => \N__61433\,
            lcout => \c0.n22134\,
            ltout => \c0.n22134_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i222_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__76694\,
            in1 => \N__79792\,
            in2 => \N__47898\,
            in3 => \N__56886\,
            lcout => \c0.data_in_frame_27_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i214_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__79355\,
            in1 => \N__79647\,
            in2 => \N__63878\,
            in3 => \N__69227\,
            lcout => \c0.data_in_frame_26_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i209_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__69226\,
            in1 => \N__56588\,
            in2 => \N__80671\,
            in3 => \N__79357\,
            lcout => \c0.data_in_frame_26_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i197_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__79354\,
            in1 => \N__71939\,
            in2 => \N__72977\,
            in3 => \N__67249\,
            lcout => \c0.data_in_frame_24_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i223_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__76695\,
            in1 => \N__73210\,
            in2 => \N__56853\,
            in3 => \N__79358\,
            lcout => \c0.data_in_frame_27_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1949_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47883\,
            in2 => \_gnd_net_\,
            in3 => \N__47829\,
            lcout => \c0.n21633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i232_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__80093\,
            in1 => \N__76317\,
            in2 => \N__52241\,
            in3 => \N__79365\,
            lcout => \c0.data_in_frame_28_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1198_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48416\,
            in2 => \_gnd_net_\,
            in3 => \N__47828\,
            lcout => \c0.n21651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i218_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__76687\,
            in1 => \N__75185\,
            in2 => \N__64139\,
            in3 => \N__79364\,
            lcout => \c0.data_in_frame_27_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19136_4_lut_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__49845\,
            in1 => \N__52408\,
            in2 => \N__48528\,
            in3 => \N__53915\,
            lcout => \c0.n5024\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1543_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__48482\,
            in1 => \N__48450\,
            in2 => \N__48432\,
            in3 => \N__53803\,
            lcout => \c0.n2119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i31_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48412\,
            in2 => \_gnd_net_\,
            in3 => \N__48980\,
            lcout => \c0.FRAME_MATCHER_state_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78744\,
            ce => 'H',
            sr => \N__48390\
        );

    \c0.select_367_Select_4_i3_2_lut_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52374\,
            in2 => \_gnd_net_\,
            in3 => \N__71553\,
            lcout => \c0.n3_adj_4428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_3_lut_adj_1941_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__60714\,
            in1 => \N__60588\,
            in2 => \_gnd_net_\,
            in3 => \N__49863\,
            lcout => \FRAME_MATCHER_state_31_N_2975_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1654_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48710\,
            in1 => \N__47904\,
            in2 => \N__64458\,
            in3 => \N__48534\,
            lcout => OPEN,
            ltout => \c0.n22_adj_4643_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1674_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55184\,
            in1 => \N__55508\,
            in2 => \N__47910\,
            in3 => \N__60548\,
            lcout => \c0.n24433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1644_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55021\,
            in1 => \N__50984\,
            in2 => \N__61541\,
            in3 => \N__50971\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4639_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1649_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55069\,
            in1 => \N__48744\,
            in2 => \N__47907\,
            in3 => \N__50945\,
            lcout => \c0.n13_adj_4640\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_1677_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57942\,
            in2 => \_gnd_net_\,
            in3 => \N__61031\,
            lcout => \c0.n12_adj_4657\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1607_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50972\,
            in1 => \N__55020\,
            in2 => \N__50988\,
            in3 => \N__50944\,
            lcout => \c0.n23666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_adj_1875_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55220\,
            in1 => \N__51085\,
            in2 => \N__57376\,
            in3 => \N__64764\,
            lcout => \c0.n20_adj_4642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i10_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__74066\,
            in1 => \N__70172\,
            in2 => \N__75254\,
            in3 => \N__51207\,
            lcout => data_in_frame_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i11_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__70170\,
            in1 => \N__74067\,
            in2 => \N__57244\,
            in3 => \N__79189\,
            lcout => data_in_frame_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i47_3_lut_4_lut_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64614\,
            in1 => \N__55664\,
            in2 => \N__55746\,
            in3 => \N__69903\,
            lcout => \c0.n128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1735_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50969\,
            in2 => \_gnd_net_\,
            in3 => \N__50943\,
            lcout => \c0.n5_adj_4268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i46_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50970\,
            in1 => \N__79628\,
            in2 => \_gnd_net_\,
            in3 => \N__69437\,
            lcout => data_in_frame_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i29_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__70171\,
            in1 => \N__76550\,
            in2 => \N__50949\,
            in3 => \N__71957\,
            lcout => \c0.data_in_frame_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1831_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51206\,
            in2 => \_gnd_net_\,
            in3 => \N__51418\,
            lcout => \c0.n22626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_adj_1603_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57228\,
            in1 => \N__51564\,
            in2 => \_gnd_net_\,
            in3 => \N__50942\,
            lcout => \c0.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i30_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__76548\,
            in1 => \N__70153\,
            in2 => \N__79677\,
            in3 => \N__51573\,
            lcout => \c0.data_in_frame_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1645_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54936\,
            in1 => \N__51211\,
            in2 => \_gnd_net_\,
            in3 => \N__57484\,
            lcout => \c0.n23305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_adj_1594_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71099\,
            in1 => \N__61030\,
            in2 => \N__60409\,
            in3 => \N__58012\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4607_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1832_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48542\,
            in1 => \N__60305\,
            in2 => \N__48558\,
            in3 => \N__48554\,
            lcout => \c0.data_out_frame_0__7__N_2626\,
            ltout => \c0.data_out_frame_0__7__N_2626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i32_4_lut_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48555\,
            in1 => \N__51335\,
            in2 => \N__48546\,
            in3 => \N__57564\,
            lcout => \c0.n88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_1830_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57232\,
            in2 => \_gnd_net_\,
            in3 => \N__60490\,
            lcout => \c0.n30_adj_4585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_4_lut_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57233\,
            in1 => \N__60386\,
            in2 => \N__60533\,
            in3 => \N__58013\,
            lcout => \c0.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_2_lut_3_lut_4_lut_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48543\,
            in1 => \N__51212\,
            in2 => \N__51465\,
            in3 => \N__55331\,
            lcout => \c0.n39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i49_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__57593\,
            in1 => \N__80655\,
            in2 => \_gnd_net_\,
            in3 => \N__68442\,
            lcout => data_in_frame_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1243_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51562\,
            in2 => \_gnd_net_\,
            in3 => \N__57592\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1244_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60835\,
            in1 => \N__60378\,
            in2 => \N__48573\,
            in3 => \N__51439\,
            lcout => \c0.n13223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1918_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__64346\,
            in1 => \N__61194\,
            in2 => \N__51099\,
            in3 => \N__61860\,
            lcout => \c0.n28_adj_4731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i31_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__76549\,
            in1 => \N__60850\,
            in2 => \N__70186\,
            in3 => \N__73156\,
            lcout => \c0.data_in_frame_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i14_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__79587\,
            in1 => \N__74104\,
            in2 => \N__60408\,
            in3 => \N__70178\,
            lcout => data_in_frame_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1860_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60834\,
            in1 => \N__60377\,
            in2 => \N__57488\,
            in3 => \N__51223\,
            lcout => \c0.n15_adj_4710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i27_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__79190\,
            in1 => \N__70174\,
            in2 => \N__76599\,
            in3 => \N__57483\,
            lcout => \c0.data_in_frame_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i24_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__76148\,
            in1 => \N__70149\,
            in2 => \N__64755\,
            in3 => \N__69117\,
            lcout => \c0.data_in_frame_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i56_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__68422\,
            in1 => \N__76149\,
            in2 => \_gnd_net_\,
            in3 => \N__64873\,
            lcout => data_in_frame_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i48_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__57638\,
            in1 => \N__76153\,
            in2 => \_gnd_net_\,
            in3 => \N__69411\,
            lcout => data_in_frame_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i80_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__76152\,
            in1 => \N__73658\,
            in2 => \N__55023\,
            in3 => \N__74021\,
            lcout => \c0.data_in_frame_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1218_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__49238\,
            in1 => \N__49303\,
            in2 => \N__48684\,
            in3 => \N__48636\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1843_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57637\,
            in2 => \_gnd_net_\,
            in3 => \N__48743\,
            lcout => \c0.n6_adj_4704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1914_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \N__51159\,
            in1 => \N__57782\,
            in2 => \N__51015\,
            in3 => \N__64377\,
            lcout => \c0.n20_adj_4729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i47_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48739\,
            in1 => \N__69410\,
            in2 => \_gnd_net_\,
            in3 => \N__73201\,
            lcout => data_in_frame_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1844_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51574\,
            in1 => \N__58199\,
            in2 => \N__48588\,
            in3 => \N__60535\,
            lcout => \c0.n14016\,
            ltout => \c0.n14016_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_adj_1640_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61552\,
            in2 => \N__48579\,
            in3 => \N__55455\,
            lcout => \c0.n13329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_1826_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__60534\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48731\,
            lcout => \c0.n20\,
            ltout => \c0.n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1347_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55512\,
            in1 => \N__57636\,
            in2 => \N__48576\,
            in3 => \N__48697\,
            lcout => \c0.n4_adj_4333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__60536\,
            in1 => \N__48732\,
            in2 => \N__71187\,
            in3 => \N__55513\,
            lcout => \c0.n23_adj_4590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i114_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__75255\,
            in1 => \N__59207\,
            in2 => \_gnd_net_\,
            in3 => \N__55429\,
            lcout => data_in_frame_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i62_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__79626\,
            in1 => \N__70147\,
            in2 => \N__64450\,
            in3 => \N__80920\,
            lcout => \c0.data_in_frame_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1717_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65184\,
            in2 => \_gnd_net_\,
            in3 => \N__65073\,
            lcout => \c0.n5_adj_4443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i55_3_lut_4_lut_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62614\,
            in1 => \N__59259\,
            in2 => \N__61987\,
            in3 => \N__51275\,
            lcout => \c0.n136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i128_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__80919\,
            in1 => \N__73669\,
            in2 => \N__61991\,
            in3 => \N__76151\,
            lcout => \c0.data_in_frame_15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i101_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__73668\,
            in1 => \N__59010\,
            in2 => \N__80099\,
            in3 => \N__71762\,
            lcout => \c0.data_in_frame_12_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i113_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__80575\,
            in1 => \N__59206\,
            in2 => \_gnd_net_\,
            in3 => \N__58614\,
            lcout => data_in_frame_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i64_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__76150\,
            in1 => \N__70148\,
            in2 => \N__48711\,
            in3 => \N__80921\,
            lcout => \c0.data_in_frame_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__71761\,
            in1 => \N__49572\,
            in2 => \N__50904\,
            in3 => \N__49385\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i7_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49186\,
            in2 => \_gnd_net_\,
            in3 => \N__49007\,
            lcout => \c0.FRAME_MATCHER_state_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78697\,
            ce => 'H',
            sr => \N__49170\
        );

    \c0.i6_4_lut_adj_1597_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57663\,
            in1 => \N__61553\,
            in2 => \N__59011\,
            in3 => \N__58892\,
            lcout => \c0.n16_adj_4608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1202_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__55727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59001\,
            lcout => \c0.n13186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1901_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__64884\,
            in1 => \N__57816\,
            in2 => \N__57671\,
            in3 => \N__64638\,
            lcout => \c0.n25_adj_4723\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64883\,
            in2 => \_gnd_net_\,
            in3 => \N__68127\,
            lcout => \c0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1900_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__64834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__64737\,
            lcout => \c0.n7_adj_4337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1973_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49143\,
            in1 => \N__49107\,
            in2 => \N__49083\,
            in3 => \N__48766\,
            lcout => \c0.n22049\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i27_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48767\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49011\,
            lcout => \c0.FRAME_MATCHER_state_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78681\,
            ce => 'H',
            sr => \N__48753\
        );

    \c0.i42_4_lut_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72689\,
            in1 => \N__72154\,
            in2 => \N__58937\,
            in3 => \N__59105\,
            lcout => \c0.n123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_9_i3_2_lut_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__71519\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52776\,
            lcout => \c0.n3_adj_4418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1348_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62445\,
            in2 => \_gnd_net_\,
            in3 => \N__65405\,
            lcout => \c0.n22463\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i3_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50480\,
            in1 => \N__49272\,
            in2 => \_gnd_net_\,
            in3 => \N__49237\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_1701_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62379\,
            in1 => \N__59018\,
            in2 => \_gnd_net_\,
            in3 => \N__58775\,
            lcout => \c0.n15_adj_4301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1919_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51291\,
            in1 => \N__58618\,
            in2 => \N__70482\,
            in3 => \N__62854\,
            lcout => \c0.n10_adj_4732\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1231_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49320\,
            in1 => \N__65460\,
            in2 => \N__69669\,
            in3 => \N__51279\,
            lcout => \c0.n21491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1920_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62931\,
            in1 => \N__64662\,
            in2 => \N__49215\,
            in3 => \N__68556\,
            lcout => OPEN,
            ltout => \c0.n26_adj_4733_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1989_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68883\,
            in1 => \N__65538\,
            in2 => \N__49206\,
            in3 => \N__68593\,
            lcout => \c0.n20409\,
            ltout => \c0.n20409_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1232_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49203\,
            in3 => \N__63542\,
            lcout => \c0.n22716\,
            ltout => \c0.n22716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_2042_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51773\,
            in1 => \N__56139\,
            in2 => \N__49323\,
            in3 => \N__59742\,
            lcout => \c0.n21389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1542_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56193\,
            in2 => \_gnd_net_\,
            in3 => \N__58833\,
            lcout => \c0.n6_adj_4577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58619\,
            in1 => \N__66228\,
            in2 => \_gnd_net_\,
            in3 => \N__60063\,
            lcout => \c0.n8_adj_4248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i26_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__75028\,
            in1 => \N__50473\,
            in2 => \_gnd_net_\,
            in3 => \N__49302\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i171_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__78978\,
            in1 => \N__67620\,
            in2 => \_gnd_net_\,
            in3 => \N__51729\,
            lcout => data_in_frame_21_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1952_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__52480\,
            in1 => \N__52410\,
            in2 => \_gnd_net_\,
            in3 => \N__52568\,
            lcout => \c0.n12989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i148_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__80318\,
            in1 => \N__77102\,
            in2 => \N__69225\,
            in3 => \N__66650\,
            lcout => \c0.data_in_frame_18_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i172_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__67621\,
            in1 => \N__77101\,
            in2 => \_gnd_net_\,
            in3 => \N__65884\,
            lcout => data_in_frame_21_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_14_i3_2_lut_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52955\,
            in2 => \_gnd_net_\,
            in3 => \N__71482\,
            lcout => \c0.n3_adj_4408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i168_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__80096\,
            in1 => \N__76389\,
            in2 => \N__56370\,
            in3 => \N__80319\,
            lcout => \c0.data_in_frame_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_16_i3_2_lut_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53054\,
            in2 => \_gnd_net_\,
            in3 => \N__71483\,
            lcout => \c0.n3_adj_4404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1642_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72219\,
            in2 => \_gnd_net_\,
            in3 => \N__72161\,
            lcout => \c0.n13756\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1478_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59876\,
            in2 => \_gnd_net_\,
            in3 => \N__56515\,
            lcout => \c0.n15_adj_4508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i25_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50484\,
            in1 => \N__80508\,
            in2 => \_gnd_net_\,
            in3 => \N__49422\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1536_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58689\,
            in1 => \N__66579\,
            in2 => \N__61962\,
            in3 => \N__66369\,
            lcout => \c0.n23718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1365_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56354\,
            in2 => \_gnd_net_\,
            in3 => \N__63560\,
            lcout => \c0.n15_adj_4344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1390_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__56815\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__77273\,
            lcout => \c0.n5_adj_4370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__49349\,
            in1 => \N__80509\,
            in2 => \N__50911\,
            in3 => \N__49378\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__75027\,
            in1 => \N__49350\,
            in2 => \N__50910\,
            in3 => \N__50719\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1401_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__49332\,
            in1 => \N__66654\,
            in2 => \N__62982\,
            in3 => \N__56736\,
            lcout => \c0.n20_adj_4441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1541_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51810\,
            in1 => \N__49473\,
            in2 => \N__52097\,
            in3 => \N__56738\,
            lcout => \c0.n14_adj_4576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1369_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51777\,
            in1 => \N__59493\,
            in2 => \N__49494\,
            in3 => \N__61934\,
            lcout => OPEN,
            ltout => \c0.n12_adj_4348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1486_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66897\,
            in1 => \N__63306\,
            in2 => \N__49476\,
            in3 => \N__66710\,
            lcout => \c0.n8_adj_4526\,
            ltout => \c0.n8_adj_4526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1489_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56737\,
            in1 => \N__52205\,
            in2 => \N__49467\,
            in3 => \N__51809\,
            lcout => \c0.n14_adj_4528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1496_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__76828\,
            in2 => \_gnd_net_\,
            in3 => \N__63241\,
            lcout => \c0.n9_adj_4536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1498_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56276\,
            in1 => \N__49464\,
            in2 => \N__59875\,
            in3 => \N__49458\,
            lcout => \c0.n24547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1550_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51870\,
            in1 => \N__51945\,
            in2 => \N__56649\,
            in3 => \N__49452\,
            lcout => \c0.n24098\,
            ltout => \c0.n24098_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1446_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__49445\,
            in1 => \N__52035\,
            in2 => \N__49434\,
            in3 => \N__51897\,
            lcout => \c0.n10_adj_4484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_adj_1736_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__77291\,
            in1 => \N__76833\,
            in2 => \N__59628\,
            in3 => \N__56752\,
            lcout => \c0.n20_adj_4512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i170_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__66426\,
            in1 => \N__75113\,
            in2 => \_gnd_net_\,
            in3 => \N__67644\,
            lcout => data_in_frame_21_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1370_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66425\,
            in2 => \_gnd_net_\,
            in3 => \N__51778\,
            lcout => \c0.n5_adj_4349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_1435_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56670\,
            in1 => \N__49500\,
            in2 => \N__49523\,
            in3 => \N__59524\,
            lcout => OPEN,
            ltout => \c0.n52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i30_4_lut_adj_1500_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59557\,
            in1 => \N__72371\,
            in2 => \N__49539\,
            in3 => \N__67038\,
            lcout => \c0.n64_adj_4539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_1513_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59556\,
            in2 => \_gnd_net_\,
            in3 => \N__59525\,
            lcout => OPEN,
            ltout => \c0.n47_adj_4537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1497_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57076\,
            in1 => \N__49508\,
            in2 => \N__49536\,
            in3 => \N__56893\,
            lcout => \c0.n24581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i234_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__75112\,
            in1 => \N__56461\,
            in2 => \N__49524\,
            in3 => \N__75407\,
            lcout => \c0.data_in_frame_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i239_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__75406\,
            in1 => \N__73346\,
            in2 => \N__56479\,
            in3 => \N__49509\,
            lcout => \c0.data_in_frame_29_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1704_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67121\,
            in1 => \N__52028\,
            in2 => \N__57021\,
            in3 => \N__51998\,
            lcout => \c0.n20793\,
            ltout => \c0.n20793_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63018\,
            in1 => \N__59912\,
            in2 => \N__49557\,
            in3 => \N__72370\,
            lcout => \c0.n70_adj_4514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_4_lut_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66430\,
            in1 => \N__56369\,
            in2 => \N__56411\,
            in3 => \N__51779\,
            lcout => \c0.n14_adj_4529\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i216_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__79362\,
            in1 => \N__69224\,
            in2 => \N__76365\,
            in3 => \N__67296\,
            lcout => \c0.data_in_frame_26_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i167_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__73298\,
            in1 => \N__56406\,
            in2 => \N__80100\,
            in3 => \N__80424\,
            lcout => \c0.data_in_frame_20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1277_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__62316\,
            in1 => \N__52407\,
            in2 => \_gnd_net_\,
            in3 => \N__49844\,
            lcout => \c0.n12927\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i211_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69223\,
            in1 => \N__79173\,
            in2 => \N__66807\,
            in3 => \N__79363\,
            lcout => \c0.data_in_frame_26_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_15_i3_2_lut_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__71348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53006\,
            lcout => \c0.n3_adj_4406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_11_i3_2_lut_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52836\,
            in2 => \_gnd_net_\,
            in3 => \N__71347\,
            lcout => \c0.n3_adj_4414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_6_i3_2_lut_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__71351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52575\,
            lcout => \c0.n3_adj_4424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i204_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__74216\,
            in1 => \N__76945\,
            in2 => \N__52204\,
            in3 => \N__79421\,
            lcout => \c0.data_in_frame_25_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_23_i3_2_lut_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__71350\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53309\,
            lcout => \c0.n3_adj_4390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_22_i3_2_lut_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53271\,
            in2 => \_gnd_net_\,
            in3 => \N__71349\,
            lcout => \c0.n3_adj_4392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_24_i3_2_lut_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53346\,
            in2 => \_gnd_net_\,
            in3 => \N__71372\,
            lcout => \c0.n3_adj_4388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1953_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__52409\,
            in1 => \N__52485\,
            in2 => \_gnd_net_\,
            in3 => \N__52561\,
            lcout => \c0.n12973\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_adj_1276_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49857\,
            in1 => \N__52140\,
            in2 => \N__52215\,
            in3 => \N__52257\,
            lcout => \c0.n13043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_1267_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__53409\,
            in1 => \N__52835\,
            in2 => \N__53058\,
            in3 => \N__53270\,
            lcout => \c0.n41_adj_4292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19124_2_lut_3_lut_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__53908\,
            in1 => \N__49830\,
            in2 => \_gnd_net_\,
            in3 => \N__49787\,
            lcout => \c0.n22885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_31_i3_2_lut_LC_17_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53881\,
            in2 => \_gnd_net_\,
            in3 => \N__71536\,
            lcout => \c0.n3_adj_4373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_102_i4_2_lut_LC_18_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49740\,
            in2 => \_gnd_net_\,
            in3 => \N__49662\,
            lcout => n4,
            ltout => \n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_18_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__79542\,
            in1 => \N__50909\,
            in2 => \N__50736\,
            in3 => \N__50733\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_18_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__50234\,
            in1 => \N__49943\,
            in2 => \N__50184\,
            in3 => \N__50679\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_2_lut_LC_18_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50198\,
            in2 => \_gnd_net_\,
            in3 => \N__50233\,
            lcout => \c0.n161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1887_LC_18_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50664\,
            in1 => \N__50634\,
            in2 => \N__50598\,
            in3 => \N__50541\,
            lcout => \c0.n21_adj_4719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_18_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50235\,
            lcout => \c0.FRAME_MATCHER_rx_data_ready_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i21281_2_lut_3_lut_LC_18_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__50179\,
            in1 => \N__50055\,
            in2 => \_gnd_net_\,
            in3 => \N__49942\,
            lcout => \c0.rx.n22094\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_adj_1940_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__50994\,
            in1 => \N__51000\,
            in2 => \N__59949\,
            in3 => \N__60327\,
            lcout => \c0.n46_adj_4739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_99_i9_2_lut_3_lut_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__74625\,
            in1 => \N__74288\,
            in2 => \_gnd_net_\,
            in3 => \N__74499\,
            lcout => \c0.n9_adj_4563\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_5_i3_2_lut_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52455\,
            in2 => \_gnd_net_\,
            in3 => \N__71545\,
            lcout => \c0.n3_adj_4426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i59_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__80871\,
            in1 => \N__70173\,
            in2 => \N__70741\,
            in3 => \N__79107\,
            lcout => \c0.data_in_frame_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_1933_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__64272\,
            in1 => \N__71032\,
            in2 => \N__68555\,
            in3 => \N__51219\,
            lcout => \c0.n39_adj_4737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1932_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__57243\,
            in1 => \N__51460\,
            in2 => \N__61064\,
            in3 => \N__58043\,
            lcout => \c0.n38_adj_4736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1663_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60229\,
            in1 => \N__51424\,
            in2 => \_gnd_net_\,
            in3 => \N__51216\,
            lcout => \c0.n4_adj_4267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51217\,
            in1 => \N__57930\,
            in2 => \N__51447\,
            in3 => \N__60230\,
            lcout => \c0.n23562\,
            ltout => \c0.n23562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__50941\,
            in1 => \_gnd_net_\,
            in2 => \N__50976\,
            in3 => \N__50973\,
            lcout => \c0.n13280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_adj_1837_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55322\,
            in2 => \_gnd_net_\,
            in3 => \N__57235\,
            lcout => \c0.n22_adj_4647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i28_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__77065\,
            in1 => \N__76595\,
            in2 => \N__57949\,
            in3 => \N__70169\,
            lcout => \c0.data_in_frame_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1851_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50940\,
            in2 => \_gnd_net_\,
            in3 => \N__57234\,
            lcout => \c0.n22511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1722_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57236\,
            in1 => \N__57507\,
            in2 => \N__60239\,
            in3 => \N__51021\,
            lcout => \c0.n13141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i16_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__70168\,
            in1 => \N__74145\,
            in2 => \N__71078\,
            in3 => \N__76285\,
            lcout => data_in_frame_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_4_lut_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55332\,
            in1 => \N__51420\,
            in2 => \N__57535\,
            in3 => \N__51218\,
            lcout => \c0.n18_adj_4228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_3_lut_4_lut_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71031\,
            in1 => \N__56013\,
            in2 => \N__60545\,
            in3 => \N__51136\,
            lcout => \c0.n23_adj_4648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_3_lut_4_lut_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60387\,
            in1 => \N__71030\,
            in2 => \N__72414\,
            in3 => \N__58014\,
            lcout => \c0.n63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_adj_1593_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55124\,
            in1 => \N__51613\,
            in2 => \_gnd_net_\,
            in3 => \N__55980\,
            lcout => \c0.n42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1853_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51563\,
            in1 => \N__60507\,
            in2 => \_gnd_net_\,
            in3 => \N__51419\,
            lcout => \c0.n22160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i12_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__77129\,
            in1 => \N__74179\,
            in2 => \N__51446\,
            in3 => \N__70179\,
            lcout => data_in_frame_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78771\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60511\,
            in2 => \_gnd_net_\,
            in3 => \N__60385\,
            lcout => \c0.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i15_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__70138\,
            in1 => \N__74068\,
            in2 => \N__58055\,
            in3 => \N__73349\,
            lcout => data_in_frame_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i13_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__71915\,
            in1 => \N__74051\,
            in2 => \N__60546\,
            in3 => \N__70140\,
            lcout => data_in_frame_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_adj_1993_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69728\,
            in1 => \N__61263\,
            in2 => \N__71220\,
            in3 => \N__71077\,
            lcout => \c0.n44_adj_4744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i63_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__73348\,
            in1 => \N__70139\,
            in2 => \N__57308\,
            in3 => \N__80888\,
            lcout => \c0.data_in_frame_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_1666_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68545\,
            in1 => \N__68126\,
            in2 => \N__67944\,
            in3 => \N__51044\,
            lcout => \c0.n13_adj_4584\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i117_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__71914\,
            in1 => \N__59208\,
            in2 => \_gnd_net_\,
            in3 => \N__55919\,
            lcout => data_in_frame_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_1263_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51150\,
            in1 => \N__51117\,
            in2 => \N__55383\,
            in3 => \N__61302\,
            lcout => OPEN,
            ltout => \c0.n38_adj_4285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51030\,
            in1 => \N__51054\,
            in2 => \N__51057\,
            in3 => \N__70233\,
            lcout => \c0.n24527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_2_lut_3_lut_4_lut_adj_2029_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51233\,
            in1 => \N__57563\,
            in2 => \N__51464\,
            in3 => \N__51138\,
            lcout => \c0.n26_adj_4289\,
            ltout => \c0.n26_adj_4289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_3_lut_4_lut_adj_1622_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51029\,
            in1 => \N__57721\,
            in2 => \N__51048\,
            in3 => \N__58169\,
            lcout => \c0.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_2_lut_3_lut_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__64839\,
            in1 => \N__64724\,
            in2 => \_gnd_net_\,
            in3 => \N__51045\,
            lcout => \c0.n20_adj_4290\,
            ltout => \c0.n20_adj_4290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_2_lut_3_lut_4_lut_adj_2026_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57562\,
            in1 => \N__51448\,
            in2 => \N__51240\,
            in3 => \N__51232\,
            lcout => \c0.n51\,
            ltout => \c0.n51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_3_lut_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__51149\,
            in1 => \_gnd_net_\,
            in2 => \N__51141\,
            in3 => \N__51137\,
            lcout => \c0.n56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_2_lut_3_lut_4_lut_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57381\,
            in1 => \N__55221\,
            in2 => \N__51108\,
            in3 => \N__64677\,
            lcout => \c0.n102\,
            ltout => \c0.n102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_3_lut_adj_1261_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55430\,
            in2 => \N__51120\,
            in3 => \N__64988\,
            lcout => \c0.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__70551\,
            in1 => \N__58751\,
            in2 => \_gnd_net_\,
            in3 => \N__58967\,
            lcout => \c0.n16_adj_4256\,
            ltout => \c0.n16_adj_4256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i45_4_lut_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51063\,
            in1 => \N__54984\,
            in2 => \N__51111\,
            in3 => \N__69800\,
            lcout => \c0.n126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_1646_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__55185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__64733\,
            lcout => \c0.n9_adj_4279\,
            ltout => \c0.n9_adj_4279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51092\,
            in1 => \N__55242\,
            in2 => \N__51069\,
            in3 => \N__64440\,
            lcout => \c0.n23574\,
            ltout => \c0.n23574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_4_lut_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55186\,
            in1 => \N__70352\,
            in2 => \N__51066\,
            in3 => \N__64606\,
            lcout => \c0.n11_adj_4257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1995_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69898\,
            in1 => \N__60159\,
            in2 => \N__64239\,
            in3 => \N__64017\,
            lcout => \c0.n41_adj_4745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_3_lut_4_lut_adj_2045_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70353\,
            in1 => \N__51328\,
            in2 => \N__69902\,
            in3 => \N__57537\,
            lcout => \c0.n38_adj_4573\,
            ltout => \c0.n38_adj_4573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_3_lut_4_lut_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58419\,
            in1 => \N__64347\,
            in2 => \N__51312\,
            in3 => \N__70298\,
            lcout => OPEN,
            ltout => \c0.n43_adj_4574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_adj_2009_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51309\,
            in1 => \N__67998\,
            in2 => \N__51300\,
            in3 => \N__51297\,
            lcout => \c0.n24048\,
            ltout => \c0.n24048_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_3_lut_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65964\,
            in2 => \N__51282\,
            in3 => \N__56043\,
            lcout => \c0.n109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i53_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__71816\,
            in1 => \N__68441\,
            in2 => \_gnd_net_\,
            in3 => \N__65193\,
            lcout => data_in_frame_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78722\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1923_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111101"
        )
    port map (
            in0 => \N__64613\,
            in1 => \N__57579\,
            in2 => \N__51264\,
            in3 => \N__58373\,
            lcout => \c0.n29_adj_4734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1829_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55125\,
            in2 => \_gnd_net_\,
            in3 => \N__55976\,
            lcout => \c0.n7_adj_4221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i35_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__79203\,
            in1 => \N__70078\,
            in2 => \N__80098\,
            in3 => \N__65069\,
            lcout => \c0.data_in_frame_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1653_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58137\,
            in1 => \N__64409\,
            in2 => \_gnd_net_\,
            in3 => \N__58080\,
            lcout => \c0.n16_adj_4641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i32_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__76315\,
            in1 => \N__76612\,
            in2 => \N__58090\,
            in3 => \N__70079\,
            lcout => \c0.data_in_frame_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1651_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65068\,
            in1 => \N__58079\,
            in2 => \_gnd_net_\,
            in3 => \N__55798\,
            lcout => \c0.n23313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i34_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__55800\,
            in1 => \N__75256\,
            in2 => \N__80097\,
            in3 => \N__70080\,
            lcout => \c0.data_in_frame_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1854_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54951\,
            in1 => \N__58078\,
            in2 => \_gnd_net_\,
            in3 => \N__55799\,
            lcout => \c0.n14_adj_4707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1195_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51467\,
            in1 => \N__51354\,
            in2 => \N__55905\,
            in3 => \N__51521\,
            lcout => \c0.n20_adj_4222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_2_lut_3_lut_4_lut_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60906\,
            in1 => \N__55901\,
            in2 => \N__51522\,
            in3 => \N__57731\,
            lcout => \c0.n58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1813_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58372\,
            in1 => \N__57900\,
            in2 => \N__60562\,
            in3 => \N__51345\,
            lcout => \c0.n23116\,
            ltout => \c0.n23116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1827_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51339\,
            in3 => \N__55899\,
            lcout => \c0.n11_adj_4614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i48_4_lut_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55900\,
            in1 => \N__51517\,
            in2 => \N__58173\,
            in3 => \N__66173\,
            lcout => OPEN,
            ltout => \c0.n129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i73_4_lut_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51507\,
            in1 => \N__55644\,
            in2 => \N__51492\,
            in3 => \N__58242\,
            lcout => \c0.n154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1611_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51581\,
            in1 => \N__60552\,
            in2 => \N__55682\,
            in3 => \N__62084\,
            lcout => OPEN,
            ltout => \c0.n16_adj_4613_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1612_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60905\,
            in1 => \N__51489\,
            in2 => \N__51483\,
            in3 => \N__51466\,
            lcout => \c0.n23390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56085\,
            in1 => \N__55566\,
            in2 => \N__73861\,
            in3 => \N__65835\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1585_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58544\,
            in1 => \N__58776\,
            in2 => \N__59243\,
            in3 => \N__56084\,
            lcout => \c0.n21_adj_4605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1584_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61616\,
            in1 => \N__61658\,
            in2 => \N__72693\,
            in3 => \N__58890\,
            lcout => \c0.n19_adj_4604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i116_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__76954\,
            in1 => \N__59197\,
            in2 => \N__55823\,
            in3 => \_gnd_net_\,
            lcout => data_in_frame_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i63_4_lut_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51372\,
            in1 => \N__58891\,
            in2 => \N__51675\,
            in3 => \N__66160\,
            lcout => OPEN,
            ltout => \c0.n144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i77_4_lut_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62151\,
            in1 => \N__51363\,
            in2 => \N__51357\,
            in3 => \N__51681\,
            lcout => \c0.n158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i119_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__59231\,
            in1 => \_gnd_net_\,
            in2 => \N__73356\,
            in3 => \N__59198\,
            lcout => data_in_frame_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1586_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51671\,
            in1 => \N__51657\,
            in2 => \N__51651\,
            in3 => \N__51642\,
            lcout => \c0.n21344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1196_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59300\,
            in1 => \N__51633\,
            in2 => \N__55275\,
            in3 => \N__55523\,
            lcout => OPEN,
            ltout => \c0.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51626\,
            in1 => \N__55741\,
            in2 => \N__51597\,
            in3 => \N__51594\,
            lcout => OPEN,
            ltout => \c0.n22_adj_4223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58263\,
            in1 => \N__51585\,
            in2 => \N__51531\,
            in3 => \N__60553\,
            lcout => \c0.n21_adj_4225\,
            ltout => \c0.n21_adj_4225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1257_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51528\,
            in3 => \N__77654\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1258_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56163\,
            in1 => \N__66309\,
            in2 => \N__51525\,
            in3 => \N__77583\,
            lcout => \c0.n13_adj_4281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1587_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61901\,
            in1 => \N__66570\,
            in2 => \N__63441\,
            in3 => \N__58871\,
            lcout => \c0.n10_adj_4591\,
            ltout => \c0.n10_adj_4591_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_1565_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51727\,
            in1 => \N__73854\,
            in2 => \N__51738\,
            in3 => \N__62711\,
            lcout => \c0.n41_adj_4592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1589_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__62712\,
            in1 => \N__51735\,
            in2 => \N__73862\,
            in3 => \N__65846\,
            lcout => OPEN,
            ltout => \c0.n12_adj_4606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1590_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51728\,
            in1 => \N__59479\,
            in2 => \N__51714\,
            in3 => \N__63471\,
            lcout => \c0.n21325\,
            ltout => \c0.n21325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1559_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51711\,
            in3 => \N__76832\,
            lcout => \c0.n4_adj_4464\,
            ltout => \c0.n4_adj_4464_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1460_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51708\,
            in1 => \N__56268\,
            in2 => \N__51693\,
            in3 => \N__74733\,
            lcout => \c0.n12_adj_4506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i189_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__59480\,
            in1 => \N__71913\,
            in2 => \N__80982\,
            in3 => \N__80324\,
            lcout => \c0.data_in_frame_23_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1569_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51687\,
            in1 => \N__51864\,
            in2 => \N__63089\,
            in3 => \N__59440\,
            lcout => \c0.n23863\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1570_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__65853\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63381\,
            lcout => \c0.n21428\,
            ltout => \c0.n21428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1566_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51834\,
            in1 => \N__58527\,
            in2 => \N__51690\,
            in3 => \N__56323\,
            lcout => \c0.n24_adj_4593\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__65854\,
            in1 => \N__66431\,
            in2 => \_gnd_net_\,
            in3 => \N__51843\,
            lcout => \c0.n23_adj_4598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1372_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77688\,
            in1 => \N__58482\,
            in2 => \N__51858\,
            in3 => \N__58794\,
            lcout => \c0.n23_adj_4353\,
            ltout => \c0.n23_adj_4353_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1393_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72360\,
            in1 => \N__56427\,
            in2 => \N__51837\,
            in3 => \N__51833\,
            lcout => \c0.n16_adj_4437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1394_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__58523\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56322\,
            lcout => OPEN,
            ltout => \c0.n11_adj_4438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1395_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59286\,
            in1 => \N__51825\,
            in2 => \N__51819\,
            in3 => \N__51816\,
            lcout => \c0.n21280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66987\,
            in1 => \N__57887\,
            in2 => \N__66900\,
            in3 => \N__59442\,
            lcout => \c0.n22420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1463_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67706\,
            in1 => \N__56272\,
            in2 => \N__51801\,
            in3 => \N__51903\,
            lcout => \c0.n24_adj_4509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_adj_1397_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57886\,
            in2 => \_gnd_net_\,
            in3 => \N__59441\,
            lcout => OPEN,
            ltout => \c0.n23187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1399_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51780\,
            in1 => \N__67194\,
            in2 => \N__51741\,
            in3 => \N__66986\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4439_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1402_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59738\,
            in1 => \N__66893\,
            in2 => \N__51960\,
            in3 => \N__66929\,
            lcout => OPEN,
            ltout => \c0.n13_adj_4442_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1403_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51957\,
            in1 => \N__63276\,
            in2 => \N__51951\,
            in3 => \N__61935\,
            lcout => \c0.n24528\,
            ltout => \c0.n24528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1551_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__73772\,
            in2 => \N__51948\,
            in3 => \N__51943\,
            lcout => \c0.n23533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1477_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62549\,
            in1 => \N__63792\,
            in2 => \N__52101\,
            in3 => \N__51924\,
            lcout => \c0.n10_adj_4513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1466_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63243\,
            in1 => \N__51915\,
            in2 => \N__62980\,
            in3 => \N__51909\,
            lcout => \c0.n24559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1462_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56854\,
            in1 => \N__52133\,
            in2 => \N__56574\,
            in3 => \N__67505\,
            lcout => \c0.n22_adj_4507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1481_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52132\,
            in1 => \N__51969\,
            in2 => \N__77292\,
            in3 => \N__56751\,
            lcout => \c0.n23627\,
            ltout => \c0.n23627_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1733_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52167\,
            in1 => \N__52206\,
            in2 => \N__51891\,
            in3 => \N__51881\,
            lcout => \c0.n21353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1540_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52166\,
            in2 => \_gnd_net_\,
            in3 => \N__63242\,
            lcout => \c0.n10_adj_4575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i205_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__74135\,
            in1 => \N__59868\,
            in2 => \N__71921\,
            in3 => \N__79397\,
            lcout => \c0.data_in_frame_25_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1519_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67140\,
            in2 => \_gnd_net_\,
            in3 => \N__52090\,
            lcout => \c0.n22505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i221_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__76655\,
            in1 => \N__71866\,
            in2 => \N__57081\,
            in3 => \N__79398\,
            lcout => \c0.data_in_frame_27_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i220_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__79396\,
            in1 => \N__76944\,
            in2 => \N__57112\,
            in3 => \N__76656\,
            lcout => \c0.data_in_frame_27_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_345_2_lut_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57102\,
            in2 => \_gnd_net_\,
            in3 => \N__57072\,
            lcout => \c0.n25467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1504_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67883\,
            in1 => \N__52029\,
            in2 => \N__52017\,
            in3 => \N__51999\,
            lcout => \c0.n10_adj_4544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1487_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52110\,
            in1 => \N__59867\,
            in2 => \N__51984\,
            in3 => \N__56753\,
            lcout => \c0.n10874\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_17_i3_2_lut_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__53099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__71471\,
            lcout => \c0.n3_adj_4402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_19_i3_2_lut_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__71472\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53180\,
            lcout => \c0.n3_adj_4398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_1755_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__56372\,
            in1 => \_gnd_net_\,
            in2 => \N__56407\,
            in3 => \N__63240\,
            lcout => \c0.n10_adj_4371\,
            ltout => \c0.n10_adj_4371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1391_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52134\,
            in2 => \N__52113\,
            in3 => \N__56522\,
            lcout => \c0.n12_adj_4372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_20_i3_2_lut_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53136\,
            in2 => \_gnd_net_\,
            in3 => \N__71473\,
            lcout => \c0.n3_adj_4396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1724_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56239\,
            in2 => \_gnd_net_\,
            in3 => \N__62317\,
            lcout => \c0.n12_adj_4671\,
            ltout => \c0.n12_adj_4671_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i235_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__79125\,
            in1 => \N__56705\,
            in2 => \N__52104\,
            in3 => \N__75393\,
            lcout => \c0.data_in_frame_29_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3725_2_lut_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56396\,
            in2 => \_gnd_net_\,
            in3 => \N__56371\,
            lcout => \c0.n6404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63906\,
            in1 => \N__56797\,
            in2 => \N__57001\,
            in3 => \N__74874\,
            lcout => \c0.n23_adj_4551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_21_i3_2_lut_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53220\,
            in2 => \_gnd_net_\,
            in3 => \N__71394\,
            lcout => \c0.n3_adj_4394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1503_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__63907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56798\,
            lcout => \c0.n22227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i208_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__74203\,
            in1 => \N__76354\,
            in2 => \N__63917\,
            in3 => \N__79440\,
            lcout => \c0.data_in_frame_25_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1453_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__74837\,
            in1 => \N__75969\,
            in2 => \N__52245\,
            in3 => \N__59901\,
            lcout => \c0.n22_adj_4498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i201_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__74202\,
            in1 => \N__80703\,
            in2 => \N__79477\,
            in3 => \N__56994\,
            lcout => \c0.data_in_frame_25_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i206_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__79439\,
            in1 => \N__74204\,
            in2 => \N__56816\,
            in3 => \N__79627\,
            lcout => \c0.data_in_frame_25_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1273_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52481\,
            in1 => \N__53376\,
            in2 => \N__53181\,
            in3 => \N__52694\,
            lcout => \c0.n45_adj_4298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1482_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52155\,
            in2 => \_gnd_net_\,
            in3 => \N__52191\,
            lcout => \c0.n22334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_1250_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__53341\,
            in1 => \N__53219\,
            in2 => \N__53103\,
            in3 => \N__53514\,
            lcout => \c0.n44_adj_4270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i203_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__79441\,
            in1 => \N__79172\,
            in2 => \N__52165\,
            in3 => \N__74209\,
            lcout => \c0.data_in_frame_25_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78770\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_12_i3_2_lut_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52905\,
            in2 => \_gnd_net_\,
            in3 => \N__71454\,
            lcout => \c0.n3_adj_4412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1269_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__53007\,
            in1 => \N__52721\,
            in2 => \N__53487\,
            in3 => \N__70400\,
            lcout => \c0.n40_adj_4294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_10_i3_2_lut_LC_18_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52722\,
            in2 => \_gnd_net_\,
            in3 => \N__71455\,
            lcout => \c0.n3_adj_4416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_25_i3_2_lut_LC_18_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53375\,
            in2 => \_gnd_net_\,
            in3 => \N__71456\,
            lcout => \c0.n3_adj_4386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_LC_18_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52552\,
            in1 => \N__71588\,
            in2 => \N__53313\,
            in3 => \N__53547\,
            lcout => OPEN,
            ltout => \c0.n42_adj_4272_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_1271_LC_18_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52251\,
            in1 => \N__52272\,
            in2 => \N__52266\,
            in3 => \N__52263\,
            lcout => \c0.n50_adj_4296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_LC_18_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52628\,
            in1 => \N__53132\,
            in2 => \N__52959\,
            in3 => \N__52904\,
            lcout => \c0.n43_adj_4275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_26_i3_2_lut_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__71457\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53408\,
            lcout => \c0.n3_adj_4384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_27_i3_2_lut_LC_18_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53441\,
            in2 => \_gnd_net_\,
            in3 => \N__71458\,
            lcout => \c0.n3_adj_4382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_28_i3_2_lut_LC_18_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__71504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53480\,
            lcout => \c0.n3_adj_4380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_29_i3_2_lut_LC_18_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53543\,
            in2 => \_gnd_net_\,
            in3 => \N__71505\,
            lcout => \c0.n3_adj_4378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_30_i3_2_lut_LC_18_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53510\,
            in2 => \_gnd_net_\,
            in3 => \N__71506\,
            lcout => \c0.n3_adj_4376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i0_LC_19_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74238\,
            in2 => \N__52284\,
            in3 => \N__53765\,
            lcout => \c0.FRAME_MATCHER_i_0\,
            ltout => OPEN,
            carryin => \bfn_19_1_0_\,
            carryout => \c0.n19625\,
            clk => \N__78825\,
            ce => 'H',
            sr => \N__54903\
        );

    \c0.add_49_2_THRU_CRY_0_LC_19_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54581\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19625\,
            carryout => \c0.n19625_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_1_LC_19_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54630\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19625_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19625_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_2_LC_19_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54585\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19625_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19625_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_3_LC_19_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54631\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19625_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19625_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_4_LC_19_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54589\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19625_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19625_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_5_LC_19_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54632\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19625_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19625_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_6_LC_19_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54593\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19625_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19625_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i1_LC_19_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53764\,
            in1 => \N__74406\,
            in2 => \_gnd_net_\,
            in3 => \N__52275\,
            lcout => \c0.FRAME_MATCHER_i_1\,
            ltout => OPEN,
            carryin => \bfn_19_2_0_\,
            carryout => \c0.n19626\,
            clk => \N__78823\,
            ce => 'H',
            sr => \N__52317\
        );

    \c0.add_49_3_THRU_CRY_0_LC_19_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54462\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19626\,
            carryout => \c0.n19626_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_1_LC_19_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54578\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19626_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19626_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_2_LC_19_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54466\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19626_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19626_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_3_LC_19_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54579\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19626_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19626_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_4_LC_19_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54470\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19626_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19626_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_5_LC_19_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54580\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19626_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19626_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_6_LC_19_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54474\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19626_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19626_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i2_LC_19_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53769\,
            in1 => \N__74562\,
            in2 => \_gnd_net_\,
            in3 => \N__52302\,
            lcout => \c0.FRAME_MATCHER_i_2\,
            ltout => OPEN,
            carryin => \bfn_19_3_0_\,
            carryout => \c0.n19627\,
            clk => \N__78821\,
            ce => 'H',
            sr => \N__52299\
        );

    \c0.add_49_4_THRU_CRY_0_LC_19_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54449\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19627\,
            carryout => \c0.n19627_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_1_LC_19_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54575\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19627_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19627_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_2_LC_19_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54453\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19627_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19627_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_3_LC_19_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54576\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19627_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19627_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_4_LC_19_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54457\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19627_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19627_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_5_LC_19_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54577\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19627_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19627_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_6_LC_19_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54461\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19627_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19627_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i3_LC_19_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53760\,
            in1 => \N__62197\,
            in2 => \_gnd_net_\,
            in3 => \N__52320\,
            lcout => \c0.FRAME_MATCHER_i_3\,
            ltout => OPEN,
            carryin => \bfn_19_4_0_\,
            carryout => \c0.n19628\,
            clk => \N__78817\,
            ce => 'H',
            sr => \N__62166\
        );

    \c0.add_49_5_THRU_CRY_0_LC_19_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54436\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19628\,
            carryout => \c0.n19628_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_1_LC_19_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54572\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19628_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19628_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_2_LC_19_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54440\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19628_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19628_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_3_LC_19_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54573\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19628_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19628_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_4_LC_19_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54444\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19628_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19628_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_5_LC_19_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54574\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19628_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19628_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_6_LC_19_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54448\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19628_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19628_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i4_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53759\,
            in1 => \N__52362\,
            in2 => \_gnd_net_\,
            in3 => \N__52335\,
            lcout => \c0.FRAME_MATCHER_i_4\,
            ltout => OPEN,
            carryin => \bfn_19_5_0_\,
            carryout => \c0.n19629\,
            clk => \N__78813\,
            ce => 'H',
            sr => \N__52332\
        );

    \c0.add_49_6_THRU_CRY_0_LC_19_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54423\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19629\,
            carryout => \c0.n19629_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_1_LC_19_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54569\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19629_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19629_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_2_LC_19_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54427\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19629_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19629_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_3_LC_19_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54570\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19629_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19629_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_4_LC_19_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54431\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19629_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19629_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_5_LC_19_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54571\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19629_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19629_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_6_LC_19_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54435\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19629_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19629_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i5_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53748\,
            in1 => \N__52454\,
            in2 => \_gnd_net_\,
            in3 => \N__52425\,
            lcout => \c0.FRAME_MATCHER_i_5\,
            ltout => OPEN,
            carryin => \bfn_19_6_0_\,
            carryout => \c0.n19630\,
            clk => \N__78804\,
            ce => 'H',
            sr => \N__52422\
        );

    \c0.add_49_7_THRU_CRY_0_LC_19_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54231\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19630\,
            carryout => \c0.n19630_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_1_LC_19_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54420\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19630_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19630_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_2_LC_19_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54235\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19630_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19630_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_3_LC_19_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54421\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19630_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19630_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_4_LC_19_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54239\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19630_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19630_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_5_LC_19_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54422\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19630_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19630_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_6_LC_19_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54243\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19630_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19630_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i6_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53747\,
            in1 => \N__52525\,
            in2 => \_gnd_net_\,
            in3 => \N__52509\,
            lcout => \c0.FRAME_MATCHER_i_6\,
            ltout => OPEN,
            carryin => \bfn_19_7_0_\,
            carryout => \c0.n19631\,
            clk => \N__78795\,
            ce => 'H',
            sr => \N__52506\
        );

    \c0.add_49_8_THRU_CRY_0_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54218\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19631\,
            carryout => \c0.n19631_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_1_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54417\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19631_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19631_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_2_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54222\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19631_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19631_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_3_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54418\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19631_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19631_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_4_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54226\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19631_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19631_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_5_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54419\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19631_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19631_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_6_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54230\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19631_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19631_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i7_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53746\,
            in1 => \N__52615\,
            in2 => \_gnd_net_\,
            in3 => \N__52599\,
            lcout => \c0.FRAME_MATCHER_i_7\,
            ltout => OPEN,
            carryin => \bfn_19_8_0_\,
            carryout => \c0.n19632\,
            clk => \N__78788\,
            ce => 'H',
            sr => \N__52596\
        );

    \c0.add_49_9_THRU_CRY_0_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54138\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19632\,
            carryout => \c0.n19632_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_1_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54314\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19632_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19632_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_2_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54142\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19632_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19632_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_3_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54315\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19632_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19632_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_4_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54146\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19632_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19632_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_5_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54316\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19632_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19632_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_6_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54150\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19632_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19632_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i8_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53745\,
            in1 => \N__52669\,
            in2 => \_gnd_net_\,
            in3 => \N__52653\,
            lcout => \c0.FRAME_MATCHER_i_8\,
            ltout => OPEN,
            carryin => \bfn_19_9_0_\,
            carryout => \c0.n19633\,
            clk => \N__78782\,
            ce => 'H',
            sr => \N__52650\
        );

    \c0.add_49_10_THRU_CRY_0_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53995\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19633\,
            carryout => \c0.n19633_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_1_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53999\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19633_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19633_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_2_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53996\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19633_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19633_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_3_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54000\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19633_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19633_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_4_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53997\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19633_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19633_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_5_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54001\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19633_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19633_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_6_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53998\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19633_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19633_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i9_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53744\,
            in1 => \N__52756\,
            in2 => \_gnd_net_\,
            in3 => \N__52740\,
            lcout => \c0.FRAME_MATCHER_i_9\,
            ltout => OPEN,
            carryin => \bfn_19_10_0_\,
            carryout => \c0.n19634\,
            clk => \N__78772\,
            ce => 'H',
            sr => \N__52737\
        );

    \c0.add_49_11_THRU_CRY_0_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54307\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19634\,
            carryout => \c0.n19634_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_1_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54311\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19634_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19634_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_2_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54308\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19634_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19634_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_3_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54312\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19634_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19634_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_4_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54309\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19634_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19634_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_5_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54313\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19634_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19634_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_6_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54310\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19634_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19634_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i10_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53743\,
            in1 => \N__52712\,
            in2 => \_gnd_net_\,
            in3 => \N__52698\,
            lcout => \c0.FRAME_MATCHER_i_10\,
            ltout => OPEN,
            carryin => \bfn_19_11_0_\,
            carryout => \c0.n19635\,
            clk => \N__78761\,
            ce => 'H',
            sr => \N__52854\
        );

    \c0.add_49_12_THRU_CRY_0_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54317\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19635\,
            carryout => \c0.n19635_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_1_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54321\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19635_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19635_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_2_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54318\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19635_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19635_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_3_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54322\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19635_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19635_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_4_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54319\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19635_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19635_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_5_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54323\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19635_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19635_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_6_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54320\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19635_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19635_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i11_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53742\,
            in1 => \N__52816\,
            in2 => \_gnd_net_\,
            in3 => \N__52800\,
            lcout => \c0.FRAME_MATCHER_i_11\,
            ltout => OPEN,
            carryin => \bfn_19_12_0_\,
            carryout => \c0.n19636\,
            clk => \N__78749\,
            ce => 'H',
            sr => \N__52797\
        );

    \c0.add_49_13_THRU_CRY_0_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54324\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19636\,
            carryout => \c0.n19636_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_1_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54328\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19636_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19636_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_2_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54325\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19636_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19636_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_3_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54329\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19636_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19636_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_4_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54326\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19636_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19636_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_5_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54330\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19636_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19636_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_6_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54327\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19636_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19636_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i12_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53741\,
            in1 => \N__52891\,
            in2 => \_gnd_net_\,
            in3 => \N__52875\,
            lcout => \c0.FRAME_MATCHER_i_12\,
            ltout => OPEN,
            carryin => \bfn_19_13_0_\,
            carryout => \c0.n19637\,
            clk => \N__78736\,
            ce => 'H',
            sr => \N__52872\
        );

    \c0.add_49_14_THRU_CRY_0_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54331\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19637\,
            carryout => \c0.n19637_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_1_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54335\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19637_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19637_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_2_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54332\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19637_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19637_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_3_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54336\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19637_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19637_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_4_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54333\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19637_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19637_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_5_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54337\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19637_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19637_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_6_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54334\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19637_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19637_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i13_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53740\,
            in1 => \N__70387\,
            in2 => \_gnd_net_\,
            in3 => \N__52908\,
            lcout => \c0.FRAME_MATCHER_i_13\,
            ltout => OPEN,
            carryin => \bfn_19_14_0_\,
            carryout => \c0.n19638\,
            clk => \N__78723\,
            ce => 'H',
            sr => \N__70368\
        );

    \c0.add_49_15_THRU_CRY_0_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54490\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19638\,
            carryout => \c0.n19638_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_1_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54494\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19638_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19638_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_2_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54491\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19638_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19638_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_3_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54495\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19638_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19638_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_4_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54492\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19638_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19638_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_5_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54496\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19638_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19638_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_6_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54493\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19638_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19638_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i14_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53768\,
            in1 => \N__52942\,
            in2 => \_gnd_net_\,
            in3 => \N__52923\,
            lcout => \c0.FRAME_MATCHER_i_14\,
            ltout => OPEN,
            carryin => \bfn_19_15_0_\,
            carryout => \c0.n19639\,
            clk => \N__78713\,
            ce => 'H',
            sr => \N__52920\
        );

    \c0.add_49_16_THRU_CRY_0_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54497\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19639\,
            carryout => \c0.n19639_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_1_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54501\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19639_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19639_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_2_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54498\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19639_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19639_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_3_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54502\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19639_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19639_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_4_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54499\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19639_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19639_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_5_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54503\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19639_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19639_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_6_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54500\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19639_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19639_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i15_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53767\,
            in1 => \N__52996\,
            in2 => \_gnd_net_\,
            in3 => \N__52977\,
            lcout => \c0.FRAME_MATCHER_i_15\,
            ltout => OPEN,
            carryin => \bfn_19_16_0_\,
            carryout => \c0.n19640\,
            clk => \N__78698\,
            ce => 'H',
            sr => \N__52974\
        );

    \c0.add_49_17_THRU_CRY_0_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54504\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19640\,
            carryout => \c0.n19640_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_1_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54508\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19640_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19640_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_2_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54505\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19640_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19640_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_3_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54509\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19640_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19640_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_4_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54506\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19640_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19640_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_5_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54510\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19640_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19640_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_6_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54507\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19640_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19640_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i16_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53766\,
            in1 => \N__53038\,
            in2 => \_gnd_net_\,
            in3 => \N__53022\,
            lcout => \c0.FRAME_MATCHER_i_16\,
            ltout => OPEN,
            carryin => \bfn_19_17_0_\,
            carryout => \c0.n19641\,
            clk => \N__78670\,
            ce => 'H',
            sr => \N__53019\
        );

    \c0.add_49_18_THRU_CRY_0_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54511\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19641\,
            carryout => \c0.n19641_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_1_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54515\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19641_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19641_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_2_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54512\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19641_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19641_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_3_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54516\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19641_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19641_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_4_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54513\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19641_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19641_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_5_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54517\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19641_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19641_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_6_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54514\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19641_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19641_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i17_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53724\,
            in1 => \N__53089\,
            in2 => \_gnd_net_\,
            in3 => \N__53073\,
            lcout => \c0.FRAME_MATCHER_i_17\,
            ltout => OPEN,
            carryin => \bfn_19_18_0_\,
            carryout => \c0.n19642\,
            clk => \N__78699\,
            ce => 'H',
            sr => \N__53070\
        );

    \c0.add_49_19_THRU_CRY_0_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54020\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19642\,
            carryout => \c0.n19642_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_1_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54024\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19642_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19642_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_2_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54021\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19642_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19642_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_3_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54025\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19642_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19642_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_4_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54022\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19642_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19642_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_5_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54026\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19642_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19642_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_6_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54023\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19642_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19642_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i18_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53749\,
            in1 => \N__71572\,
            in2 => \_gnd_net_\,
            in3 => \N__53106\,
            lcout => \c0.FRAME_MATCHER_i_18\,
            ltout => OPEN,
            carryin => \bfn_19_19_0_\,
            carryout => \c0.n19643\,
            clk => \N__78714\,
            ce => 'H',
            sr => \N__71295\
        );

    \c0.add_49_20_THRU_CRY_0_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54594\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19643\,
            carryout => \c0.n19643_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_1_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54598\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19643_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19643_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_2_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54595\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19643_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19643_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_3_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54599\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19643_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19643_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_4_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54596\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19643_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19643_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_5_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54600\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19643_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19643_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_6_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54597\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19643_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19643_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i19_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53713\,
            in1 => \N__53170\,
            in2 => \_gnd_net_\,
            in3 => \N__53154\,
            lcout => \c0.FRAME_MATCHER_i_19\,
            ltout => OPEN,
            carryin => \bfn_19_20_0_\,
            carryout => \c0.n19644\,
            clk => \N__78724\,
            ce => 'H',
            sr => \N__53151\
        );

    \c0.add_49_21_THRU_CRY_0_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54601\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19644\,
            carryout => \c0.n19644_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_1_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54605\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19644_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19644_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_2_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54602\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19644_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19644_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_3_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54606\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19644_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19644_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_4_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54603\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19644_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19644_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_5_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54607\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19644_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19644_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_6_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54604\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19644_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19644_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i20_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53712\,
            in1 => \N__53125\,
            in2 => \_gnd_net_\,
            in3 => \N__53109\,
            lcout => \c0.FRAME_MATCHER_i_20\,
            ltout => OPEN,
            carryin => \bfn_19_21_0_\,
            carryout => \c0.n19645\,
            clk => \N__78737\,
            ce => 'H',
            sr => \N__53232\
        );

    \c0.add_49_22_THRU_CRY_0_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54608\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19645\,
            carryout => \c0.n19645_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_1_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54612\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19645_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19645_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_2_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54609\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19645_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19645_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_3_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54613\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19645_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19645_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_4_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54610\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19645_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19645_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_5_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54614\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19645_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19645_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_6_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54611\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19645_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19645_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i21_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53698\,
            in1 => \N__53212\,
            in2 => \_gnd_net_\,
            in3 => \N__53196\,
            lcout => \c0.FRAME_MATCHER_i_21\,
            ltout => OPEN,
            carryin => \bfn_19_22_0_\,
            carryout => \c0.n19646\,
            clk => \N__78750\,
            ce => 'H',
            sr => \N__53193\
        );

    \c0.add_49_23_THRU_CRY_0_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54714\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19646\,
            carryout => \c0.n19646_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_1_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54718\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19646_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19646_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_2_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54715\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19646_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19646_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_3_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54719\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19646_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19646_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_4_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54716\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19646_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19646_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_5_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54720\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19646_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19646_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_6_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54717\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19646_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19646_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i22_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53697\,
            in1 => \N__53263\,
            in2 => \_gnd_net_\,
            in3 => \N__53247\,
            lcout => \c0.FRAME_MATCHER_i_22\,
            ltout => OPEN,
            carryin => \bfn_19_23_0_\,
            carryout => \c0.n19647\,
            clk => \N__78762\,
            ce => 'H',
            sr => \N__53244\
        );

    \c0.add_49_24_THRU_CRY_0_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54827\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19647\,
            carryout => \c0.n19647_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_1_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54724\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19647_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19647_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_2_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54828\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19647_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19647_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_3_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54728\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19647_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19647_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_4_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54829\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19647_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19647_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_5_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54732\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19647_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19647_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_6_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54830\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19647_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19647_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i23_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53696\,
            in1 => \N__53302\,
            in2 => \_gnd_net_\,
            in3 => \N__53283\,
            lcout => \c0.FRAME_MATCHER_i_23\,
            ltout => OPEN,
            carryin => \bfn_19_24_0_\,
            carryout => \c0.n19648\,
            clk => \N__78773\,
            ce => 'H',
            sr => \N__53280\
        );

    \c0.add_49_25_THRU_CRY_0_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54736\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19648\,
            carryout => \c0.n19648_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_1_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54740\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19648_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19648_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_2_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54737\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19648_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19648_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_3_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54741\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19648_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19648_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_4_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54738\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19648_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19648_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_5_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54742\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19648_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19648_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_6_LC_19_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54739\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19648_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19648_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i24_LC_19_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53695\,
            in1 => \N__53342\,
            in2 => \_gnd_net_\,
            in3 => \N__53325\,
            lcout => \c0.FRAME_MATCHER_i_24\,
            ltout => OPEN,
            carryin => \bfn_19_25_0_\,
            carryout => \c0.n19649\,
            clk => \N__78781\,
            ce => 'H',
            sr => \N__53322\
        );

    \c0.add_49_26_THRU_CRY_0_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54831\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19649\,
            carryout => \c0.n19649_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_1_LC_19_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54746\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19649_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19649_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_2_LC_19_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54832\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19649_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19649_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_3_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54750\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19649_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19649_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_4_LC_19_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54833\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19649_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19649_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_5_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54754\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19649_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19649_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_6_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__54834\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19649_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19649_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i25_LC_19_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53694\,
            in1 => \N__53374\,
            in2 => \_gnd_net_\,
            in3 => \N__53355\,
            lcout => \c0.FRAME_MATCHER_i_25\,
            ltout => OPEN,
            carryin => \bfn_19_26_0_\,
            carryout => \c0.n19650\,
            clk => \N__78787\,
            ce => 'H',
            sr => \N__53352\
        );

    \c0.add_49_27_THRU_CRY_0_LC_19_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54835\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19650\,
            carryout => \c0.n19650_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_1_LC_19_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54839\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19650_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19650_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_2_LC_19_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54836\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19650_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19650_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_3_LC_19_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54840\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19650_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19650_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_4_LC_19_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54837\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19650_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19650_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_5_LC_19_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54841\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19650_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19650_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_6_LC_19_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54838\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19650_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19650_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i26_LC_19_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53693\,
            in1 => \N__53404\,
            in2 => \_gnd_net_\,
            in3 => \N__53385\,
            lcout => \c0.FRAME_MATCHER_i_26\,
            ltout => OPEN,
            carryin => \bfn_19_27_0_\,
            carryout => \c0.n19651\,
            clk => \N__78794\,
            ce => 'H',
            sr => \N__53382\
        );

    \c0.add_49_28_THRU_CRY_0_LC_19_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54842\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19651\,
            carryout => \c0.n19651_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_1_LC_19_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54846\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19651_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19651_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_2_LC_19_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54843\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19651_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19651_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_3_LC_19_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54847\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19651_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19651_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_4_LC_19_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54844\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19651_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19651_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_5_LC_19_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54848\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19651_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19651_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_6_LC_19_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54845\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19651_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19651_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i27_LC_19_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53692\,
            in1 => \N__53440\,
            in2 => \_gnd_net_\,
            in3 => \N__53421\,
            lcout => \c0.FRAME_MATCHER_i_27\,
            ltout => OPEN,
            carryin => \bfn_19_28_0_\,
            carryout => \c0.n19652\,
            clk => \N__78803\,
            ce => 'H',
            sr => \N__53418\
        );

    \c0.add_49_29_THRU_CRY_0_LC_19_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54849\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19652\,
            carryout => \c0.n19652_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_1_LC_19_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54853\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19652_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19652_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_2_LC_19_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54850\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19652_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19652_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_3_LC_19_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54854\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19652_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19652_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_4_LC_19_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54851\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19652_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19652_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_5_LC_19_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54855\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19652_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19652_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_6_LC_19_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54852\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19652_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19652_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i28_LC_19_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53699\,
            in1 => \N__53479\,
            in2 => \_gnd_net_\,
            in3 => \N__53460\,
            lcout => \c0.FRAME_MATCHER_i_28\,
            ltout => OPEN,
            carryin => \bfn_19_29_0_\,
            carryout => \c0.n19653\,
            clk => \N__78812\,
            ce => 'H',
            sr => \N__53457\
        );

    \c0.add_49_30_THRU_CRY_0_LC_19_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54856\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19653\,
            carryout => \c0.n19653_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_1_LC_19_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54860\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19653_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19653_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_2_LC_19_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54857\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19653_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19653_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_3_LC_19_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54861\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19653_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19653_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_4_LC_19_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54858\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19653_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19653_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_5_LC_19_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54862\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19653_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19653_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_6_LC_19_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54859\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19653_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19653_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i29_LC_19_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53665\,
            in1 => \N__53542\,
            in2 => \_gnd_net_\,
            in3 => \N__53523\,
            lcout => \c0.FRAME_MATCHER_i_29\,
            ltout => OPEN,
            carryin => \bfn_19_30_0_\,
            carryout => \c0.n19654\,
            clk => \N__78816\,
            ce => 'H',
            sr => \N__53520\
        );

    \c0.add_49_31_THRU_CRY_0_LC_19_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54131\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19654\,
            carryout => \c0.n19654_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_1_LC_19_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54135\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19654_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19654_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_2_LC_19_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54132\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19654_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19654_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_3_LC_19_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54136\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19654_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19654_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_4_LC_19_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54133\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19654_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19654_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_5_LC_19_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54137\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19654_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19654_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_6_LC_19_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54134\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19654_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19654_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i30_LC_19_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53640\,
            in1 => \N__53509\,
            in2 => \_gnd_net_\,
            in3 => \N__53490\,
            lcout => \c0.FRAME_MATCHER_i_30\,
            ltout => OPEN,
            carryin => \bfn_19_31_0_\,
            carryout => \c0.n19655\,
            clk => \N__78820\,
            ce => 'H',
            sr => \N__54894\
        );

    \c0.add_49_32_THRU_CRY_0_LC_19_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54879\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19655\,
            carryout => \c0.n19655_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_1_LC_19_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54883\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19655_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19655_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_2_LC_19_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54880\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19655_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19655_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_3_LC_19_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54884\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19655_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19655_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_4_LC_19_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54881\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19655_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19655_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_5_LC_19_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54885\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19655_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19655_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_6_LC_19_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54882\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19655_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19655_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i31_LC_19_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__53641\,
            in1 => \N__53877\,
            in2 => \_gnd_net_\,
            in3 => \N__53919\,
            lcout => \c0.FRAME_MATCHER_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78824\,
            ce => 'H',
            sr => \N__53823\
        );

    \c0.i14251_1_lut_LC_19_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53814\,
            lcout => \c0.n1306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_0_i3_2_lut_LC_20_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74302\,
            in2 => \_gnd_net_\,
            in3 => \N__71552\,
            lcout => \c0.n3_adj_4436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1610_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60131\,
            in1 => \N__60686\,
            in2 => \N__58403\,
            in3 => \N__60116\,
            lcout => \c0.n23677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i81_LC_20_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__73709\,
            in1 => \N__69183\,
            in2 => \N__80736\,
            in3 => \N__58399\,
            lcout => \c0.data_in_frame_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i41_4_lut_LC_20_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55100\,
            in1 => \N__58395\,
            in2 => \N__69362\,
            in3 => \N__64529\,
            lcout => \c0.n97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i75_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__64530\,
            in1 => \N__79108\,
            in2 => \N__73719\,
            in3 => \N__74115\,
            lcout => \c0.data_in_frame_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i74_LC_20_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__75249\,
            in1 => \N__74111\,
            in2 => \N__69363\,
            in3 => \N__73715\,
            lcout => \c0.data_in_frame_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13936_4_lut_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__57030\,
            in1 => \N__68757\,
            in2 => \N__60312\,
            in3 => \N__59931\,
            lcout => \c0.n17537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i66_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__75248\,
            in1 => \N__72880\,
            in2 => \N__55113\,
            in3 => \N__73714\,
            lcout => \c0.data_in_frame_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i83_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__73710\,
            in1 => \N__69184\,
            in2 => \N__55045\,
            in3 => \N__79109\,
            lcout => \c0.data_in_frame_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1613_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57322\,
            in1 => \N__54909\,
            in2 => \N__55329\,
            in3 => \N__60295\,
            lcout => \c0.n10_adj_4615\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1836_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60631\,
            in1 => \N__54968\,
            in2 => \_gnd_net_\,
            in3 => \N__61036\,
            lcout => \c0.n22196\,
            ltout => \c0.n22196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57323\,
            in1 => \N__60296\,
            in2 => \N__54987\,
            in3 => \N__60741\,
            lcout => \c0.n12_adj_4299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1878_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__64581\,
            in1 => \N__70348\,
            in2 => \_gnd_net_\,
            in3 => \N__57399\,
            lcout => \c0.n10_adj_4283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1648_LC_20_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57355\,
            in2 => \_gnd_net_\,
            in3 => \N__55206\,
            lcout => \c0.n11_adj_4280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i8_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__70155\,
            in1 => \N__72862\,
            in2 => \N__60243\,
            in3 => \N__76316\,
            lcout => \c0.data_in_frame_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1874_LC_20_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57365\,
            in1 => \N__55207\,
            in2 => \N__57409\,
            in3 => \N__64768\,
            lcout => \c0.n12_adj_4258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i25_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__70154\,
            in1 => \N__54969\,
            in2 => \N__76630\,
            in3 => \N__80711\,
            lcout => \c0.data_in_frame_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1620_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68510\,
            in2 => \N__54960\,
            in3 => \N__60742\,
            lcout => \c0.n13523\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1549_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__54943\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60186\,
            lcout => \c0.n7_adj_4300\,
            ltout => \c0.n7_adj_4300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1278_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70742\,
            in1 => \N__55251\,
            in2 => \N__55245\,
            in3 => \N__68511\,
            lcout => \c0.n22316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1694_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55134\,
            in1 => \N__55188\,
            in2 => \N__55241\,
            in3 => \N__64773\,
            lcout => \c0.n23655\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1643_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60187\,
            in1 => \N__60635\,
            in2 => \_gnd_net_\,
            in3 => \N__60297\,
            lcout => \c0.n23251\,
            ltout => \c0.n23251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_4_lut_adj_1664_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57377\,
            in1 => \N__55187\,
            in2 => \N__55152\,
            in3 => \N__64772\,
            lcout => \c0.n7_adj_4282\,
            ltout => \c0.n7_adj_4282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1260_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55630\,
            in1 => \N__55149\,
            in2 => \N__55137\,
            in3 => \N__55133\,
            lcout => \c0.n22472\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1686_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55338\,
            in1 => \N__60235\,
            in2 => \N__57263\,
            in3 => \N__57298\,
            lcout => OPEN,
            ltout => \c0.n13_adj_4638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1639_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55049\,
            in1 => \N__55114\,
            in2 => \N__55080\,
            in3 => \N__57435\,
            lcout => \c0.n13_adj_4610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_2_lut_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57297\,
            in2 => \_gnd_net_\,
            in3 => \N__60234\,
            lcout => \c0.n68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i42_4_lut_adj_1409_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57416\,
            in1 => \N__55077\,
            in2 => \N__55050\,
            in3 => \N__55022\,
            lcout => \c0.n98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1249_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57958\,
            in1 => \N__55362\,
            in2 => \N__55564\,
            in3 => \N__55350\,
            lcout => \c0.n4_adj_4269\,
            ltout => \c0.n4_adj_4269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i33_4_lut_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55330\,
            in1 => \N__61859\,
            in2 => \N__55290\,
            in3 => \N__60148\,
            lcout => OPEN,
            ltout => \c0.n89_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i45_4_lut_adj_1408_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55287\,
            in1 => \N__60547\,
            in2 => \N__55281\,
            in3 => \N__71093\,
            lcout => \c0.n101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1619_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71092\,
            in1 => \N__57186\,
            in2 => \N__69252\,
            in3 => \N__70602\,
            lcout => \c0.n22_adj_4622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58548\,
            in1 => \N__57662\,
            in2 => \N__59265\,
            in3 => \N__60818\,
            lcout => OPEN,
            ltout => \c0.n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58281\,
            in1 => \N__55478\,
            in2 => \N__55278\,
            in3 => \N__55767\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_1787_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60817\,
            in2 => \_gnd_net_\,
            in3 => \N__58280\,
            lcout => \c0.n13075\,
            ltout => \c0.n13075_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i37_4_lut_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60792\,
            in1 => \N__68970\,
            in2 => \N__55257\,
            in3 => \N__61294\,
            lcout => OPEN,
            ltout => \c0.n93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i47_4_lut_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55766\,
            in1 => \N__60924\,
            in2 => \N__55254\,
            in3 => \N__68750\,
            lcout => \c0.n103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_3_lut_4_lut_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71091\,
            in1 => \N__58054\,
            in2 => \N__57783\,
            in3 => \N__60080\,
            lcout => \c0.n23156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i66_4_lut_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62123\,
            in1 => \N__55434\,
            in2 => \N__55392\,
            in3 => \N__55410\,
            lcout => OPEN,
            ltout => \c0.n147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i74_4_lut_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61094\,
            in1 => \N__70229\,
            in2 => \N__55401\,
            in3 => \N__55398\,
            lcout => \c0.n155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i53_4_lut_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57684\,
            in1 => \N__55632\,
            in2 => \N__57672\,
            in3 => \N__56005\,
            lcout => \c0.n134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i50_4_lut_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70445\,
            in1 => \N__65576\,
            in2 => \N__71280\,
            in3 => \N__62858\,
            lcout => \c0.n131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1262_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69837\,
            in1 => \N__70444\,
            in2 => \N__62859\,
            in3 => \N__55839\,
            lcout => \c0.n31_adj_4284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_3_lut_4_lut_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57667\,
            in1 => \N__57683\,
            in2 => \N__56009\,
            in3 => \N__60957\,
            lcout => \c0.n38_adj_4448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1411_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__64986\,
            in1 => \N__70443\,
            in2 => \N__70787\,
            in3 => \N__57822\,
            lcout => \c0.n36_adj_4447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_1414_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57732\,
            in1 => \N__58162\,
            in2 => \N__58458\,
            in3 => \N__55368\,
            lcout => OPEN,
            ltout => \c0.n41_adj_4452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_adj_1416_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55587\,
            in1 => \N__55593\,
            in2 => \N__55635\,
            in3 => \N__57966\,
            lcout => \c0.n24540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1415_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60416\,
            in1 => \N__55631\,
            in2 => \N__70677\,
            in3 => \N__59366\,
            lcout => \c0.n39_adj_4453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1413_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58051\,
            in1 => \N__70854\,
            in2 => \N__64059\,
            in3 => \N__57801\,
            lcout => \c0.n40_adj_4451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_4_lut_adj_1606_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71114\,
            in1 => \N__69585\,
            in2 => \N__60427\,
            in3 => \N__58053\,
            lcout => \c0.n22_adj_4244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1673_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58049\,
            in1 => \N__60414\,
            in2 => \_gnd_net_\,
            in3 => \N__71113\,
            lcout => \c0.n23178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_adj_1828_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__60415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58050\,
            lcout => \c0.n31_adj_4701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_3_lut_4_lut_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58052\,
            in1 => \N__60417\,
            in2 => \N__65040\,
            in3 => \N__71115\,
            lcout => \c0.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1847_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61334\,
            in1 => \N__55760\,
            in2 => \N__55581\,
            in3 => \N__55565\,
            lcout => \c0.n13721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1599_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55533\,
            in1 => \N__55524\,
            in2 => \N__55482\,
            in3 => \N__55454\,
            lcout => \c0.n23611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i85_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__71936\,
            in1 => \N__69195\,
            in2 => \N__55779\,
            in3 => \N__73610\,
            lcout => \c0.data_in_frame_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1741_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55797\,
            in2 => \_gnd_net_\,
            in3 => \N__60413\,
            lcout => \c0.n8_adj_4673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i68_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__72898\,
            in1 => \N__73608\,
            in2 => \N__72309\,
            in3 => \N__77123\,
            lcout => \c0.data_in_frame_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i84_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__69194\,
            in1 => \N__77122\,
            in2 => \N__73684\,
            in3 => \N__55972\,
            lcout => \c0.data_in_frame_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i69_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__71937\,
            in1 => \N__73609\,
            in2 => \N__76047\,
            in3 => \N__72899\,
            lcout => \c0.data_in_frame_8_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__72283\,
            in1 => \N__55775\,
            in2 => \_gnd_net_\,
            in3 => \N__55882\,
            lcout => \c0.n22455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_4_lut_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55740\,
            in1 => \N__55686\,
            in2 => \N__74964\,
            in3 => \N__55653\,
            lcout => \c0.n65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i77_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__71875\,
            in1 => \N__61245\,
            in2 => \N__73685\,
            in3 => \N__74180\,
            lcout => \c0.data_in_frame_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i46_4_lut_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77446\,
            in1 => \N__55931\,
            in2 => \N__72006\,
            in3 => \N__55944\,
            lcout => \c0.n127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1805_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58136\,
            in2 => \_gnd_net_\,
            in3 => \N__58097\,
            lcout => \c0.n5_adj_4311\,
            ltout => \c0.n5_adj_4311_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_4_lut_adj_1357_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70885\,
            in1 => \N__61235\,
            in2 => \N__55983\,
            in3 => \N__55965\,
            lcout => \c0.n85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1785_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55943\,
            in1 => \N__65010\,
            in2 => \N__55932\,
            in3 => \N__58767\,
            lcout => \c0.n22644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i67_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__72935\,
            in1 => \N__73611\,
            in2 => \N__55898\,
            in3 => \N__79110\,
            lcout => \c0.data_in_frame_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i39_2_lut_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__62528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62666\,
            lcout => OPEN,
            ltout => \c0.n120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i71_4_lut_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61890\,
            in1 => \N__62638\,
            in2 => \N__55866\,
            in3 => \N__55863\,
            lcout => OPEN,
            ltout => \c0.n152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i79_4_lut_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69760\,
            in1 => \N__58554\,
            in2 => \N__55851\,
            in3 => \N__55848\,
            lcout => \c0.n160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_4_lut_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64340\,
            in1 => \N__70297\,
            in2 => \N__70449\,
            in3 => \N__55838\,
            lcout => OPEN,
            ltout => \c0.n30_adj_4571_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_1573_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58966\,
            in1 => \N__55824\,
            in2 => \N__55803\,
            in3 => \N__69804\,
            lcout => OPEN,
            ltout => \c0.n34_adj_4600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_1574_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56112\,
            in1 => \N__69759\,
            in2 => \N__56103\,
            in3 => \N__56100\,
            lcout => \c0.n24333\,
            ltout => \c0.n24333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1698_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__62527\,
            in1 => \_gnd_net_\,
            in2 => \N__56088\,
            in3 => \N__62476\,
            lcout => \c0.n23661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1396_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56038\,
            in1 => \N__72001\,
            in2 => \N__56073\,
            in3 => \N__65927\,
            lcout => \c0.n22173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i132_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__72965\,
            in1 => \N__80262\,
            in2 => \N__77098\,
            in3 => \N__56039\,
            lcout => \c0.data_in_frame_16_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i139_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__80259\,
            in1 => \N__74146\,
            in2 => \N__79182\,
            in3 => \N__58669\,
            lcout => \c0.data_in_frame_17_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i131_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__72964\,
            in1 => \N__80261\,
            in2 => \N__65960\,
            in3 => \N__79140\,
            lcout => \c0.data_in_frame_16_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i158_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__80260\,
            in1 => \N__76611\,
            in2 => \N__71635\,
            in3 => \N__79784\,
            lcout => \c0.data_in_frame_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i156_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__76610\,
            in1 => \N__80263\,
            in2 => \N__77099\,
            in3 => \N__59129\,
            lcout => \c0.data_in_frame_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1588_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__72002\,
            in1 => \N__62667\,
            in2 => \_gnd_net_\,
            in3 => \N__60048\,
            lcout => \c0.n22540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i80_4_lut_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56022\,
            in1 => \N__58560\,
            in2 => \N__61212\,
            in3 => \N__56247\,
            lcout => \c0.n24520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1866_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__56240\,
            in1 => \N__61429\,
            in2 => \_gnd_net_\,
            in3 => \N__62294\,
            lcout => \c0.n22104\,
            ltout => \c0.n22104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i141_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__74207\,
            in1 => \N__71958\,
            in2 => \N__56196\,
            in3 => \N__72238\,
            lcout => \c0.data_in_frame_17_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i140_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__77100\,
            in1 => \N__74208\,
            in2 => \N__58829\,
            in3 => \N__80264\,
            lcout => \c0.data_in_frame_17_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1176_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72237\,
            in2 => \_gnd_net_\,
            in3 => \N__58821\,
            lcout => \c0.n22822\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1708_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__77639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__77579\,
            lcout => OPEN,
            ltout => \c0.n22347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1311_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56192\,
            in1 => \N__59125\,
            in2 => \N__56166\,
            in3 => \N__56159\,
            lcout => \c0.n10_adj_4315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_3_lut_adj_2043_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56147\,
            in1 => \N__59730\,
            in2 => \_gnd_net_\,
            in3 => \N__75784\,
            lcout => \c0.n39_adj_4341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1204_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63141\,
            in2 => \_gnd_net_\,
            in3 => \N__72299\,
            lcout => \c0.n10_adj_4230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_3_lut_4_lut_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67376\,
            in1 => \N__67362\,
            in2 => \N__67415\,
            in3 => \N__59433\,
            lcout => \c0.n45_adj_4476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__59280\,
            in1 => \N__58715\,
            in2 => \_gnd_net_\,
            in3 => \N__58843\,
            lcout => \c0.n14_adj_4356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_4_lut_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59333\,
            in1 => \N__62682\,
            in2 => \N__58848\,
            in3 => \N__60062\,
            lcout => \c0.n22_adj_4350\,
            ltout => \c0.n22_adj_4350_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_3_lut_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__59281\,
            in1 => \_gnd_net_\,
            in2 => \N__56418\,
            in3 => \N__56324\,
            lcout => \c0.n59_adj_4351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_2_lut_adj_1991_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__58847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59282\,
            lcout => \c0.n11_adj_4505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_3_lut_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56415\,
            in1 => \N__56373\,
            in2 => \_gnd_net_\,
            in3 => \N__56325\,
            lcout => \c0.n28_adj_4504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i104_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__73598\,
            in1 => \N__80044\,
            in2 => \N__76275\,
            in3 => \N__63148\,
            lcout => \c0.data_in_frame_12_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_adj_1951_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59348\,
            in1 => \N__58500\,
            in2 => \N__58671\,
            in3 => \N__81058\,
            lcout => \c0.n20_adj_4596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1473_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__75795\,
            in1 => \N__56610\,
            in2 => \N__56298\,
            in3 => \N__56280\,
            lcout => \c0.n23975\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1994_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__74679\,
            in1 => \N__74529\,
            in2 => \N__74387\,
            in3 => \N__73597\,
            lcout => n22118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1746_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56573\,
            in1 => \N__56595\,
            in2 => \N__70818\,
            in3 => \N__66709\,
            lcout => \c0.n9_adj_4521\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1568_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56493\,
            in1 => \N__56604\,
            in2 => \N__81114\,
            in3 => \N__59031\,
            lcout => \c0.n23733\,
            ltout => \c0.n23733_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1591_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__56598\,
            in3 => \N__56594\,
            lcout => \c0.n20314\,
            ltout => \c0.n20314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1512_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56894\,
            in1 => \N__56572\,
            in2 => \N__56529\,
            in3 => \N__56858\,
            lcout => \c0.n13_adj_4492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1424_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__74817\,
            in1 => \N__56526\,
            in2 => \N__59636\,
            in3 => \N__56499\,
            lcout => \c0.n37_adj_4458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_4_lut_adj_1702_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72321\,
            in1 => \N__77872\,
            in2 => \N__73401\,
            in3 => \N__77816\,
            lcout => \c0.n22_adj_4597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i105_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__75493\,
            in1 => \N__75421\,
            in2 => \N__58304\,
            in3 => \N__80615\,
            lcout => \c0.data_in_frame_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i233_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__75420\,
            in1 => \N__56483\,
            in2 => \N__80673\,
            in3 => \N__56684\,
            lcout => \c0.data_in_frame_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i240_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__56482\,
            in1 => \N__76227\,
            in2 => \N__75426\,
            in3 => \N__56904\,
            lcout => \c0.data_in_frame_29_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1429_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56903\,
            in1 => \N__56895\,
            in2 => \_gnd_net_\,
            in3 => \N__56862\,
            lcout => \c0.n12_adj_4466\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1745_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__56817\,
            in1 => \N__77287\,
            in2 => \_gnd_net_\,
            in3 => \N__59561\,
            lcout => OPEN,
            ltout => \c0.n11_adj_4474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1433_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56766\,
            in1 => \N__63226\,
            in2 => \N__56760\,
            in3 => \N__56757\,
            lcout => \c0.n18_adj_4475\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i112_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__75494\,
            in1 => \N__75422\,
            in2 => \N__62847\,
            in3 => \N__76228\,
            lcout => \c0.data_in_frame_13_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1455_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58719\,
            in1 => \N__64134\,
            in2 => \N__56712\,
            in3 => \N__56691\,
            lcout => \c0.n44_adj_4501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_324_2_lut_3_lut_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__56652\,
            in1 => \_gnd_net_\,
            in2 => \N__67152\,
            in3 => \N__57014\,
            lcout => \c0.n25446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1748_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57015\,
            in1 => \N__67147\,
            in2 => \N__56685\,
            in3 => \N__56650\,
            lcout => OPEN,
            ltout => \c0.n43_adj_4463_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i32_4_lut_adj_1426_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__76742\,
            in1 => \N__56669\,
            in2 => \N__56655\,
            in3 => \N__63786\,
            lcout => \c0.n74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_adj_1744_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57016\,
            in1 => \N__67148\,
            in2 => \N__67327\,
            in3 => \N__56651\,
            lcout => \c0.n42_adj_4540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1234_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__67149\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57017\,
            lcout => \c0.n13911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i33_4_lut_adj_1505_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63264\,
            in1 => \N__56973\,
            in2 => \N__59796\,
            in3 => \N__59808\,
            lcout => OPEN,
            ltout => \c0.n23921_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1508_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111101101111"
        )
    port map (
            in0 => \N__56964\,
            in1 => \N__56955\,
            in2 => \N__56949\,
            in3 => \N__57113\,
            lcout => \c0.n21_adj_4547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_2_lut_4_lut_adj_1732_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67559\,
            in1 => \N__68366\,
            in2 => \N__75938\,
            in3 => \N__68280\,
            lcout => \c0.n31_adj_4542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1493_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110111"
        )
    port map (
            in0 => \N__66768\,
            in1 => \N__56934\,
            in2 => \N__68295\,
            in3 => \N__57120\,
            lcout => \c0.n32_adj_4533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i210_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69204\,
            in1 => \N__75138\,
            in2 => \N__63731\,
            in3 => \N__79457\,
            lcout => \c0.data_in_frame_26_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i40_4_lut_adj_1468_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63263\,
            in1 => \N__56910\,
            in2 => \N__75636\,
            in3 => \N__59505\,
            lcout => \c0.n82_adj_4517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i194_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__72989\,
            in1 => \N__75137\,
            in2 => \N__64179\,
            in3 => \N__79456\,
            lcout => \c0.data_in_frame_24_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_1494_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__67297\,
            in1 => \N__77341\,
            in2 => \_gnd_net_\,
            in3 => \N__66831\,
            lcout => \c0.n32_adj_4534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_3_lut_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__64085\,
            in1 => \N__59782\,
            in2 => \_gnd_net_\,
            in3 => \N__59896\,
            lcout => OPEN,
            ltout => \c0.n71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i39_4_lut_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57174\,
            in1 => \N__67033\,
            in2 => \N__57162\,
            in3 => \N__59985\,
            lcout => OPEN,
            ltout => \c0.n81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1480_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111110"
        )
    port map (
            in0 => \N__57155\,
            in1 => \N__59955\,
            in2 => \N__57129\,
            in3 => \N__57126\,
            lcout => \c0.n28_adj_4523\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1492_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57114\,
            in1 => \N__57080\,
            in2 => \_gnd_net_\,
            in3 => \N__67506\,
            lcout => OPEN,
            ltout => \c0.n23_adj_4532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1495_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67797\,
            in1 => \N__77898\,
            in2 => \N__57048\,
            in3 => \N__67819\,
            lcout => OPEN,
            ltout => \c0.n38_adj_4535_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_adj_1502_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67748\,
            in1 => \N__57045\,
            in2 => \N__57039\,
            in3 => \N__57036\,
            lcout => \c0.n15_adj_4497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1978_LC_20_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61380\,
            in2 => \_gnd_net_\,
            in3 => \N__62318\,
            lcout => \c0.n12_adj_4672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1833_LC_21_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69354\,
            in2 => \_gnd_net_\,
            in3 => \N__64531\,
            lcout => \c0.n13998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_adj_1767_LC_21_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__60594\,
            in1 => \N__60204\,
            in2 => \_gnd_net_\,
            in3 => \N__68120\,
            lcout => \c0.n8_adj_4677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i79_LC_21_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__73717\,
            in1 => \N__74150\,
            in2 => \N__57417\,
            in3 => \N__73291\,
            lcout => \c0.data_in_frame_9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i44_LC_21_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__77106\,
            in1 => \N__69462\,
            in2 => \_gnd_net_\,
            in3 => \N__57366\,
            lcout => data_in_frame_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i87_LC_21_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__73718\,
            in1 => \N__69185\,
            in2 => \N__61781\,
            in3 => \N__73292\,
            lcout => \c0.data_in_frame_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i43_LC_21_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__57324\,
            in1 => \N__69461\,
            in2 => \_gnd_net_\,
            in3 => \N__79106\,
            lcout => data_in_frame_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1582_LC_21_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64049\,
            in2 => \_gnd_net_\,
            in3 => \N__69330\,
            lcout => \c0.n7_adj_4603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1609_LC_21_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61044\,
            in1 => \N__57192\,
            in2 => \N__57309\,
            in3 => \N__57245\,
            lcout => \c0.n23554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i45_LC_21_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__57461\,
            in1 => \N__71968\,
            in2 => \_gnd_net_\,
            in3 => \N__69459\,
            lcout => data_in_frame_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1608_LC_21_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57951\,
            in1 => \N__60634\,
            in2 => \N__57447\,
            in3 => \N__60203\,
            lcout => \c0.n12_adj_4612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_4_lut_adj_1662_LC_21_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68928\,
            in1 => \N__64490\,
            in2 => \N__72585\,
            in3 => \N__69584\,
            lcout => \c0.n15_adj_4444\,
            ltout => \c0.n15_adj_4444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i46_4_lut_adj_1407_LC_21_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61466\,
            in1 => \N__57428\,
            in2 => \N__57510\,
            in3 => \N__69492\,
            lcout => \c0.n102_adj_4445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_1672_LC_21_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__60632\,
            in1 => \_gnd_net_\,
            in2 => \N__57462\,
            in3 => \N__57494\,
            lcout => \c0.n11_adj_4656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1668_LC_21_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__57495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57460\,
            lcout => \c0.n6_adj_4611\,
            ltout => \c0.n6_adj_4611_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i35_2_lut_4_lut_LC_21_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60633\,
            in1 => \N__57950\,
            in2 => \N__57438\,
            in3 => \N__61043\,
            lcout => \c0.n91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i57_LC_21_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__80922\,
            in1 => \N__70166\,
            in2 => \N__64502\,
            in3 => \N__80737\,
            lcout => \c0.data_in_frame_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i7_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__70165\,
            in1 => \N__73294\,
            in2 => \N__60648\,
            in3 => \N__72924\,
            lcout => \c0.data_in_frame_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i23_LC_21_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__73293\,
            in1 => \N__70167\,
            in2 => \N__60746\,
            in3 => \N__69150\,
            lcout => \c0.data_in_frame_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1631_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60283\,
            in1 => \N__60737\,
            in2 => \_gnd_net_\,
            in3 => \N__68495\,
            lcout => \c0.n23302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i5_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__68496\,
            in1 => \N__71959\,
            in2 => \N__72966\,
            in3 => \N__70022\,
            lcout => \c0.data_in_frame_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i165_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__79986\,
            in1 => \N__59702\,
            in2 => \N__71969\,
            in3 => \N__80426\,
            lcout => \c0.data_in_frame_20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i6_LC_21_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__60301\,
            in1 => \N__79646\,
            in2 => \N__72967\,
            in3 => \N__70023\,
            lcout => \c0.data_in_frame_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i4_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__70164\,
            in1 => \N__77111\,
            in2 => \N__68121\,
            in3 => \N__72923\,
            lcout => \c0.data_in_frame_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1898_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__67915\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68096\,
            lcout => \c0.n10_adj_4722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1873_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65678\,
            in2 => \_gnd_net_\,
            in3 => \N__57957\,
            lcout => \c0.n15_adj_4450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i22_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69156\,
            in1 => \N__70141\,
            in2 => \N__67943\,
            in3 => \N__79589\,
            lcout => \c0.data_in_frame_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1595_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__67914\,
            in1 => \N__68497\,
            in2 => \_gnd_net_\,
            in3 => \N__68095\,
            lcout => \c0.n13453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i50_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__75186\,
            in1 => \N__68437\,
            in2 => \_gnd_net_\,
            in3 => \N__58128\,
            lcout => data_in_frame_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i164_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__79953\,
            in1 => \N__80425\,
            in2 => \N__75765\,
            in3 => \N__77130\,
            lcout => \c0.data_in_frame_20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_2_lut_4_lut_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57536\,
            in1 => \N__64827\,
            in2 => \N__64902\,
            in3 => \N__64779\,
            lcout => \c0.n61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_1233_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60884\,
            in2 => \_gnd_net_\,
            in3 => \N__62070\,
            lcout => \c0.n17_adj_4224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i54_4_lut_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57864\,
            in1 => \N__57855\,
            in2 => \N__61503\,
            in3 => \N__57849\,
            lcout => OPEN,
            ltout => \c0.n110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i55_4_lut_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57843\,
            in1 => \N__57837\,
            in2 => \N__57825\,
            in3 => \N__57738\,
            lcout => \c0.n24465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1621_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__62071\,
            in1 => \N__57730\,
            in2 => \N__60895\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_frame_0__7__N_2579\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_2_lut_3_lut_4_lut_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57728\,
            in1 => \N__58155\,
            in2 => \N__57800\,
            in3 => \N__60942\,
            lcout => \c0.n87\,
            ltout => \c0.n87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i50_4_lut_adj_1410_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57765\,
            in1 => \N__57753\,
            in2 => \N__57741\,
            in3 => \N__64389\,
            lcout => \c0.n106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1780_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57729\,
            in1 => \N__60883\,
            in2 => \N__61596\,
            in3 => \N__62069\,
            lcout => \c0.n7_adj_4304\,
            ltout => \c0.n7_adj_4304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1283_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__57675\,
            in3 => \N__57661\,
            lcout => \c0.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1902_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58048\,
            in1 => \N__57606\,
            in2 => \N__61083\,
            in3 => \N__71080\,
            lcout => \c0.n27_adj_4725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i49_3_lut_4_lut_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72397\,
            in1 => \N__58253\,
            in2 => \N__72483\,
            in3 => \N__60029\,
            lcout => \c0.n130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1863_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58230\,
            in1 => \N__58212\,
            in2 => \N__58200\,
            in3 => \N__65096\,
            lcout => \c0.n22_adj_4259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_LC_21_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__65706\,
            in1 => \_gnd_net_\,
            in2 => \N__60953\,
            in3 => \N__57960\,
            lcout => \c0.n18_adj_4314\,
            ltout => \c0.n18_adj_4314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_3_lut_4_lut_adj_1678_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71095\,
            in1 => \N__58132\,
            in2 => \N__58101\,
            in3 => \N__58098\,
            lcout => \c0.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_1895_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__71079\,
            in1 => \N__58047\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n22230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1412_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70225\,
            in1 => \N__64345\,
            in2 => \N__65295\,
            in3 => \N__57972\,
            lcout => \c0.n42_adj_4449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_4_lut_4_lut_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65705\,
            in1 => \N__71094\,
            in2 => \N__60952\,
            in3 => \N__57959\,
            lcout => \c0.n24_adj_4689\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_1377_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__78852\,
            in1 => \N__66863\,
            in2 => \N__73038\,
            in3 => \N__57888\,
            lcout => \c0.n41_adj_4360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_2040_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__58447\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__70439\,
            lcout => \c0.n31\,
            ltout => \c0.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_adj_1228_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61293\,
            in1 => \N__58331\,
            in2 => \N__58410\,
            in3 => \N__58407\,
            lcout => \c0.n53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58377\,
            in1 => \N__60558\,
            in2 => \N__58350\,
            in3 => \N__58341\,
            lcout => \c0.n23267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i115_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__79168\,
            in1 => \N__59205\,
            in2 => \_gnd_net_\,
            in3 => \N__58332\,
            lcout => data_in_frame_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1747_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58313\,
            in1 => \N__60557\,
            in2 => \N__58323\,
            in3 => \N__61292\,
            lcout => \c0.n23491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i51_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__68433\,
            in1 => \_gnd_net_\,
            in2 => \N__79193\,
            in3 => \N__58314\,
            lcout => data_in_frame_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__76037\,
            in1 => \N__77845\,
            in2 => \N__76070\,
            in3 => \N__81032\,
            lcout => \c0.n22205\,
            ltout => \c0.n22205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1696_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58305\,
            in1 => \N__60819\,
            in2 => \N__58284\,
            in3 => \N__58279\,
            lcout => \c0.n22589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_3_lut_4_lut_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66053\,
            in1 => \N__77846\,
            in2 => \N__76048\,
            in3 => \N__77776\,
            lcout => \c0.n22_adj_4243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1652_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__72577\,
            in1 => \N__66052\,
            in2 => \_gnd_net_\,
            in3 => \N__69580\,
            lcout => \c0.n23598\,
            ltout => \c0.n23598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1723_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__77844\,
            in2 => \N__58503\,
            in3 => \N__81031\,
            lcout => \c0.n13128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63032\,
            in2 => \_gnd_net_\,
            in3 => \N__72284\,
            lcout => \c0.n9_adj_4208\,
            ltout => \c0.n9_adj_4208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1890_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__73400\,
            in1 => \N__58496\,
            in2 => \N__58485\,
            in3 => \N__77777\,
            lcout => \c0.n22304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61122\,
            in1 => \N__68190\,
            in2 => \N__68879\,
            in3 => \N__62875\,
            lcout => \c0.n107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1883_LC_21_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59260\,
            in1 => \N__59053\,
            in2 => \N__62615\,
            in3 => \N__58472\,
            lcout => \c0.n13892\,
            ltout => \c0.n13892_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1789_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__74714\,
            in1 => \N__66097\,
            in2 => \N__58461\,
            in3 => \N__58872\,
            lcout => \c0.n6215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1604_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__61648\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62808\,
            lcout => \c0.n22662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i95_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76654\,
            in1 => \N__73705\,
            in2 => \N__58451\,
            in3 => \N__73299\,
            lcout => \c0.data_in_frame_11_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1948_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59352\,
            in1 => \N__59081\,
            in2 => \N__58670\,
            in3 => \N__58425\,
            lcout => \c0.n13797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1538_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__74713\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58662\,
            lcout => \c0.n14088\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1223_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72631\,
            in1 => \N__72581\,
            in2 => \N__65748\,
            in3 => \N__65798\,
            lcout => \c0.n22547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1623_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65112\,
            in1 => \N__70926\,
            in2 => \N__58638\,
            in3 => \N__65154\,
            lcout => \c0.n22825\,
            ltout => \c0.n22825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1730_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__72165\,
            in1 => \_gnd_net_\,
            in2 => \N__58623\,
            in3 => \N__72210\,
            lcout => \c0.n22751\,
            ltout => \c0.n22751_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i68_4_lut_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58620\,
            in1 => \N__58587\,
            in2 => \N__58572\,
            in3 => \N__58569\,
            lcout => \c0.n149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1632_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65370\,
            in1 => \N__74962\,
            in2 => \_gnd_net_\,
            in3 => \N__61815\,
            lcout => \c0.n22586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i59_4_lut_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65717\,
            in1 => \N__71116\,
            in2 => \N__65779\,
            in3 => \N__77792\,
            lcout => \c0.n140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1575_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__66096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66565\,
            lcout => \c0.n22843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1224_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61796\,
            in1 => \N__63152\,
            in2 => \N__74718\,
            in3 => \N__61698\,
            lcout => \c0.n22_adj_4245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1279_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__66006\,
            in1 => \N__58700\,
            in2 => \_gnd_net_\,
            in3 => \N__72078\,
            lcout => \c0.n22514\,
            ltout => \c0.n22514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1871_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__58704\,
            in3 => \N__72103\,
            lcout => \c0.n22803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i129_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__80746\,
            in1 => \N__72982\,
            in2 => \N__72110\,
            in3 => \N__80265\,
            lcout => \c0.data_in_frame_16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i130_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__75253\,
            in1 => \N__58701\,
            in2 => \N__72992\,
            in3 => \N__80266\,
            lcout => \c0.data_in_frame_16_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i110_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__79727\,
            in1 => \N__75499\,
            in2 => \N__66016\,
            in3 => \N__75373\,
            lcout => \c0.data_in_frame_13_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i111_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__75498\,
            in1 => \N__73335\,
            in2 => \N__72088\,
            in3 => \N__75374\,
            lcout => \c0.data_in_frame_13_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1534_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__73944\,
            in1 => \N__59724\,
            in2 => \_gnd_net_\,
            in3 => \N__66336\,
            lcout => \c0.n14_adj_4566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1729_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58980\,
            in1 => \N__72681\,
            in2 => \N__58782\,
            in3 => \N__70549\,
            lcout => \c0.n14165\,
            ltout => \c0.n14165_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1521_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__58674\,
            in3 => \N__62360\,
            lcout => \c0.n4_adj_4345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1681_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__58777\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59025\,
            lcout => OPEN,
            ltout => \c0.n4_adj_4658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1786_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__62407\,
            in1 => \N__62483\,
            in2 => \N__58983\,
            in3 => \N__58979\,
            lcout => OPEN,
            ltout => \c0.n12_adj_4682_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1788_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58938\,
            in1 => \N__58725\,
            in2 => \N__58902\,
            in3 => \N__58899\,
            lcout => \c0.n22249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1903_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63430\,
            in1 => \N__63347\,
            in2 => \N__71631\,
            in3 => \N__58854\,
            lcout => \c0.n24534\,
            ltout => \c0.n24534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1366_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58828\,
            in1 => \N__58803\,
            in2 => \N__58797\,
            in3 => \N__62009\,
            lcout => \c0.n12_adj_4346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1618_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__70548\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58778\,
            lcout => \c0.n4_adj_4621\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_1561_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77674\,
            in1 => \N__72123\,
            in2 => \N__77705\,
            in3 => \N__77812\,
            lcout => \c0.n44_adj_4588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_4_lut_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__60061\,
            in1 => \N__72347\,
            in2 => \N__59334\,
            in3 => \N__62687\,
            lcout => \c0.n12_adj_4500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_1892_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65787\,
            in1 => \N__61746\,
            in2 => \N__59058\,
            in3 => \N__61797\,
            lcout => \c0.n6_adj_4587\,
            ltout => \c0.n6_adj_4587_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1889_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77673\,
            in1 => \N__59370\,
            in2 => \N__59355\,
            in3 => \N__77811\,
            lcout => \c0.n13461\,
            ltout => \c0.n13461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1697_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66496\,
            in1 => \N__59329\,
            in2 => \N__59310\,
            in3 => \N__72242\,
            lcout => \c0.n6227\,
            ltout => \c0.n6227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1398_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62686\,
            in2 => \N__59307\,
            in3 => \N__59304\,
            lcout => \c0.n21301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1265_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62424\,
            in1 => \N__62411\,
            in2 => \N__66501\,
            in3 => \N__60060\,
            lcout => \c0.n19_adj_4291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1879_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59261\,
            in1 => \N__62720\,
            in2 => \N__62603\,
            in3 => \N__59088\,
            lcout => \c0.n21414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i120_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__76385\,
            in1 => \N__59148\,
            in2 => \_gnd_net_\,
            in3 => \N__62591\,
            lcout => data_in_frame_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78752\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1548_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59130\,
            in1 => \N__59109\,
            in2 => \N__62331\,
            in3 => \N__62010\,
            lcout => \c0.n23300\,
            ltout => \c0.n23300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1567_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59082\,
            in1 => \N__59057\,
            in2 => \N__59034\,
            in3 => \N__62721\,
            lcout => \c0.n21_adj_4594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1388_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59456\,
            in2 => \_gnd_net_\,
            in3 => \N__67180\,
            lcout => \c0.n4_adj_4347\,
            ltout => \c0.n4_adj_4347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1376_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59484\,
            in1 => \N__80136\,
            in2 => \N__59463\,
            in3 => \N__77229\,
            lcout => \c0.n40_adj_4359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i186_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__80328\,
            in1 => \N__80966\,
            in2 => \N__59460\,
            in3 => \N__75224\,
            lcout => \c0.data_in_frame_23_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78752\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1700_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__73034\,
            in1 => \N__65904\,
            in2 => \_gnd_net_\,
            in3 => \N__63299\,
            lcout => \c0.n22698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_adj_1576_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__66661\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66597\,
            lcout => \c0.n30_adj_4357\,
            ltout => \c0.n30_adj_4357_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1375_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59720\,
            in1 => \N__66950\,
            in2 => \N__59445\,
            in3 => \N__59434\,
            lcout => OPEN,
            ltout => \c0.n42_adj_4358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59403\,
            in1 => \N__61926\,
            in2 => \N__59397\,
            in3 => \N__59394\,
            lcout => \c0.n34_adj_4361\,
            ltout => \c0.n34_adj_4361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1464_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59385\,
            in1 => \N__59376\,
            in2 => \N__59379\,
            in3 => \N__63170\,
            lcout => \c0.n42_adj_4510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1553_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__75847\,
            in2 => \_gnd_net_\,
            in3 => \N__66751\,
            lcout => \c0.n14148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1421_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61927\,
            in1 => \N__66525\,
            in2 => \N__59731\,
            in3 => \N__59676\,
            lcout => \c0.n22426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1527_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67313\,
            in2 => \_gnd_net_\,
            in3 => \N__67260\,
            lcout => \c0.n5_adj_4486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_334_2_lut_4_lut_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67251\,
            in1 => \N__59589\,
            in2 => \N__64168\,
            in3 => \N__67550\,
            lcout => \c0.n25456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1509_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67499\,
            in1 => \N__59663\,
            in2 => \N__59640\,
            in3 => \N__73943\,
            lcout => \c0.n26_adj_4548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1718_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__64158\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59588\,
            lcout => \c0.n13468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1518_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67549\,
            in2 => \_gnd_net_\,
            in3 => \N__67250\,
            lcout => \c0.n13490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_3_lut_4_lut_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__78026\,
            in1 => \N__59562\,
            in2 => \N__59532\,
            in3 => \N__67500\,
            lcout => OPEN,
            ltout => \c0.n66_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i33_4_lut_adj_1427_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67314\,
            in1 => \N__59499\,
            in2 => \N__59508\,
            in3 => \N__63599\,
            lcout => \c0.n75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__77376\,
            in1 => \N__74893\,
            in2 => \_gnd_net_\,
            in3 => \N__67593\,
            lcout => \c0.n46_adj_4461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_adj_1927_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__63230\,
            in1 => \N__68312\,
            in2 => \_gnd_net_\,
            in3 => \N__63636\,
            lcout => \c0.n25_adj_4469\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1499_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67089\,
            in1 => \N__59919\,
            in2 => \N__59787\,
            in3 => \N__59897\,
            lcout => \c0.n53_adj_4538\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1510_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__74778\,
            in1 => \N__67592\,
            in2 => \N__59880\,
            in3 => \N__63598\,
            lcout => OPEN,
            ltout => \c0.n24_adj_4550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1511_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59838\,
            in1 => \N__59826\,
            in2 => \N__59820\,
            in3 => \N__73773\,
            lcout => \c0.n21010\,
            ltout => \c0.n21010_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64089\,
            in1 => \N__63686\,
            in2 => \N__59817\,
            in3 => \N__59814\,
            lcout => \c0.n61_adj_4543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_adj_1501_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59802\,
            in1 => \N__63567\,
            in2 => \N__63739\,
            in3 => \N__63849\,
            lcout => \c0.n62_adj_4541\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_adj_1450_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64138\,
            in2 => \N__67873\,
            in3 => \N__59786\,
            lcout => \c0.n18_adj_4493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1454_LC_21_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59763\,
            in1 => \N__63791\,
            in2 => \N__75702\,
            in3 => \N__63642\,
            lcout => OPEN,
            ltout => \c0.n26_adj_4499_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1458_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62553\,
            in1 => \N__59754\,
            in2 => \N__59745\,
            in3 => \N__63848\,
            lcout => OPEN,
            ltout => \c0.n24441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1506_LC_21_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__63453\,
            in1 => \N__63855\,
            in2 => \N__60003\,
            in3 => \N__67398\,
            lcout => \c0.n30_adj_4545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i30_4_lut_adj_1467_LC_21_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63680\,
            in1 => \N__63847\,
            in2 => \N__63741\,
            in3 => \N__63653\,
            lcout => \c0.n72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i177_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__63499\,
            in1 => \N__80672\,
            in2 => \_gnd_net_\,
            in3 => \N__78915\,
            lcout => data_in_frame_22_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1469_LC_21_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__59979\,
            in1 => \N__67005\,
            in2 => \N__59967\,
            in3 => \N__63810\,
            lcout => \c0.n20_adj_4518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i227_LC_21_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__80079\,
            in1 => \N__79167\,
            in2 => \N__63828\,
            in3 => \N__79482\,
            lcout => \c0.data_in_frame_28_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78797\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20984_4_lut_LC_22_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__67941\,
            in1 => \N__60644\,
            in2 => \N__60798\,
            in3 => \N__60304\,
            lcout => \c0.n24751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1839_LC_22_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64033\,
            in2 => \_gnd_net_\,
            in3 => \N__61767\,
            lcout => \c0.n6_adj_4632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1766_LC_22_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__60303\,
            in1 => \N__60208\,
            in2 => \N__68543\,
            in3 => \N__60637\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1768_LC_22_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__69582\,
            in1 => \N__64068\,
            in2 => \N__59934\,
            in3 => \N__68094\,
            lcout => \c0.data_out_frame_0__7__N_2777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1762_LC_22_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__68849\,
            in1 => \N__60636\,
            in2 => \N__68542\,
            in3 => \N__69581\,
            lcout => \c0.n24016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20982_4_lut_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__69583\,
            in1 => \N__64778\,
            in2 => \N__60228\,
            in3 => \N__68795\,
            lcout => \c0.n24749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1935_LC_22_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__68848\,
            in1 => \N__60566\,
            in2 => \N__72586\,
            in3 => \N__60431\,
            lcout => \c0.n37_adj_4738\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1881_LC_22_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72570\,
            in1 => \N__60302\,
            in2 => \N__60227\,
            in3 => \N__68093\,
            lcout => \c0.n24_adj_4717\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_2049_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__60155\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61262\,
            lcout => OPEN,
            ltout => \c0.n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60012\,
            in1 => \N__60135\,
            in2 => \N__60120\,
            in3 => \N__60117\,
            lcout => OPEN,
            ltout => \c0.n54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_4_lut_adj_1230_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60099\,
            in1 => \N__60654\,
            in2 => \N__60087\,
            in3 => \N__60084\,
            lcout => \c0.n13821\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69894\,
            in1 => \N__64008\,
            in2 => \N__64229\,
            in3 => \N__68141\,
            lcout => \c0.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_adj_1865_LC_22_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68840\,
            in2 => \_gnd_net_\,
            in3 => \N__68081\,
            lcout => \c0.n37\,
            ltout => \c0.n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1869_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64012\,
            in1 => \N__68028\,
            in2 => \N__60753\,
            in3 => \N__68140\,
            lcout => \c0.n22647\,
            ltout => \c0.n22647_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1877_LC_22_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__60750\,
            in3 => \N__68958\,
            lcout => \c0.n16_adj_4716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20980_4_lut_LC_22_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__68082\,
            in1 => \N__68752\,
            in2 => \N__60747\,
            in3 => \N__68029\,
            lcout => \c0.n24747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_adj_1614_LC_22_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68733\,
            in1 => \N__68512\,
            in2 => \N__65696\,
            in3 => \N__68846\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4616_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1899_LC_22_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68781\,
            in1 => \N__60699\,
            in2 => \N__60693\,
            in3 => \N__64006\,
            lcout => \c0.data_out_frame_0__7__N_2743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i38_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__79588\,
            in1 => \N__79988\,
            in2 => \N__65697\,
            in3 => \N__70146\,
            lcout => \c0.data_in_frame_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_LC_22_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64293\,
            in1 => \N__60690\,
            in2 => \N__60666\,
            in3 => \N__68034\,
            lcout => \c0.n55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i33_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__80742\,
            in1 => \N__79987\,
            in2 => \N__60899\,
            in3 => \N__70145\,
            lcout => \c0.data_in_frame_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1864_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__68780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68671\,
            lcout => \c0.n5_adj_4711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_LC_22_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60891\,
            in1 => \N__61101\,
            in2 => \_gnd_net_\,
            in3 => \N__60854\,
            lcout => \c0.n24_adj_4724\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i39_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__70144\,
            in1 => \N__73289\,
            in2 => \N__80032\,
            in3 => \N__64007\,
            lcout => \c0.data_in_frame_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1882_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61057\,
            in1 => \N__60987\,
            in2 => \N__60796\,
            in3 => \N__60912\,
            lcout => OPEN,
            ltout => \c0.n28_adj_4718_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1891_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60981\,
            in1 => \N__68531\,
            in2 => \N__60969\,
            in3 => \N__60966\,
            lcout => \c0.n23_adj_4599\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1872_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64259\,
            in2 => \_gnd_net_\,
            in3 => \N__69546\,
            lcout => \c0.n4_adj_4446\,
            ltout => \c0.n4_adj_4446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_1876_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68727\,
            in2 => \N__60915\,
            in3 => \N__61288\,
            lcout => \c0.n26_adj_4714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i17_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__80741\,
            in1 => \N__70018\,
            in2 => \N__60797\,
            in3 => \N__69091\,
            lcout => \c0.data_in_frame_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1757_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60774\,
            in1 => \N__60882\,
            in2 => \_gnd_net_\,
            in3 => \N__60855\,
            lcout => \c0.n23597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1705_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68959\,
            in1 => \N__60773\,
            in2 => \N__61298\,
            in3 => \N__64260\,
            lcout => \c0.n10_adj_4664\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_3_lut_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__61255\,
            in1 => \N__70694\,
            in2 => \_gnd_net_\,
            in3 => \N__67985\,
            lcout => \c0.n48_adj_4227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i69_4_lut_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61113\,
            in1 => \N__70715\,
            in2 => \N__65369\,
            in3 => \N__69700\,
            lcout => \c0.n150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_1179_LC_22_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65201\,
            in2 => \_gnd_net_\,
            in3 => \N__65220\,
            lcout => \c0.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_1665_LC_22_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65221\,
            in1 => \N__65202\,
            in2 => \_gnd_net_\,
            in3 => \N__65108\,
            lcout => \c0.n13651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1200_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64562\,
            in1 => \N__61111\,
            in2 => \N__64686\,
            in3 => \N__71119\,
            lcout => OPEN,
            ltout => \c0.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_3_lut_LC_22_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61175\,
            in2 => \N__61152\,
            in3 => \N__61149\,
            lcout => \c0.n23528\,
            ltout => \c0.n23528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_22_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65988\,
            in1 => \N__64967\,
            in2 => \N__61128\,
            in3 => \N__61341\,
            lcout => OPEN,
            ltout => \c0.n34_adj_4278_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1259_LC_22_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66227\,
            in1 => \N__68604\,
            in2 => \N__61125\,
            in3 => \N__68532\,
            lcout => \c0.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_2_lut_LC_22_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__64563\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61112\,
            lcout => \c0.n60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1848_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62119\,
            in1 => \N__71209\,
            in2 => \N__64966\,
            in3 => \N__71118\,
            lcout => OPEN,
            ltout => \c0.n30_adj_4705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1850_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69758\,
            in1 => \N__69693\,
            in2 => \N__61347\,
            in3 => \N__62033\,
            lcout => \c0.n23523\,
            ltout => \c0.n23523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65591\,
            in2 => \N__61344\,
            in3 => \N__65549\,
            lcout => \c0.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1728_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__66246\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65525\,
            lcout => \c0.n4_adj_4261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i99_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__80060\,
            in1 => \N__73665\,
            in2 => \N__65039\,
            in3 => \N__79209\,
            lcout => \c0.data_in_frame_12_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_2013_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__64191\,
            in1 => \N__70672\,
            in2 => \_gnd_net_\,
            in3 => \N__65638\,
            lcout => \c0.n6_adj_4209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i72_LC_22_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__76378\,
            in1 => \N__65639\,
            in2 => \N__72978\,
            in3 => \N__73666\,
            lcout => \c0.data_in_frame_8_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1838_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65631\,
            in1 => \N__61333\,
            in2 => \N__61479\,
            in3 => \N__61488\,
            lcout => \c0.n7_adj_4634\,
            ltout => \c0.n7_adj_4634_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1775_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71177\,
            in1 => \N__70958\,
            in2 => \N__61305\,
            in3 => \N__65297\,
            lcout => \c0.n5807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1776_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65296\,
            in1 => \N__64506\,
            in2 => \N__71176\,
            in3 => \N__61738\,
            lcout => \c0.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i40_4_lut_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61589\,
            in1 => \N__61782\,
            in2 => \N__61745\,
            in3 => \N__65630\,
            lcout => OPEN,
            ltout => \c0.n96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i48_4_lut_adj_1406_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61475\,
            in1 => \N__61487\,
            in2 => \N__61560\,
            in3 => \N__61557\,
            lcout => \c0.n104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1242_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69301\,
            in2 => \_gnd_net_\,
            in3 => \N__70618\,
            lcout => \c0.n7_adj_4253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i52_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__68432\,
            in1 => \_gnd_net_\,
            in2 => \N__77121\,
            in3 => \N__77856\,
            lcout => data_in_frame_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1241_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__76036\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65327\,
            lcout => \c0.n5_adj_4252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1676_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61852\,
            in1 => \N__61467\,
            in2 => \N__65337\,
            in3 => \N__65226\,
            lcout => \c0.n13734\,
            ltout => \c0.n13734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_1675_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__61741\,
            in1 => \_gnd_net_\,
            in2 => \N__61440\,
            in3 => \N__65772\,
            lcout => \c0.n18_adj_4580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1719_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__61437\,
            in1 => \N__61392\,
            in2 => \_gnd_net_\,
            in3 => \N__62271\,
            lcout => \c0.n22120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1656_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65331\,
            in2 => \_gnd_net_\,
            in3 => \N__61851\,
            lcout => \c0.n22176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1583_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64373\,
            in1 => \N__65150\,
            in2 => \N__61833\,
            in3 => \N__65111\,
            lcout => \c0.n13738\,
            ltout => \c0.n13738_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1893_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61811\,
            in1 => \N__61739\,
            in2 => \N__61800\,
            in3 => \N__61792\,
            lcout => \c0.n22782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1667_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__61740\,
            in1 => \N__61691\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n5_adj_4310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_1855_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62141\,
            in2 => \_gnd_net_\,
            in3 => \N__62132\,
            lcout => OPEN,
            ltout => \c0.n39_adj_4708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_adj_1857_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66161\,
            in1 => \N__62799\,
            in2 => \N__61680\,
            in3 => \N__61629\,
            lcout => OPEN,
            ltout => \c0.n64_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i34_4_lut_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61677\,
            in1 => \N__69765\,
            in2 => \N__61662\,
            in3 => \N__69701\,
            lcout => \c0.n70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1856_LC_22_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72468\,
            in1 => \N__66010\,
            in2 => \N__61659\,
            in3 => \N__65435\,
            lcout => \c0.n55_adj_4709\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1227_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68982\,
            in1 => \N__65009\,
            in2 => \N__61623\,
            in3 => \N__64655\,
            lcout => \c0.n10_adj_4247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i43_4_lut_LC_22_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__73392\,
            in1 => \N__62742\,
            in2 => \N__62806\,
            in3 => \N__66464\,
            lcout => \c0.n124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1417_LC_22_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65436\,
            in1 => \N__62142\,
            in2 => \N__62807\,
            in3 => \N__62133\,
            lcout => \c0.n12_adj_4455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62124\,
            in1 => \N__62886\,
            in2 => \N__64989\,
            in3 => \N__62091\,
            lcout => OPEN,
            ltout => \c0.n59_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i35_4_lut_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62052\,
            in1 => \N__62037\,
            in2 => \N__62022\,
            in3 => \N__62019\,
            lcout => \c0.n24444\,
            ltout => \c0.n24444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__62919\,
            in1 => \N__62887\,
            in2 => \N__62013\,
            in3 => \N__62756\,
            lcout => \c0.n13604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1523_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__62757\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62356\,
            lcout => \c0.n21282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1264_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61995\,
            in2 => \N__62361\,
            in3 => \N__62758\,
            lcout => \c0.n23224\,
            ltout => \c0.n23224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_2028_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__61949\,
            in1 => \N__66608\,
            in2 => \N__61938\,
            in3 => \N__66364\,
            lcout => \c0.n21409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1577_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__61902\,
            in1 => \N__62710\,
            in2 => \N__66117\,
            in3 => \N__62688\,
            lcout => \c0.n10_adj_4602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_2027_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__72021\,
            in1 => \N__66335\,
            in2 => \N__69645\,
            in3 => \N__66365\,
            lcout => \c0.n21404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1630_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__62355\,
            in1 => \N__62613\,
            in2 => \N__62643\,
            in3 => \N__66133\,
            lcout => \c0.n10_adj_4630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_2034_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__62639\,
            in1 => \N__62994\,
            in2 => \N__62616\,
            in3 => \N__62354\,
            lcout => \c0.n12_adj_4246\,
            ltout => \c0.n12_adj_4246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1419_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71646\,
            in1 => \N__62766\,
            in2 => \N__62559\,
            in3 => \N__66134\,
            lcout => \c0.n23691\,
            ltout => \c0.n23691_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1371_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__62556\,
            in3 => \N__66871\,
            lcout => \c0.n20543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1581_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__62532\,
            in1 => \N__62493\,
            in2 => \_gnd_net_\,
            in3 => \N__62487\,
            lcout => \c0.n14189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_1706_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__62463\,
            in1 => \N__62423\,
            in2 => \N__62412\,
            in3 => \N__62353\,
            lcout => \c0.n7_adj_4581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_3_i3_2_lut_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62295\,
            in2 => \_gnd_net_\,
            in3 => \N__71537\,
            lcout => \c0.n3_adj_4430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_1852_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62920\,
            in2 => \_gnd_net_\,
            in3 => \N__62894\,
            lcout => \c0.n20467\,
            ltout => \c0.n20467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_adj_1754_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__62768\,
            in1 => \N__62939\,
            in2 => \N__62985\,
            in3 => \N__75939\,
            lcout => \c0.n17_adj_4354\,
            ltout => \c0.n17_adj_4354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_1373_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63522\,
            in1 => \N__62981\,
            in2 => \N__62943\,
            in3 => \N__67351\,
            lcout => \c0.n58_adj_4355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1689_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62769\,
            in1 => \N__62940\,
            in2 => \N__62927\,
            in3 => \N__62895\,
            lcout => \c0.n21295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3286_2_lut_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__72089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62848\,
            lcout => \c0.n5965\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i103_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__80016\,
            in1 => \N__73708\,
            in2 => \N__73347\,
            in3 => \N__62795\,
            lcout => \c0.data_in_frame_12_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i183_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__63523\,
            in1 => \N__73331\,
            in2 => \_gnd_net_\,
            in3 => \N__78904\,
            lcout => data_in_frame_22_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1225_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62767\,
            in1 => \N__66135\,
            in2 => \N__77209\,
            in3 => \N__62727\,
            lcout => \c0.n21299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1547_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63108\,
            in1 => \N__63120\,
            in2 => \N__72594\,
            in3 => \N__66033\,
            lcout => \c0.n23453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_2_lut_4_lut_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72319\,
            in1 => \N__77879\,
            in2 => \N__63156\,
            in3 => \N__77810\,
            lcout => \c0.n25_adj_4579\,
            ltout => \c0.n25_adj_4579_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1707_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63096\,
            in1 => \N__66032\,
            in2 => \N__63114\,
            in3 => \N__65385\,
            lcout => \c0.n23433\,
            ltout => \c0.n23433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_4_lut_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__72320\,
            in1 => \_gnd_net_\,
            in2 => \N__63111\,
            in3 => \N__77578\,
            lcout => \c0.n43_adj_4661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_3_lut_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__63107\,
            in1 => \_gnd_net_\,
            in2 => \N__74963\,
            in3 => \N__65427\,
            lcout => \c0.n24_adj_4655\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_1910_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63090\,
            in1 => \N__63069\,
            in2 => \N__63063\,
            in3 => \N__65814\,
            lcout => OPEN,
            ltout => \c0.n50_adj_4340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_adj_1361_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63051\,
            in1 => \N__63039\,
            in2 => \N__63021\,
            in3 => \N__66375\,
            lcout => \c0.n28_adj_4343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1571_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65903\,
            in2 => \_gnd_net_\,
            in3 => \N__63295\,
            lcout => \c0.n22375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1448_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63011\,
            in1 => \N__67082\,
            in2 => \N__75700\,
            in3 => \N__63790\,
            lcout => \c0.n39_adj_4487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1965_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__63345\,
            in1 => \N__63379\,
            in2 => \_gnd_net_\,
            in3 => \N__66919\,
            lcout => \c0.n12559\,
            ltout => \c0.n12559_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_1731_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__73033\,
            in1 => \N__66750\,
            in2 => \N__63474\,
            in3 => \N__63464\,
            lcout => \c0.n21316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1457_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__68365\,
            in1 => \N__77307\,
            in2 => \_gnd_net_\,
            in3 => \N__66827\,
            lcout => \c0.n24451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1966_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__66985\,
            in1 => \N__63346\,
            in2 => \_gnd_net_\,
            in3 => \N__63380\,
            lcout => \c0.n6_adj_4459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63440\,
            in1 => \N__63378\,
            in2 => \N__63348\,
            in3 => \N__65862\,
            lcout => \c0.n21275\,
            ltout => \c0.n21275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1400_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__63279\,
            in3 => \N__80135\,
            lcout => \c0.n14_adj_4440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_2_lut_4_lut_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63635\,
            in1 => \N__67056\,
            in2 => \N__63174\,
            in3 => \N__77955\,
            lcout => \c0.n63_adj_4516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__78018\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__67491\,
            lcout => \c0.n48_adj_4365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_2_lut_3_lut_adj_1921_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__63211\,
            in1 => \N__67163\,
            in2 => \_gnd_net_\,
            in3 => \N__68311\,
            lcout => \c0.n46\,
            ltout => \c0.n46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_3_lut_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__77938\,
            in2 => \N__63159\,
            in3 => \N__63634\,
            lcout => OPEN,
            ltout => \c0.n57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1381_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72366\,
            in1 => \N__66998\,
            in2 => \N__63621\,
            in3 => \N__63618\,
            lcout => \c0.n21426\,
            ltout => \c0.n21426_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1753_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74815\,
            in2 => \N__63612\,
            in3 => \N__63782\,
            lcout => \c0.n23032\,
            ltout => \c0.n23032_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1532_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__73809\,
            in1 => \N__73797\,
            in2 => \N__63582\,
            in3 => \N__67591\,
            lcout => \c0.n23209\,
            ltout => \c0.n23209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_adj_1441_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__78019\,
            in1 => \N__63579\,
            in2 => \N__63570\,
            in3 => \N__67492\,
            lcout => \c0.n56_adj_4479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1928_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77190\,
            in1 => \N__77730\,
            in2 => \N__73908\,
            in3 => \N__63561\,
            lcout => \c0.n20802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_1555_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63543\,
            in2 => \_gnd_net_\,
            in3 => \N__67164\,
            lcout => \c0.n26_adj_4470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i175_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67214\,
            in1 => \N__73326\,
            in2 => \_gnd_net_\,
            in3 => \N__67664\,
            lcout => data_in_frame_21_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1558_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63506\,
            in1 => \N__77151\,
            in2 => \N__67218\,
            in3 => \N__66899\,
            lcout => \c0.n22340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1380_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74811\,
            in2 => \_gnd_net_\,
            in3 => \N__63787\,
            lcout => OPEN,
            ltout => \c0.n7_adj_4364_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1422_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__67213\,
            in1 => \N__63972\,
            in2 => \N__63945\,
            in3 => \N__63932\,
            lcout => \c0.n23031\,
            ltout => \c0.n23031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_1430_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__77958\,
            in1 => \N__63727\,
            in2 => \N__63921\,
            in3 => \N__63918\,
            lcout => \c0.n39_adj_4467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1461_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63685\,
            in1 => \N__74904\,
            in2 => \N__63888\,
            in3 => \N__68247\,
            lcout => \c0.n24482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1425_LC_22_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63803\,
            in1 => \N__63788\,
            in2 => \N__63740\,
            in3 => \N__63846\,
            lcout => OPEN,
            ltout => \c0.n36_adj_4460_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_1465_LC_22_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63824\,
            in1 => \N__77957\,
            in2 => \N__63813\,
            in3 => \N__72372\,
            lcout => \c0.n41_adj_4511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1431_LC_22_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63804\,
            in1 => \N__74816\,
            in2 => \N__63687\,
            in3 => \N__63789\,
            lcout => \c0.n38_adj_4468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1554_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__64177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66811\,
            lcout => \c0.n5_adj_4472\,
            ltout => \c0.n5_adj_4472_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1452_LC_22_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63735\,
            in1 => \N__63684\,
            in2 => \N__63657\,
            in3 => \N__63654\,
            lcout => \c0.n24_adj_4496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1738_LC_22_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64178\,
            in1 => \N__66812\,
            in2 => \N__67863\,
            in3 => \N__64143\,
            lcout => \c0.n39_adj_4515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_87_i9_2_lut_3_lut_LC_23_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__74348\,
            in1 => \N__74642\,
            in2 => \_gnd_net_\,
            in3 => \N__74507\,
            lcout => \c0.n9_adj_4552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1764_LC_23_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68751\,
            in2 => \_gnd_net_\,
            in3 => \N__68850\,
            lcout => \c0.n10_adj_4675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i89_LC_23_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76629\,
            in1 => \N__73716\,
            in2 => \N__64048\,
            in3 => \N__80740\,
            lcout => \c0.data_in_frame_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_2022_LC_23_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68108\,
            in1 => \N__68030\,
            in2 => \N__64013\,
            in3 => \N__68841\,
            lcout => \c0.n23282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1605_LC_23_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__68842\,
            in1 => \_gnd_net_\,
            in2 => \N__68039\,
            in3 => \N__68110\,
            lcout => \c0.n23283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1969_LC_23_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67968\,
            in1 => \N__64491\,
            in2 => \N__64544\,
            in3 => \N__68215\,
            lcout => \c0.n8_adj_4216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i37_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__70081\,
            in1 => \N__68677\,
            in2 => \N__79954\,
            in3 => \N__71945\,
            lcout => \c0.data_in_frame_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i20_LC_23_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__77110\,
            in1 => \N__70082\,
            in2 => \N__68796\,
            in3 => \N__69211\,
            lcout => \c0.data_in_frame_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i21_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__69210\,
            in1 => \N__68038\,
            in2 => \N__70150\,
            in3 => \N__71944\,
            lcout => \c0.data_in_frame_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i3_LC_23_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__72925\,
            in1 => \N__70083\,
            in2 => \N__79204\,
            in3 => \N__68843\,
            lcout => \c0.data_in_frame_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1330_LC_23_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67942\,
            in1 => \N__68527\,
            in2 => \N__64901\,
            in3 => \N__68109\,
            lcout => \c0.n21_adj_4327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1602_LC_23_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68161\,
            in1 => \N__64819\,
            in2 => \N__70277\,
            in3 => \N__64212\,
            lcout => \c0.n7_adj_4226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1546_LC_23_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__64818\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68162\,
            lcout => \c0.n4_adj_4211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i40_LC_23_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__70142\,
            in1 => \N__80030\,
            in2 => \N__76294\,
            in3 => \N__64820\,
            lcout => \c0.data_in_frame_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i36_LC_23_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__80029\,
            in1 => \N__70143\,
            in2 => \N__68969\,
            in3 => \N__77131\,
            lcout => \c0.data_in_frame_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1713_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__68160\,
            in1 => \N__64817\,
            in2 => \_gnd_net_\,
            in3 => \N__64211\,
            lcout => \c0.n13904\,
            ltout => \c0.n13904_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1328_LC_23_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67967\,
            in1 => \N__69480\,
            in2 => \N__64203\,
            in3 => \N__68645\,
            lcout => OPEN,
            ltout => \c0.n19_adj_4324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_1343_LC_23_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64200\,
            in2 => \N__64194\,
            in3 => \N__68889\,
            lcout => \c0.n22417\,
            ltout => \c0.n22417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i30_4_lut_LC_23_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64457\,
            in1 => \N__64360\,
            in2 => \N__64416\,
            in3 => \N__64413\,
            lcout => \c0.n86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_4_lut_LC_23_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69549\,
            in1 => \N__69481\,
            in2 => \N__68927\,
            in3 => \N__72563\,
            lcout => \c0.n13085\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_3_lut_4_lut_LC_23_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69788\,
            in1 => \N__70215\,
            in2 => \N__69832\,
            in3 => \N__64341\,
            lcout => \c0.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1997_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__74525\,
            in1 => \N__74632\,
            in2 => \N__74381\,
            in3 => \N__70014\,
            lcout => n22121,
            ltout => \n22121_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i55_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__64283\,
            in1 => \_gnd_net_\,
            in2 => \N__64287\,
            in3 => \N__73290\,
            lcout => data_in_frame_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i2_LC_23_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__72936\,
            in1 => \N__70016\,
            in2 => \N__68756\,
            in3 => \N__75250\,
            lcout => \c0.data_in_frame_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_LC_23_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68726\,
            in1 => \N__69548\,
            in2 => \N__64284\,
            in3 => \N__64261\,
            lcout => \c0.n22322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i19_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__64262\,
            in1 => \N__79205\,
            in2 => \N__69170\,
            in3 => \N__70017\,
            lcout => \c0.data_in_frame_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i1_LC_23_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__70015\,
            in1 => \N__72937\,
            in2 => \N__80735\,
            in3 => \N__69550\,
            lcout => \c0.data_in_frame_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_3_lut_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__64897\,
            in1 => \_gnd_net_\,
            in2 => \N__64838\,
            in3 => \N__64777\,
            lcout => \c0.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_2001_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__70659\,
            in1 => \N__65637\,
            in2 => \_gnd_net_\,
            in3 => \N__67986\,
            lcout => \c0.n20_adj_4260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64965\,
            in2 => \_gnd_net_\,
            in3 => \N__64673\,
            lcout => \c0.n7_adj_4229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_23_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65336\,
            in1 => \N__70915\,
            in2 => \N__69384\,
            in3 => \N__77857\,
            lcout => \c0.n17_adj_4219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_1194_LC_23_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__64634\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__70887\,
            lcout => \c0.n9_adj_4220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_2_lut_3_lut_4_lut_LC_23_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70886\,
            in1 => \N__64633\,
            in2 => \N__69884\,
            in3 => \N__64605\,
            lcout => \c0.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1711_LC_23_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68732\,
            in2 => \N__64554\,
            in3 => \N__69557\,
            lcout => \c0.n23406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i125_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__80923\,
            in1 => \N__73667\,
            in2 => \N__66273\,
            in3 => \N__71781\,
            lcout => \c0.data_in_frame_15_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1190_LC_23_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64545\,
            in2 => \_gnd_net_\,
            in3 => \N__64501\,
            lcout => \c0.n22650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1598_LC_23_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65222\,
            in1 => \N__65200\,
            in2 => \N__70598\,
            in3 => \N__65110\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4609_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1615_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70498\,
            in1 => \N__65160\,
            in2 => \N__65163\,
            in3 => \N__69321\,
            lcout => \c0.n22748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1974_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65633\,
            in1 => \N__70645\,
            in2 => \_gnd_net_\,
            in3 => \N__65127\,
            lcout => \c0.n10_adj_4617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_2014_LC_23_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70591\,
            in1 => \N__65632\,
            in2 => \N__70658\,
            in3 => \N__65143\,
            lcout => OPEN,
            ltout => \c0.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1192_LC_23_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69320\,
            in1 => \N__65126\,
            in2 => \N__65115\,
            in3 => \N__65109\,
            lcout => \c0.n5813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1201_LC_23_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__70527\,
            in1 => \_gnd_net_\,
            in2 => \N__65035\,
            in3 => \_gnd_net_\,
            lcout => \c0.n13809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i94_LC_23_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76674\,
            in1 => \N__73696\,
            in2 => \N__64987\,
            in3 => \N__79698\,
            lcout => \c0.data_in_frame_11_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i127_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__73692\,
            in1 => \N__80941\,
            in2 => \N__70506\,
            in3 => \N__73336\,
            lcout => \c0.data_in_frame_15_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1515_LC_23_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64914\,
            in1 => \N__69609\,
            in2 => \N__70458\,
            in3 => \N__70469\,
            lcout => \c0.n22508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i73_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__73694\,
            in1 => \N__74178\,
            in2 => \N__80747\,
            in3 => \N__70620\,
            lcout => \c0.data_in_frame_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_adj_1861_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72559\,
            in1 => \N__71268\,
            in2 => \N__72482\,
            in3 => \N__72396\,
            lcout => \c0.n23_adj_4665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i123_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__80940\,
            in1 => \N__73695\,
            in2 => \N__65368\,
            in3 => \N__79185\,
            lcout => \c0.data_in_frame_15_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i71_LC_23_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__73693\,
            in1 => \N__72940\,
            in2 => \N__69325\,
            in3 => \N__73337\,
            lcout => \c0.data_in_frame_8_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i70_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__73688\,
            in1 => \N__72941\,
            in2 => \N__79728\,
            in3 => \N__65335\,
            lcout => \c0.data_in_frame_8_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1637_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68634\,
            in1 => \N__70899\,
            in2 => \N__65304\,
            in3 => \N__65654\,
            lcout => OPEN,
            ltout => \c0.n28_adj_4637_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1638_LC_23_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65253\,
            in1 => \N__65244\,
            in2 => \N__65247\,
            in3 => \N__65232\,
            lcout => \c0.n22319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1636_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65493\,
            in1 => \N__69380\,
            in2 => \N__65511\,
            in3 => \N__70848\,
            lcout => \c0.n24_adj_4636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1635_LC_23_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__66271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65238\,
            lcout => \c0.n16_adj_4635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1807_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__68679\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65704\,
            lcout => \c0.n5_adj_4631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1596_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65703\,
            in1 => \N__68633\,
            in2 => \N__65655\,
            in3 => \N__68678\,
            lcout => \c0.n13474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1191_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69313\,
            in2 => \_gnd_net_\,
            in3 => \N__65640\,
            lcout => \c0.n22602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1984_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68189\,
            in1 => \N__65595\,
            in2 => \N__65580\,
            in3 => \N__65553\,
            lcout => \c0.n31_adj_4743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1193_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70847\,
            in1 => \N__65526\,
            in2 => \N__65510\,
            in3 => \N__65492\,
            lcout => OPEN,
            ltout => \c0.n16_adj_4218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_4_lut_adj_1769_LC_23_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__76082\,
            in1 => \N__65475\,
            in2 => \N__65466\,
            in3 => \N__81057\,
            lcout => \c0.n13767\,
            ltout => \c0.n13767_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1716_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71675\,
            in1 => \N__72196\,
            in2 => \N__65463\,
            in3 => \N__65453\,
            lcout => \c0.n6_adj_4454\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1679_LC_23_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74961\,
            in2 => \_gnd_net_\,
            in3 => \N__65419\,
            lcout => \c0.n14_adj_4619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1418_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66018\,
            in1 => \N__66189\,
            in2 => \N__66183\,
            in3 => \N__66162\,
            lcout => \c0.n23507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i169_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__80733\,
            in1 => \N__66116\,
            in2 => \_gnd_net_\,
            in3 => \N__67657\,
            lcout => data_in_frame_21_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i137_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__74187\,
            in1 => \N__80395\,
            in2 => \N__66098\,
            in3 => \N__80734\,
            lcout => \c0.data_in_frame_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_2_lut_3_lut_adj_2024_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__72638\,
            in1 => \N__76052\,
            in2 => \_gnd_net_\,
            in3 => \N__66060\,
            lcout => \c0.n26_adj_4578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1239_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65980\,
            in2 => \_gnd_net_\,
            in3 => \N__66017\,
            lcout => \c0.n22518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i144_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__74188\,
            in1 => \N__76393\,
            in2 => \N__65987\,
            in3 => \N__80396\,
            lcout => \c0.data_in_frame_17_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1350_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__65959\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65931\,
            lcout => \c0.n5_adj_4335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1562_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__71645\,
            in1 => \N__72036\,
            in2 => \N__65902\,
            in3 => \N__65861\,
            lcout => \c0.n42_adj_4589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_4_lut_adj_1693_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65805\,
            in1 => \N__65786\,
            in2 => \N__65747\,
            in3 => \N__65721\,
            lcout => \c0.n24_adj_4618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i180_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__77044\,
            in1 => \N__73750\,
            in2 => \_gnd_net_\,
            in3 => \N__78895\,
            lcout => data_in_frame_22_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1240_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72017\,
            in2 => \_gnd_net_\,
            in3 => \N__66355\,
            lcout => \c0.n7_adj_4251\,
            ltout => \c0.n7_adj_4251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1537_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__75778\,
            in1 => \N__69630\,
            in2 => \N__66339\,
            in3 => \N__66333\,
            lcout => \c0.n4_adj_4568\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1516_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66334\,
            in1 => \N__66393\,
            in2 => \N__69640\,
            in3 => \N__66315\,
            lcout => \c0.n21412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i184_LC_23_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__78896\,
            in1 => \N__76289\,
            in2 => \_gnd_net_\,
            in3 => \N__66302\,
            lcout => data_in_frame_22_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i142_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__74205\,
            in1 => \N__79759\,
            in2 => \N__66500\,
            in3 => \N__80415\,
            lcout => \c0.data_in_frame_17_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1626_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66288\,
            in1 => \N__66272\,
            in2 => \N__67071\,
            in3 => \N__69608\,
            lcout => \c0.n15_adj_4624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i147_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__69180\,
            in1 => \N__80416\,
            in2 => \N__79051\,
            in3 => \N__66242\,
            lcout => \c0.data_in_frame_18_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i149_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__80412\,
            in1 => \N__69181\,
            in2 => \N__66220\,
            in3 => \N__71953\,
            lcout => \c0.data_in_frame_18_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1535_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66666\,
            in1 => \N__66612\,
            in2 => \N__66521\,
            in3 => \N__66593\,
            lcout => \c0.n15_adj_4569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i152_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__80413\,
            in1 => \N__69182\,
            in2 => \N__76325\,
            in3 => \N__66552\,
            lcout => \c0.data_in_frame_18_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i182_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__66517\,
            in1 => \N__79758\,
            in2 => \_gnd_net_\,
            in3 => \N__78891\,
            lcout => data_in_frame_22_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i187_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__80414\,
            in1 => \N__78994\,
            in2 => \N__80986\,
            in3 => \N__77266\,
            lcout => \c0.data_in_frame_23_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i181_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__71943\,
            in1 => \N__75558\,
            in2 => \_gnd_net_\,
            in3 => \N__78897\,
            lcout => data_in_frame_22_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1625_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__66495\,
            in1 => \N__71247\,
            in2 => \_gnd_net_\,
            in3 => \N__66465\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4623_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1627_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77573\,
            in1 => \N__72489\,
            in2 => \N__66444\,
            in3 => \N__66441\,
            lcout => \c0.n13963\,
            ltout => \c0.n13963_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1563_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66435\,
            in1 => \N__66756\,
            in2 => \N__66396\,
            in3 => \N__66392\,
            lcout => \c0.n40_adj_4342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1526_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__68262\,
            in1 => \N__67151\,
            in2 => \_gnd_net_\,
            in3 => \N__75962\,
            lcout => \c0.n22495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i162_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__79983\,
            in1 => \N__80397\,
            in2 => \N__75229\,
            in3 => \N__67070\,
            lcout => \c0.data_in_frame_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_2_lut_adj_1379_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67055\,
            in2 => \_gnd_net_\,
            in3 => \N__67037\,
            lcout => \c0.n28_adj_4363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1483_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77150\,
            in1 => \N__66984\,
            in2 => \N__66957\,
            in3 => \N__66930\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1485_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__75946\,
            in2 => \N__66903\,
            in3 => \N__66898\,
            lcout => \c0.n24576\,
            ltout => \c0.n24576_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1471_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__66813\,
            in1 => \N__78025\,
            in2 => \N__66771\,
            in3 => \N__66687\,
            lcout => \c0.n14_adj_4519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1703_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__66752\,
            in1 => \_gnd_net_\,
            in2 => \N__75857\,
            in3 => \N__66714\,
            lcout => \c0.n22686\,
            ltout => \c0.n22686_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1432_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70575\,
            in1 => \N__66681\,
            in2 => \N__66669\,
            in3 => \N__78024\,
            lcout => \c0.n37_adj_4473\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i198_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__72991\,
            in1 => \N__79703\,
            in2 => \N__74870\,
            in3 => \N__79489\,
            lcout => \c0.data_in_frame_24_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1737_LC_23_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67552\,
            in1 => \N__67255\,
            in2 => \N__77394\,
            in3 => \N__67501\,
            lcout => OPEN,
            ltout => \c0.n30_adj_4489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67328\,
            in1 => \N__67461\,
            in2 => \N__67455\,
            in3 => \N__67452\,
            lcout => OPEN,
            ltout => \c0.n45_adj_4490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_adj_1456_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67335\,
            in1 => \N__67793\,
            in2 => \N__67446\,
            in3 => \N__67386\,
            lcout => OPEN,
            ltout => \c0.n48_adj_4503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_1459_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67443\,
            in1 => \N__67434\,
            in2 => \N__67422\,
            in3 => \N__67419\,
            lcout => \c0.n24573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_3_lut_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__78020\,
            in1 => \N__77956\,
            in2 => \_gnd_net_\,
            in3 => \N__67820\,
            lcout => \c0.n41_adj_4488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_1552_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67380\,
            in2 => \_gnd_net_\,
            in3 => \N__67361\,
            lcout => \c0.n27_adj_4502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1740_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67551\,
            in1 => \N__77391\,
            in2 => \N__67329\,
            in3 => \N__67256\,
            lcout => \c0.n21_adj_4481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1930_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__73899\,
            in1 => \N__67212\,
            in2 => \N__77189\,
            in3 => \N__67193\,
            lcout => \c0.n23_adj_4582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i219_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__76693\,
            in1 => \N__67862\,
            in2 => \N__79191\,
            in3 => \N__79476\,
            lcout => \c0.data_in_frame_27_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_3_lut_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__67824\,
            in1 => \N__67792\,
            in2 => \_gnd_net_\,
            in3 => \N__67773\,
            lcout => OPEN,
            ltout => \c0.n44_adj_4471_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_adj_1434_LC_23_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67767\,
            in1 => \N__67761\,
            in2 => \N__67752\,
            in3 => \N__67749\,
            lcout => OPEN,
            ltout => \c0.n24362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1490_LC_23_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111001"
        )
    port map (
            in0 => \N__67725\,
            in1 => \N__67716\,
            in2 => \N__67695\,
            in3 => \N__67692\,
            lcout => \c0.n26_adj_4530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i176_LC_23_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__77187\,
            in1 => \N__76274\,
            in2 => \_gnd_net_\,
            in3 => \N__67665\,
            lcout => data_in_frame_21_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1517_LC_23_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__73751\,
            in2 => \_gnd_net_\,
            in3 => \N__75732\,
            lcout => \c0.n22632\,
            ltout => \c0.n22632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1525_LC_23_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__73900\,
            in2 => \N__67566\,
            in3 => \N__81006\,
            lcout => \c0.n20358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1479_LC_23_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__68278\,
            in1 => \N__67563\,
            in2 => \_gnd_net_\,
            in3 => \N__75951\,
            lcout => OPEN,
            ltout => \c0.n22362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1488_LC_23_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68228\,
            in1 => \N__68370\,
            in2 => \N__68319\,
            in3 => \N__68316\,
            lcout => \c0.n13_adj_4527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1449_LC_23_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68279\,
            in1 => \N__77351\,
            in2 => \N__68241\,
            in3 => \N__68261\,
            lcout => \c0.n12_adj_4491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i231_LC_23_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__79471\,
            in1 => \N__68240\,
            in2 => \N__80080\,
            in3 => \N__73330\,
            lcout => \c0.data_in_frame_28_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i229_LC_23_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__80031\,
            in1 => \N__68229\,
            in2 => \N__71970\,
            in3 => \N__79472\,
            lcout => \c0.data_in_frame_28_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1870_LC_24_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69491\,
            in1 => \N__68923\,
            in2 => \N__68216\,
            in3 => \N__68646\,
            lcout => \c0.n28_adj_4286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i41_LC_24_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__80748\,
            in1 => \N__69460\,
            in2 => \_gnd_net_\,
            in3 => \N__68163\,
            lcout => data_in_frame_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_3_lut_4_lut_LC_24_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68145\,
            in1 => \N__68122\,
            in2 => \N__68040\,
            in3 => \N__68847\,
            lcout => \c0.n42_adj_4746\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i58_LC_24_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__75261\,
            in1 => \N__80843\,
            in2 => \N__67984\,
            in3 => \N__70187\,
            lcout => \c0.data_in_frame_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_2_lut_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68901\,
            in2 => \_gnd_net_\,
            in3 => \N__67934\,
            lcout => \c0.n24_adj_4213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1802_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68957\,
            in2 => \_gnd_net_\,
            in3 => \N__68669\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4687_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1803_LC_24_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68793\,
            in1 => \N__68728\,
            in2 => \N__68931\,
            in3 => \N__68844\,
            lcout => \c0.n23274\,
            ltout => \c0.n23274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1319_LC_24_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68900\,
            in1 => \N__69500\,
            in2 => \N__68892\,
            in3 => \N__68622\,
            lcout => \c0.n20_adj_4316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_3_lut_adj_1721_LC_24_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__68624\,
            in1 => \_gnd_net_\,
            in2 => \N__69504\,
            in3 => \N__68571\,
            lcout => \c0.n29_adj_4287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_4_lut_adj_1695_LC_24_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68845\,
            in1 => \N__68794\,
            in2 => \N__68749\,
            in3 => \N__68670\,
            lcout => \c0.n23276\,
            ltout => \c0.n23276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1183_LC_24_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__68623\,
            in1 => \_gnd_net_\,
            in2 => \N__68607\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_24_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__68600\,
            in1 => \N__68570\,
            in2 => \N__68559\,
            in3 => \N__68544\,
            lcout => \c0.n23343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i54_LC_24_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__79622\,
            in1 => \N__68395\,
            in2 => \_gnd_net_\,
            in3 => \N__69264\,
            lcout => data_in_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1302_LC_24_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72528\,
            in2 => \_gnd_net_\,
            in3 => \N__69547\,
            lcout => \c0.n22701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1804_LC_24_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69262\,
            in2 => \_gnd_net_\,
            in3 => \N__71117\,
            lcout => \c0.n5_adj_4323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i42_LC_24_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__69450\,
            in1 => \N__75251\,
            in2 => \_gnd_net_\,
            in3 => \N__70284\,
            lcout => data_in_frame_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_89_i9_2_lut_3_lut_LC_24_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__74358\,
            in1 => \N__74631\,
            in2 => \_gnd_net_\,
            in3 => \N__74500\,
            lcout => \c0.n9\,
            ltout => \c0.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i145_LC_24_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__80696\,
            in1 => \N__80427\,
            in2 => \N__69387\,
            in3 => \N__69275\,
            lcout => \c0.data_in_frame_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1617_LC_24_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69376\,
            in1 => \N__69329\,
            in2 => \N__69276\,
            in3 => \N__69263\,
            lcout => \c0.n19_adj_4620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i18_LC_24_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__69068\,
            in1 => \N__75252\,
            in2 => \N__70087\,
            in3 => \N__72529\,
            lcout => \c0.data_in_frame_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i61_LC_24_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__70193\,
            in1 => \N__80944\,
            in2 => \N__70347\,
            in3 => \N__71902\,
            lcout => \c0.data_in_frame_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1203_LC_24_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69825\,
            in2 => \_gnd_net_\,
            in3 => \N__69792\,
            lcout => \c0.n22392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i78_LC_24_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__70425\,
            in1 => \N__73703\,
            in2 => \N__79649\,
            in3 => \N__74117\,
            lcout => \c0.data_in_frame_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_13_i3_2_lut_LC_24_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__70401\,
            in2 => \_gnd_net_\,
            in3 => \N__71529\,
            lcout => \c0.n3_adj_4410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_2_lut_3_lut_LC_24_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__69860\,
            in1 => \N__70328\,
            in2 => \_gnd_net_\,
            in3 => \N__70264\,
            lcout => \c0.n40_adj_4288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i60_LC_24_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__80943\,
            in1 => \N__70194\,
            in2 => \N__77132\,
            in3 => \N__69861\,
            lcout => \c0.data_in_frame_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i97_LC_24_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__80718\,
            in1 => \N__79948\,
            in2 => \N__69833\,
            in3 => \N__73704\,
            lcout => \c0.data_in_frame_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i98_LC_24_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__73702\,
            in1 => \N__75257\,
            in2 => \N__80009\,
            in3 => \N__69793\,
            lcout => \c0.data_in_frame_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_2020_LC_24_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70683\,
            in1 => \N__69761\,
            in2 => \N__70971\,
            in3 => \N__69702\,
            lcout => \c0.n13253\,
            ltout => \c0.n13253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1624_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__69648\,
            in3 => \N__69644\,
            lcout => \c0.n22828\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_2018_LC_24_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70788\,
            in1 => \N__70749\,
            in2 => \N__70716\,
            in3 => \N__70701\,
            lcout => \c0.n27_adj_4748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i92_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__73690\,
            in1 => \N__76530\,
            in2 => \N__70673\,
            in3 => \N__77091\,
            lcout => \c0.data_in_frame_11_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1178_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__70850\,
            in2 => \_gnd_net_\,
            in3 => \N__70619\,
            lcout => \c0.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i159_LC_24_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__80399\,
            in1 => \N__76529\,
            in2 => \N__77649\,
            in3 => \N__73276\,
            lcout => \c0.data_in_frame_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i228_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__79491\,
            in1 => \N__79952\,
            in2 => \N__70571\,
            in3 => \N__77090\,
            lcout => \c0.data_in_frame_28_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i126_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__73689\,
            in1 => \N__80942\,
            in2 => \N__71246\,
            in3 => \N__79702\,
            lcout => \c0.data_in_frame_15_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i100_LC_24_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__77092\,
            in1 => \N__73691\,
            in2 => \N__70550\,
            in3 => \N__79947\,
            lcout => \c0.data_in_frame_12_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1727_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__70505\,
            in2 => \_gnd_net_\,
            in3 => \N__71674\,
            lcout => \c0.n22379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1514_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__73055\,
            in2 => \_gnd_net_\,
            in3 => \N__71269\,
            lcout => \c0.n6_adj_4559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i143_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__74116\,
            in1 => \N__80385\,
            in2 => \N__73307\,
            in3 => \N__71270\,
            lcout => \c0.data_in_frame_17_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1715_LC_24_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__71242\,
            in1 => \N__72195\,
            in2 => \_gnd_net_\,
            in3 => \N__71673\,
            lcout => \c0.n22605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_2016_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__71219\,
            in1 => \N__71175\,
            in2 => \N__71148\,
            in3 => \N__71126\,
            lcout => \c0.n30_adj_4747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1634_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__70959\,
            in1 => \N__70932\,
            in2 => \N__72464\,
            in3 => \N__70922\,
            lcout => \c0.n25_adj_4633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i76_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__74157\,
            in1 => \N__73687\,
            in2 => \N__77133\,
            in3 => \N__70876\,
            lcout => \c0.data_in_frame_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i91_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__73686\,
            in1 => \N__76525\,
            in2 => \N__79184\,
            in3 => \N__70849\,
            lcout => \c0.data_in_frame_11_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i226_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__79490\,
            in1 => \N__75178\,
            in2 => \N__70808\,
            in3 => \N__80008\,
            lcout => \c0.data_in_frame_28_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i108_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__75399\,
            in1 => \N__77124\,
            in2 => \N__72215\,
            in3 => \N__75507\,
            lcout => \c0.data_in_frame_13_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1236_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__77440\,
            in2 => \_gnd_net_\,
            in3 => \N__77405\,
            lcout => \c0.n14081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i107_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__75398\,
            in1 => \N__75506\,
            in2 => \N__79183\,
            in3 => \N__72463\,
            lcout => \c0.data_in_frame_13_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_4_lut_adj_2033_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72152\,
            in1 => \N__72252\,
            in2 => \N__72214\,
            in3 => \N__72318\,
            lcout => \c0.n16_adj_4627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1685_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__72251\,
            in1 => \N__72206\,
            in2 => \_gnd_net_\,
            in3 => \N__72153\,
            lcout => \c0.n4_adj_4586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1238_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72111\,
            in1 => \N__72090\,
            in2 => \N__72060\,
            in3 => \N__72032\,
            lcout => \c0.n10_adj_4250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i133_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__72938\,
            in1 => \N__80431\,
            in2 => \N__71946\,
            in3 => \N__71988\,
            lcout => \c0.data_in_frame_16_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i109_LC_24_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__75500\,
            in1 => \N__75415\,
            in2 => \N__71679\,
            in3 => \N__71906\,
            lcout => \c0.data_in_frame_13_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1709_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__73081\,
            in2 => \_gnd_net_\,
            in3 => \N__71627\,
            lcout => \c0.n16_adj_4666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_367_Select_18_i3_2_lut_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__71589\,
            in2 => \_gnd_net_\,
            in3 => \N__71544\,
            lcout => \c0.n3_adj_4400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i178_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__75177\,
            in2 => \N__73083\,
            in3 => \N__78890\,
            lcout => data_in_frame_22_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i121_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__80973\,
            in1 => \N__73706\,
            in2 => \N__73396\,
            in3 => \N__80719\,
            lcout => \c0.data_in_frame_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i191_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__73300\,
            in1 => \N__80323\,
            in2 => \N__75830\,
            in3 => \N__80974\,
            lcout => \c0.data_in_frame_23_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1378_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__75566\,
            in1 => \N__73734\,
            in2 => \N__73082\,
            in3 => \N__75823\,
            lcout => \c0.n29_adj_4362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i163_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__80007\,
            in1 => \N__80322\,
            in2 => \N__73059\,
            in3 => \N__79148\,
            lcout => \c0.data_in_frame_20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i190_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__80320\,
            in1 => \N__80975\,
            in2 => \N__79756\,
            in3 => \N__73020\,
            lcout => \c0.data_in_frame_23_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i136_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__72939\,
            in1 => \N__80321\,
            in2 => \N__72682\,
            in3 => \N__76293\,
            lcout => \c0.data_in_frame_16_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1616_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__72642\,
            in1 => \N__72612\,
            in2 => \N__72606\,
            in3 => \N__72587\,
            lcout => \c0.n22288\,
            ltout => \c0.n22288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1862_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72472\,
            in2 => \N__72417\,
            in3 => \N__72413\,
            lcout => \c0.n14160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i138_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__80401\,
            in1 => \N__74156\,
            in2 => \N__74712\,
            in3 => \N__75047\,
            lcout => \c0.data_in_frame_17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1998_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__74678\,
            in1 => \N__74524\,
            in2 => \N__74388\,
            in3 => \N__80400\,
            lcout => n22110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i202_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__74206\,
            in1 => \N__75046\,
            in2 => \N__73939\,
            in3 => \N__79481\,
            lcout => \c0.data_in_frame_25_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i161_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__80095\,
            in1 => \N__80617\,
            in2 => \N__73901\,
            in3 => \N__80403\,
            lcout => \c0.data_in_frame_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i153_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76683\,
            in1 => \N__80402\,
            in2 => \N__73863\,
            in3 => \N__80618\,
            lcout => \c0.data_in_frame_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1528_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__75614\,
            in1 => \N__74772\,
            in2 => \N__75562\,
            in3 => \N__75708\,
            lcout => \c0.n12_adj_4564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1726_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__75785\,
            in1 => \N__73796\,
            in2 => \_gnd_net_\,
            in3 => \N__75729\,
            lcout => \c0.n6_adj_4462\,
            ltout => \c0.n6_adj_4462_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_2_lut_3_lut_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__75548\,
            in2 => \N__73776\,
            in3 => \N__75612\,
            lcout => \c0.n22562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_rep_362_2_lut_3_lut_LC_24_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__74773\,
            in1 => \_gnd_net_\,
            in2 => \N__73752\,
            in3 => \N__75731\,
            lcout => \c0.n25484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__75549\,
            in1 => \N__75613\,
            in2 => \N__75996\,
            in3 => \N__76726\,
            lcout => \c0.n22769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1428_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__75947\,
            in1 => \N__75873\,
            in2 => \N__75858\,
            in3 => \N__75810\,
            lcout => \c0.n14_adj_4465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1389_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__75786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__75730\,
            lcout => \c0.n4_adj_4369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_3_lut_4_lut_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__74768\,
            in1 => \N__75553\,
            in2 => \N__75701\,
            in3 => \N__75620\,
            lcout => \c0.n73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_2_lut_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__75621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__75554\,
            lcout => \c0.n62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i106_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__75492\,
            in1 => \N__75416\,
            in2 => \N__75228\,
            in3 => \N__74933\,
            lcout => \c0.data_in_frame_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1592_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77392\,
            in1 => \N__74903\,
            in2 => \N__74866\,
            in3 => \N__74841\,
            lcout => \c0.n6718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1714_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__81002\,
            in1 => \N__77298\,
            in2 => \N__74774\,
            in3 => \N__74745\,
            lcout => \c0.n20239\,
            ltout => \c0.n20239_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1423_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77393\,
            in1 => \N__79226\,
            in2 => \N__77355\,
            in3 => \N__77352\,
            lcout => \c0.n10_adj_4457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1773_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__77188\,
            in1 => \N__77726\,
            in2 => \_gnd_net_\,
            in3 => \N__77217\,
            lcout => \c0.n6_adj_4668\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1560_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__77280\,
            in2 => \_gnd_net_\,
            in3 => \N__76797\,
            lcout => \c0.n13314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1774_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__77216\,
            in1 => \N__77180\,
            in2 => \_gnd_net_\,
            in3 => \N__77638\,
            lcout => \c0.n20350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i188_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__80987\,
            in1 => \N__77058\,
            in2 => \N__76815\,
            in3 => \N__80433\,
            lcout => \c0.data_in_frame_23_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1444_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__76776\,
            in1 => \N__76767\,
            in2 => \N__76758\,
            in3 => \N__76741\,
            lcout => \c0.n30_adj_4482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i160_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__76582\,
            in1 => \N__80432\,
            in2 => \N__77569\,
            in3 => \N__76394\,
            lcout => \c0.data_in_frame_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_adj_1647_LC_26_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__76086\,
            in2 => \_gnd_net_\,
            in3 => \N__76053\,
            lcout => \c0.n19_adj_4595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_LC_26_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__77883\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__77817\,
            lcout => \c0.n18\,
            ltout => \c0.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1710_LC_26_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__81103\,
            in1 => \N__77501\,
            in2 => \N__77754\,
            in3 => \N__77489\,
            lcout => \c0.n28_adj_4667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_4_lut_LC_26_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77453\,
            in1 => \N__77508\,
            in2 => \N__77655\,
            in3 => \N__77417\,
            lcout => OPEN,
            ltout => \c0.n24_adj_4653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1712_LC_26_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77751\,
            in1 => \N__77739\,
            in2 => \N__77733\,
            in3 => \N__81071\,
            lcout => \c0.n22369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_1650_LC_26_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__77709\,
            in2 => \_gnd_net_\,
            in3 => \N__77687\,
            lcout => \c0.n17_adj_4626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1669_LC_26_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__77650\,
            in1 => \N__77574\,
            in2 => \_gnd_net_\,
            in3 => \N__77517\,
            lcout => \c0.n15_adj_4625\,
            ltout => \c0.n15_adj_4625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1628_LC_26_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__77502\,
            in1 => \N__77490\,
            in2 => \N__77466\,
            in3 => \N__77463\,
            lcout => \c0.n24_adj_4628\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1692_LC_26_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__78841\,
            in1 => \N__77457\,
            in2 => \_gnd_net_\,
            in3 => \N__77421\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4629_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1629_LC_26_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__81104\,
            in1 => \N__81081\,
            in2 => \N__81075\,
            in3 => \N__81072\,
            lcout => \c0.n22234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i185_LC_26_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__80918\,
            in1 => \N__80729\,
            in2 => \N__80131\,
            in3 => \N__80430\,
            lcout => \c0.data_in_frame_23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i230_LC_26_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__80051\,
            in1 => \N__79757\,
            in2 => \N__79227\,
            in3 => \N__79488\,
            lcout => \c0.data_in_frame_28_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i179_LC_26_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__79192\,
            in1 => \N__78842\,
            in2 => \_gnd_net_\,
            in3 => \N__78911\,
            lcout => data_in_frame_22_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__78811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_1491_LC_26_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__78027\,
            in2 => \_gnd_net_\,
            in3 => \N__77954\,
            lcout => \c0.n24_adj_4531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
