-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Aug 25 2019 21:15:49

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : out std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : in std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : out std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__20080\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \VCCG0\ : std_logic;
signal \PIN_2_c\ : std_logic;
signal \c0.rx.r_Rx_Data_RZ0\ : std_logic;
signal \bfn_5_22_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_i_1\ : std_logic;
signal \c0.tx.r_Clock_Count12_cry_0\ : std_logic;
signal \c0.tx.r_Clock_Count_i_2\ : std_logic;
signal \c0.tx.r_Clock_Count12_cry_1\ : std_logic;
signal \c0.tx.r_Clock_Count_i_3\ : std_logic;
signal \c0.tx.r_Clock_Count12_cry_2\ : std_logic;
signal \c0.tx.r_Clock_Count12\ : std_logic;
signal \c0.tx.r_Clock_Count_i_0\ : std_logic;
signal \c0.rx.r_Rx_Bytece_0_4_cascade_\ : std_logic;
signal \c0.rx.N_336_cascade_\ : std_logic;
signal \c0.rx.r_Rx_Bytece_0_1\ : std_logic;
signal \c0.rx.r_SM_Main_RNI58REZ0Z_0_cascade_\ : std_logic;
signal \c0.rx.rx_data_ready\ : std_logic;
signal \blink_counterZ0Z_0\ : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal \blink_counterZ0Z_1\ : std_logic;
signal blink_counter_cry_0 : std_logic;
signal \blink_counterZ0Z_2\ : std_logic;
signal blink_counter_cry_1 : std_logic;
signal \blink_counterZ0Z_3\ : std_logic;
signal blink_counter_cry_2 : std_logic;
signal \blink_counterZ0Z_4\ : std_logic;
signal blink_counter_cry_3 : std_logic;
signal \blink_counterZ0Z_5\ : std_logic;
signal blink_counter_cry_4 : std_logic;
signal \blink_counterZ0Z_6\ : std_logic;
signal blink_counter_cry_5 : std_logic;
signal \blink_counterZ0Z_7\ : std_logic;
signal blink_counter_cry_6 : std_logic;
signal blink_counter_cry_7 : std_logic;
signal \blink_counterZ0Z_8\ : std_logic;
signal \bfn_6_22_0_\ : std_logic;
signal \blink_counterZ0Z_9\ : std_logic;
signal blink_counter_cry_8 : std_logic;
signal \blink_counterZ0Z_10\ : std_logic;
signal blink_counter_cry_9 : std_logic;
signal \blink_counterZ0Z_11\ : std_logic;
signal blink_counter_cry_10 : std_logic;
signal \blink_counterZ0Z_12\ : std_logic;
signal blink_counter_cry_11 : std_logic;
signal \blink_counterZ0Z_13\ : std_logic;
signal blink_counter_cry_12 : std_logic;
signal \blink_counterZ0Z_14\ : std_logic;
signal blink_counter_cry_13 : std_logic;
signal \blink_counterZ0Z_15\ : std_logic;
signal blink_counter_cry_14 : std_logic;
signal blink_counter_cry_15 : std_logic;
signal \blink_counterZ0Z_16\ : std_logic;
signal \bfn_6_23_0_\ : std_logic;
signal \blink_counterZ0Z_17\ : std_logic;
signal blink_counter_cry_16 : std_logic;
signal \blink_counterZ0Z_18\ : std_logic;
signal blink_counter_cry_17 : std_logic;
signal \blink_counterZ0Z_19\ : std_logic;
signal blink_counter_cry_18 : std_logic;
signal \blink_counterZ0Z_20\ : std_logic;
signal blink_counter_cry_19 : std_logic;
signal blink_counter_cry_20 : std_logic;
signal blink_counter_cry_21 : std_logic;
signal blink_counter_cry_22 : std_logic;
signal blink_counter_cry_23 : std_logic;
signal \bfn_6_24_0_\ : std_logic;
signal blink_counter_cry_24 : std_logic;
signal \c0.rx.r_Rx_Bytece_0_2_cascade_\ : std_logic;
signal \c0.rx.N_325\ : std_logic;
signal \c0.rx.N_325_cascade_\ : std_logic;
signal \c0.rx.r_Rx_Bytece_0_5_cascade_\ : std_logic;
signal \c0.rx.N_388\ : std_logic;
signal \c0.rx.r_Rx_Bytece_0_6_cascade_\ : std_logic;
signal \c0.rx.r_Rx_Byte_1_sqmuxa\ : std_logic;
signal \c0.rx.r_Rx_Bytece_0_0\ : std_logic;
signal \c0.rx.r_Rx_Byte_1_sqmuxa_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_RNO_0_0_0\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \c0.rx.r_Clock_Count_RNO_0_0_1\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_cry_0\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_cry_1\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_cry_2\ : std_logic;
signal \c0.rx.r_Clock_Count_RNO_0Z0Z_4\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_cry_3\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_cry_4\ : std_logic;
signal \c0.rx.r_Clock_Count_RNO_0Z0Z_6\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_cry_5\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_cry_6\ : std_logic;
signal \c0.rx.r_Clock_Count_RNO_0Z0Z_7\ : std_logic;
signal \c0.rx.r_Clock_CountZ1Z_1\ : std_logic;
signal \c0.rx.r_Clock_CountZ1Z_0\ : std_logic;
signal \c0.rx.N_320_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_8_f0_0_o2_0_2_cascade_\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_2_sqmuxa_0_i\ : std_logic;
signal \c0.rx.r_Clock_Count_8_f0_0_o2_0_2\ : std_logic;
signal \c0.rx.r_Clock_Count_RNO_0_0_2\ : std_logic;
signal \c0.rx.N_332_cascade_\ : std_logic;
signal \c0.rx.r_Clock_CountZ1Z_2\ : std_logic;
signal \c0.rx.r_Clock_CountZ1Z_6\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_7\ : std_logic;
signal \c0.rx.r_Clock_CountZ1Z_4\ : std_logic;
signal \c0.rx.r_Clock_Count_RNO_0Z0Z_5\ : std_logic;
signal \c0.rx.r_Clock_CountZ1Z_5\ : std_logic;
signal \c0.rx.N_320\ : std_logic;
signal \c0.rx.N_317\ : std_logic;
signal \c0.rx.N_337\ : std_logic;
signal \c0.rx.N_383_cascade_\ : std_logic;
signal \c0.rx.N_138r_0_i_1_cascade_\ : std_logic;
signal \c0.rx.r_SM_MainZ0Z_0\ : std_logic;
signal \c0.rx.N_91_0_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_illegal_0\ : std_logic;
signal \c0.rx.r_SM_Main_ns_0_i_a2_0_3_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_ns_0_i_a2_1_0_2\ : std_logic;
signal \c0.rx.r_SM_Main_dup_1\ : std_logic;
signal \c0.rx.un1_r_Rx_DV7_i_0_cascade_\ : std_logic;
signal \c0.rx.r_Rx_DV_RNOZ0Z_0\ : std_logic;
signal \c0.rx.r_SM_Main_dup_2\ : std_logic;
signal \c0.rx.r_SM_Main_ns_0_i_0_0_2\ : std_logic;
signal \c0.rx.r_Rx_DataZ0\ : std_logic;
signal \c0.rx.N_383\ : std_logic;
signal \c0.rx.N_321\ : std_logic;
signal \c0.rx.r_Clock_Count_8_f0_0_a2_0_0_2_cascade_\ : std_logic;
signal \c0.rx.N_371\ : std_logic;
signal \c0.rx.N_332\ : std_logic;
signal \c0.rx.r_SM_Main_RNI58REZ0Z_0\ : std_logic;
signal \c0.rx.N_361\ : std_logic;
signal \c0.rx.r_Clock_Count_RNO_0_0_3\ : std_logic;
signal \c0.rx.r_Clock_CountZ1Z_3\ : std_logic;
signal \c0.rx.N_386\ : std_logic;
signal \c0.rx.r_SM_Main_dup_3\ : std_logic;
signal \c0.rx.N_98_dup\ : std_logic;
signal \c0.rx.r_SM_Main_dup_4\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \c0.i12_0\ : std_logic;
signal \c0.i12_1\ : std_logic;
signal \c0.i12_2\ : std_logic;
signal \c0.i12_3\ : std_logic;
signal \c0.i12_4\ : std_logic;
signal \c0.i12_5\ : std_logic;
signal \c0.i12_7_and\ : std_logic;
signal \c0.i12_6\ : std_logic;
signal \c0.i12\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \c0.i12_0_and\ : std_logic;
signal \c0.i12_1_and\ : std_logic;
signal \blink_counterZ0Z_21\ : std_logic;
signal \blink_counterZ0Z_22\ : std_logic;
signal \blink_counterZ0Z_24\ : std_logic;
signal \N_12\ : std_logic;
signal \blink_counterZ0Z_25\ : std_logic;
signal \N_8_0_cascade_\ : std_logic;
signal \blink_counterZ0Z_23\ : std_logic;
signal \LED_c\ : std_logic;
signal \c0.tx.N_90_ip_RNIVJLQZ0_cascade_\ : std_logic;
signal \c0.tx.r_SM_Main_illegal_0\ : std_logic;
signal \c0.tx.N_90_dup_cascade_\ : std_logic;
signal \c0.tx.N_83_0\ : std_logic;
signal \c0.tx.r_Clock_Count_0_sqmuxa\ : std_logic;
signal \c0.tx.r_Clock_Count_RNO_0Z0Z_0\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_RNO_0Z0Z_1\ : std_logic;
signal \c0.tx.un1_r_Clock_Count_cry_0\ : std_logic;
signal \c0.tx.r_Clock_Count_RNO_0Z0Z_2\ : std_logic;
signal \c0.tx.un1_r_Clock_Count_cry_1\ : std_logic;
signal \c0.tx.un1_r_Clock_Count_cry_2\ : std_logic;
signal \c0.tx.r_Clock_Count_RNO_0Z0Z_3\ : std_logic;
signal \c0.tx.r_Clock_CountZ0Z_2\ : std_logic;
signal \c0.tx.r_Clock_CountZ0Z_1\ : std_logic;
signal \c0.tx.r_Clock_CountZ0Z_3\ : std_logic;
signal \c0.tx.r_Clock_CountZ0Z_0\ : std_logic;
signal \c0.tx.r_SM_Main_RNO_0Z0Z_1\ : std_logic;
signal \c0.tx.N_171_0_cascade_\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_8_cascade_\ : std_logic;
signal \c0.data_out_6_Z0Z_0\ : std_logic;
signal \c0.N_71\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \c0.dataZ0Z_1\ : std_logic;
signal \c0.data_cry_0\ : std_logic;
signal \c0.data_cry_1\ : std_logic;
signal \c0.dataZ0Z_3\ : std_logic;
signal \c0.data_cry_2\ : std_logic;
signal \c0.data_cry_3\ : std_logic;
signal \c0.dataZ0Z_5\ : std_logic;
signal \c0.data_cry_4\ : std_logic;
signal \c0.data_cry_5\ : std_logic;
signal \c0.dataZ0Z_7\ : std_logic;
signal \c0.data_cry_6\ : std_logic;
signal \c0.data_cry_7\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \c0.dataZ0Z_9\ : std_logic;
signal \c0.data_cry_8\ : std_logic;
signal \c0.dataZ0Z_10\ : std_logic;
signal \c0.data_cry_9\ : std_logic;
signal \c0.data_cry_10\ : std_logic;
signal \c0.data_cry_11\ : std_logic;
signal \c0.dataZ0Z_13\ : std_logic;
signal \c0.data_cry_12\ : std_logic;
signal \c0.data_cry_13\ : std_logic;
signal \c0.data_cry_14\ : std_logic;
signal \c0.i12_3_and\ : std_logic;
signal \c0.i12_6_and\ : std_logic;
signal \c0.i12_2_and\ : std_logic;
signal \c0.i12_5_and\ : std_logic;
signal \c0.i12_4_and\ : std_logic;
signal \c0.tx.r_Bit_Index_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \c0.tx.r_Tx_Active_1_sqmuxa_cascade_\ : std_logic;
signal \c0.tx.N_90_ip_RNIVJLQZ0\ : std_logic;
signal \c0.tx_active\ : std_logic;
signal \c0.tx.N_90_ip_RNI1U1EZ0_cascade_\ : std_logic;
signal \c0.tx.r_SM_Main_dup_4\ : std_logic;
signal \c0.tx_transmitZ0\ : std_logic;
signal \c0.tx.r_SM_Main_RNO_0Z0Z_0\ : std_logic;
signal \c0.tx.N_171_0\ : std_logic;
signal \c0.tx.r_SM_Main_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \c0.tx.r_SM_MainZ0Z_0\ : std_logic;
signal \c0.tx.N_90_dup\ : std_logic;
signal \c0.tx.r_Clock_Count12_THRU_CO\ : std_logic;
signal \c0.tx.r_SM_Main_RNIVDI71Z0Z_2\ : std_logic;
signal \c0.nextCRC16_3_0_a2_6_0_15\ : std_logic;
signal \c0.nextCRC16_3_9_cascade_\ : std_logic;
signal \c0.N_106_cascade_\ : std_logic;
signal \c0.N_92\ : std_logic;
signal \c0.N_106\ : std_logic;
signal \c0.data_out_7_Z0Z_0\ : std_logic;
signal \c0.nextCRC16_3_0_a2_0_10\ : std_logic;
signal \c0.dataZ0Z_12\ : std_logic;
signal \c0.N_77\ : std_logic;
signal \c0.N_76\ : std_logic;
signal \c0.dataZ0Z_0\ : std_logic;
signal \c0.dataZ0Z_14\ : std_logic;
signal \c0.dataZ0Z_11\ : std_logic;
signal \c0.dataZ0Z_2\ : std_logic;
signal \c0.dataZ0Z_15\ : std_logic;
signal \c0.dataZ0Z_4\ : std_logic;
signal \c0.dataZ0Z_8\ : std_logic;
signal \c0.data_in_0_Z0Z_4\ : std_logic;
signal \c0.data_in_1_Z0Z_0\ : std_logic;
signal \c0.rx_data_3\ : std_logic;
signal \c0.rx_data_1\ : std_logic;
signal \c0.rx_data_0\ : std_logic;
signal \c0.tx.o_Tx_Serial_2_3_i_m2_ns_1_cascade_\ : std_logic;
signal \c0.tx.N_90_ip_RNI1U1EZ0\ : std_logic;
signal \c0.tx.o_Tx_Serial_2_6_i_m2_ns_1_cascade_\ : std_logic;
signal \c0.tx.o_Tx_Serial_RNO_3_0\ : std_logic;
signal \c0.tx.o_Tx_Serial_RNO_2_0_cascade_\ : std_logic;
signal \c0.tx.r_SM_Main_RNI522EZ0Z_4\ : std_logic;
signal \c0.tx.o_Tx_Serial_RNOZ0Z_1_cascade_\ : std_logic;
signal \c0.tx.r_SM_Main_dup_3\ : std_logic;
signal \PIN_1_c\ : std_logic;
signal \c0.tx.N_390_i\ : std_logic;
signal \c0.tx.r_SM_Main_dup_2\ : std_logic;
signal \c0.tx.r_SM_Main_recr_i_0_a2_0_2_0_1_3\ : std_logic;
signal \c0.tx.r_Bit_IndexZ0Z_1\ : std_logic;
signal \c0.tx.r_Bit_IndexZ0Z_2\ : std_logic;
signal \c0.tx.r_SM_Main_dup_1\ : std_logic;
signal \c0.tx.r_Bit_IndexZ0Z_0\ : std_logic;
signal \c0.tx.r_SM_Main_recr_i_i_a2_0_1_2\ : std_logic;
signal \c0.data_out_7_Z0Z_5\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_3_cascade_\ : std_logic;
signal \c0.d_2_19\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_3\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_2_cascade_\ : std_logic;
signal \c0.dataZ0Z_6\ : std_logic;
signal \c0.N_99_cascade_\ : std_logic;
signal \c0.nextCRC16_3_0_a2_0_0\ : std_logic;
signal \c0.nextCRC16_3_0_a2_3_0_cascade_\ : std_logic;
signal \c0.nextCRC16_3_0_a2_4_0\ : std_logic;
signal \c0.d_2_27\ : std_logic;
signal \c0.N_81_cascade_\ : std_logic;
signal \c0.N_105\ : std_logic;
signal \c0.N_105_cascade_\ : std_logic;
signal \c0.data_out_6_Z0Z_5\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_15_cascade_\ : std_logic;
signal \c0.N_99\ : std_logic;
signal \c0.nextCRC16_3_0_a2_5_15\ : std_logic;
signal \c0.nextCRC16_3_0_a2_2_15\ : std_logic;
signal \c0.N_95_cascade_\ : std_logic;
signal \c0.N_85\ : std_logic;
signal \c0.nextCRC16_3_2_1\ : std_logic;
signal \c0.d_2_3\ : std_logic;
signal \c0.N_75\ : std_logic;
signal \c0.N_75_cascade_\ : std_logic;
signal \c0.N_93\ : std_logic;
signal \c0.d_2_35\ : std_logic;
signal \c0.rx_data_7\ : std_logic;
signal \c0.data_in_2_Z0Z_5\ : std_logic;
signal \c0.data_in_2_Z0Z_3\ : std_logic;
signal \c0.data_in_0_Z0Z_7\ : std_logic;
signal \c0.data_in_2_Z0Z_7\ : std_logic;
signal \c0.data_in_6_Z0Z_0\ : std_logic;
signal \c0.data_in_2_Z0Z_4\ : std_logic;
signal \c0.data_in_4_Z0Z_2\ : std_logic;
signal \c0.data_in_4_Z0Z_5\ : std_logic;
signal \c0.data_in_0_Z0Z_0\ : std_logic;
signal \c0.data_in_1_Z0Z_3\ : std_logic;
signal \c0.data_in_1_Z0Z_7\ : std_logic;
signal \c0.data_in_3_Z0Z_0\ : std_logic;
signal \c0.data_in_3_Z0Z_5\ : std_logic;
signal \c0.data_in_4_Z0Z_1\ : std_logic;
signal \c0.data_in_4_Z0Z_7\ : std_logic;
signal \c0.data_in_5_Z0Z_3\ : std_logic;
signal \c0.N_108_cascade_\ : std_logic;
signal \c0.N_122_cascade_\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_2_cascade_\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_4_cascade_\ : std_logic;
signal \c0.data_in_7_Z0Z_3\ : std_logic;
signal \c0.data_in_2_Z0Z_1\ : std_logic;
signal \c0.data_in_3_Z0Z_6\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_3\ : std_logic;
signal \c0.data_in_6_Z0Z_3\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_3\ : std_logic;
signal \c0.d_4_17\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_1\ : std_logic;
signal \c0.m161_ns_1_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_1\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_2\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_2\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_2\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_3\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_3\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_3\ : std_logic;
signal \c0.d_2_7\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_7_cascade_\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_7\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_7_cascade_\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_7\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_4\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_5\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_5\ : std_logic;
signal \c0.N_24_0\ : std_logic;
signal \c0.un144_newcrc_2\ : std_logic;
signal \c0.un144_newcrc_5_cascade_\ : std_logic;
signal \c0.data_out_7_Z0Z_6\ : std_logic;
signal \c0.N_81\ : std_logic;
signal \c0.data_out_6_Z0Z_6\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_4_cascade_\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_4\ : std_logic;
signal \c0.d_2_20\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_4\ : std_logic;
signal \c0.N_95\ : std_logic;
signal \c0.d_2_8\ : std_logic;
signal \c0.d_2_0\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_0_cascade_\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_0\ : std_logic;
signal \c0.d_2_33\ : std_logic;
signal \c0.d_2_34\ : std_logic;
signal \c0.d_2_15\ : std_logic;
signal \c0.d_2_43\ : std_logic;
signal \c0.un105_newcrc_0_a2_0_cascade_\ : std_logic;
signal \c0.N_100\ : std_logic;
signal \c0.d_2_31\ : std_logic;
signal \c0.un105_newcrc_0_a2_3\ : std_logic;
signal \c0.d_2_32\ : std_logic;
signal \c0.d_2_24\ : std_logic;
signal \c0.nextCRC16_3_3_12\ : std_logic;
signal \c0.nextCRC16_3_4_12_cascade_\ : std_logic;
signal \c0.d_2_41\ : std_logic;
signal \c0.N_94\ : std_logic;
signal \c0.N_94_cascade_\ : std_logic;
signal \c0.d_2_23\ : std_logic;
signal \c0.d_2_40\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_11\ : std_logic;
signal \c0.data_out_6_Z0Z_4\ : std_logic;
signal \c0.data_out_7_Z0Z_4\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_4\ : std_logic;
signal \c0.data_in_5_Z0Z_5\ : std_logic;
signal \c0.rx_data_4\ : std_logic;
signal \c0.rx_data_2\ : std_logic;
signal \c0.d_4_34\ : std_logic;
signal \c0.un1_data_in_7__7_0_a2_0_a2_2_cascade_\ : std_logic;
signal \c0.un1_data_in_6__0_0_a2_5_a2_2\ : std_logic;
signal \c0.un1_data_in_7__7_i_cascade_\ : std_logic;
signal \c0.data_in_5_Z0Z_7\ : std_logic;
signal \c0.data_in_4_Z0Z_3\ : std_logic;
signal \c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_\ : std_logic;
signal \c0.data_in_3_Z0Z_4\ : std_logic;
signal \c0.data_in_1_Z0Z_5\ : std_logic;
signal \c0.data_in_3_Z0Z_2\ : std_logic;
signal \c0.data_in_5_Z0Z_1\ : std_logic;
signal \c0.data_in_5_Z0Z_0\ : std_logic;
signal \c0.N_132\ : std_logic;
signal \c0.un1_data_in_7__0_0_a2_1_a2_5_cascade_\ : std_logic;
signal \c0.N_121_cascade_\ : std_logic;
signal \c0.N_125\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_4_3_cascade_\ : std_logic;
signal \c0.N_136\ : std_logic;
signal \c0.N_136_cascade_\ : std_logic;
signal \c0.un1_data_in_7__0_0_a2_1_a2_2\ : std_logic;
signal \c0.data_in_3_Z0Z_3\ : std_logic;
signal \c0.un1_data_in_7__1_0_a2_24_a2_3_cascade_\ : std_logic;
signal \c0.un1_data_in_7__1_0_a2_24_a2_4\ : std_logic;
signal \c0.data_in_5_Z0Z_4\ : std_logic;
signal \c0.data_in_5_Z0Z_2\ : std_logic;
signal \c0.data_in_2_Z0Z_0\ : std_logic;
signal \c0.d_4_33\ : std_logic;
signal \c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_\ : std_logic;
signal \c0.N_124\ : std_logic;
signal \c0.N_124_cascade_\ : std_logic;
signal \c0.N_108\ : std_logic;
signal \c0.un1_data_in_7__6_0_a2_5_a2_2_cascade_\ : std_logic;
signal \c0.un1_data_in_7__4_0_a2_0_a2_4\ : std_logic;
signal \c0.data_in_0_Z0Z_3\ : std_logic;
signal \c0.data_in_0_Z0Z_5\ : std_logic;
signal \c0.data_in_2_Z0Z_2\ : std_logic;
signal \c0.d_4_18\ : std_logic;
signal \c0.d_2_38\ : std_logic;
signal \c0.d_2_46\ : std_logic;
signal \c0.data_out_6_Z0Z_7\ : std_logic;
signal \c0.data_out_7_Z0Z_7\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_7\ : std_logic;
signal \c0.d_2_37\ : std_logic;
signal \c0.d_2_45\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_5\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_6_cascade_\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_6\ : std_logic;
signal \c0.d_2_42\ : std_logic;
signal \c0.nextCRC16_3_3_1\ : std_logic;
signal \c0.d_2_4\ : std_logic;
signal \c0.nextCRC16_3_3_1_cascade_\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_1\ : std_logic;
signal \c0.d_2_28\ : std_logic;
signal \c0.d_2_5\ : std_logic;
signal \c0.d_2_13\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_5_cascade_\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_5\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_5\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_0\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_0\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_0\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_0\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_2\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_2\ : std_logic;
signal \c0.d_2_25\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_1_cascade_\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_1\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_1_cascade_\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_1\ : std_logic;
signal \c0.data_out_7_Z0Z_2\ : std_logic;
signal \c0.data_out_6_Z0Z_2\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_2\ : std_logic;
signal \c0.d_2_1\ : std_logic;
signal \c0.d_2_9\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_1\ : std_logic;
signal \c0.d_2_2\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_2_cascade_\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_2\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_2\ : std_logic;
signal \c0.d_2_39\ : std_logic;
signal \c0.d_2_47\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_7\ : std_logic;
signal \c0.d_2_36\ : std_logic;
signal \c0.d_2_44\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_4\ : std_logic;
signal \c0.data_out_6_Z0Z_1\ : std_logic;
signal \c0.data_out_7_Z0Z_1\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_1\ : std_logic;
signal \c0.m2_e_1_cascade_\ : std_logic;
signal \c0.data_out_7_Z0Z_3\ : std_logic;
signal \c0.data_out_6_Z0Z_3\ : std_logic;
signal \c0.N_132_mux_cascade_\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_3\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_5\ : std_logic;
signal \c0.data_in_6_Z0Z_7\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_7\ : std_logic;
signal \c0.data_in_7_Z0Z_7\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_7\ : std_logic;
signal \c0.data_in_0_Z0Z_6\ : std_logic;
signal \c0.d_4_6\ : std_logic;
signal \c0.N_109\ : std_logic;
signal \c0.data_in_1_Z0Z_6\ : std_logic;
signal \c0.d_4_7\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_7\ : std_logic;
signal \c0.data_in_4_Z0Z_4\ : std_logic;
signal \c0.data_in_6_Z0Z_1\ : std_logic;
signal \c0.N_34_cascade_\ : std_logic;
signal \c0.data_in_2_Z0Z_6\ : std_logic;
signal \c0.d_4_44\ : std_logic;
signal \c0.d_4_36\ : std_logic;
signal \c0.N_104\ : std_logic;
signal \c0.un1_data_in_6__3_0_a2_5_a2_2\ : std_logic;
signal \c0.un1_data_in_6__5_cascade_\ : std_logic;
signal \c0.un1_data_in_6__6\ : std_logic;
signal \c0.un1_data_in_6__1_0_a2_4_a2_2\ : std_logic;
signal \c0.m163_2_cascade_\ : std_logic;
signal \c0.N_126\ : std_logic;
signal \c0.m163_7_cascade_\ : std_logic;
signal \c0.m163_0\ : std_logic;
signal \c0.un1_data_in_6__5_0_a2_5_a2_2\ : std_logic;
signal \c0.N_120\ : std_logic;
signal \c0.data_in_1_Z0Z_4\ : std_logic;
signal \c0.N_121\ : std_logic;
signal \c0.m163_4\ : std_logic;
signal \c0.un1_data_in_7__1_0_a2_24_a2_7\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_6\ : std_logic;
signal \c0.m163_8_cascade_\ : std_logic;
signal \c0.un1_data_in_7__1_3\ : std_logic;
signal \c0.m163_10\ : std_logic;
signal \c0.m163_1_cascade_\ : std_logic;
signal \c0.un1_data_in_7__0\ : std_logic;
signal \c0.N_164_0_cascade_\ : std_logic;
signal \c0.N_173_0_cascade_\ : std_logic;
signal \c0.data_in_3_Z0Z_7\ : std_logic;
signal \c0.d_4_RNIB3JJZ0Z_2\ : std_logic;
signal \c0.data_in_0_Z0Z_2\ : std_logic;
signal \c0.data_in_4_Z0Z_0\ : std_logic;
signal \c0.d_4_23\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_7\ : std_logic;
signal \c0.d_4_2\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_2\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_2_cascade_\ : std_logic;
signal \c0.m131_ns_1\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_6\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_6\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_6\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_6\ : std_logic;
signal \c0.tx.N_398_i\ : std_logic;
signal \c0.rx.r_Bit_IndexZ0Z_1\ : std_logic;
signal \c0.rx.r_Bit_IndexZ0Z_2\ : std_logic;
signal \c0.rx.r_Bit_IndexZ0Z_0\ : std_logic;
signal \c0.rx.N_335\ : std_logic;
signal \c0.d_4_35\ : std_logic;
signal \c0.d_4_27\ : std_logic;
signal \c0.d_4_19\ : std_logic;
signal \c0.d_4_3\ : std_logic;
signal \c0.d_4_11\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_3\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_3_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_3\ : std_logic;
signal \c0.m105_ns_1_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_3\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_3\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_7\ : std_logic;
signal \c0.m60_0_ns_1\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_7\ : std_logic;
signal \c0.d_2_6\ : std_logic;
signal \c0.d_2_22\ : std_logic;
signal \c0.d_2_14\ : std_logic;
signal \c0.d_2_30\ : std_logic;
signal \c0.d_2_16\ : std_logic;
signal \c0.d_2_17\ : std_logic;
signal \c0.d_2_12\ : std_logic;
signal \c0.d_2_21\ : std_logic;
signal \c0.d_2_11\ : std_logic;
signal \c0.d_2_26\ : std_logic;
signal \c0.d_2_18\ : std_logic;
signal \c0.d_2_10\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_6\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_7\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_3\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_4\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_1\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_0\ : std_logic;
signal \c0.N_132_mux\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_2\ : std_logic;
signal \c0.N_5_1_cascade_\ : std_logic;
signal \c0.byte_transmit_counter15\ : std_logic;
signal \c0.data_out_0__1_sqmuxa\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_4\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_4\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_4\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_4\ : std_logic;
signal \c0.m120_ns_1_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_6\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_6\ : std_logic;
signal \c0.m90_ns_1_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_6\ : std_logic;
signal \c0.data_in_7_Z0Z_4\ : std_logic;
signal \c0.rx_data_5\ : std_logic;
signal \c0.data_in_4_Z0Z_6\ : std_logic;
signal \c0.data_in_5_Z0Z_6\ : std_logic;
signal \c0.rx_data_6\ : std_logic;
signal \c0.d_4_26\ : std_logic;
signal \c0.data_in_6_Z0Z_4\ : std_logic;
signal \c0.d_4_41\ : std_logic;
signal \c0.un1_data_in_6__4_0_a2_5_a2_1\ : std_logic;
signal \c0.data_in_1_Z0Z_2\ : std_logic;
signal \c0.d_4_10\ : std_logic;
signal \c0.N_127\ : std_logic;
signal \c0.data_in_1_Z0Z_1\ : std_logic;
signal \c0.data_in_3_Z0Z_1\ : std_logic;
signal \c0.d_4_25\ : std_logic;
signal \c0.d_4_38\ : std_logic;
signal \c0.N_107\ : std_logic;
signal \c0.un1_data_in_6__2_0_a2_6_a2_2_cascade_\ : std_logic;
signal \c0.un1_data_in_6__2\ : std_logic;
signal \c0.d_4_46\ : std_logic;
signal \c0.d_4_42\ : std_logic;
signal \c0.N_133\ : std_logic;
signal \c0.un1_data_in_7__2_0_a2_0_a2_5_cascade_\ : std_logic;
signal \c0.un1_data_in_7__2\ : std_logic;
signal \c0.d_4_14\ : std_logic;
signal \c0.d_4_31\ : std_logic;
signal \c0.un1_data_in_7__2_0_a2_0_a2_4\ : std_logic;
signal \c0.un1_data_in_7__3_0_a2_0_a2_3\ : std_logic;
signal \c0.d_4_43\ : std_logic;
signal \c0.N_128\ : std_logic;
signal \c0.un1_data_in_7__3_0_a2_0_a2_4_cascade_\ : std_logic;
signal \c0.un1_data_in_7__5_0_a2_0_a2_1\ : std_logic;
signal \c0.m163_9\ : std_logic;
signal \c0.data_in_0_Z0Z_1\ : std_logic;
signal \c0.N_123\ : std_logic;
signal \c0.d_4_15\ : std_logic;
signal \c0.N_129\ : std_logic;
signal \c0.N_18\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_cry_0\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_cry_1\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_cry_2\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_cry_3\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_cry_4\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_cry_5\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_cry_6\ : std_logic;
signal \c0.d_4_1\ : std_logic;
signal \c0.d_4_9\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_1\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_1\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_1\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_1\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_4\ : std_logic;
signal \c0.N_173_0\ : std_logic;
signal \c0.tx2.r_Clock_Count_i_0\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \c0.tx2.r_Clock_Count_i_1\ : std_logic;
signal \c0.tx2.r_Clock_Count12_cry_0\ : std_logic;
signal \c0.tx2.r_Clock_Count_i_2\ : std_logic;
signal \c0.tx2.r_Clock_Count12_cry_1\ : std_logic;
signal \c0.tx2.r_Clock_Count_i_3\ : std_logic;
signal \c0.tx2.r_Clock_Count12_cry_2\ : std_logic;
signal \c0.tx2.r_Clock_Count12\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \c0.d_2_29\ : std_logic;
signal \c0.data_out_0__1_sqmuxa_g\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_6\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_2\ : std_logic;
signal \c0.tx2.o_Tx_Serial_RNOZ0Z_6_cascade_\ : std_logic;
signal \c0.tx2.o_Tx_Serial_RNOZ0Z_5\ : std_logic;
signal \c0.tx2.o_Tx_Serial_RNOZ0Z_3\ : std_logic;
signal \c0.tx2.m195_ns_1_cascade_\ : std_logic;
signal \c0.tx2.o_Tx_Serial_RNOZ0Z_2\ : std_logic;
signal \c0.tx2.N_196_0_cascade_\ : std_logic;
signal \c0.tx2.N_493_cascade_\ : std_logic;
signal \c0.tx2.N_205_mux\ : std_logic;
signal \PIN_3_c\ : std_logic;
signal \c0.data_in_7_Z0Z_0\ : std_logic;
signal \c0.data_in_7_Z0Z_1\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_1\ : std_logic;
signal \c0.data_in_6_Z0Z_5\ : std_logic;
signal \c0.data_in_7_Z0Z_5\ : std_logic;
signal \c0.data_in_7_Z0Z_6\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_6\ : std_logic;
signal \c0.data_in_6_Z0Z_6\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_6\ : std_logic;
signal \c0.data_in_frame_0__0_sqmuxa_g\ : std_logic;
signal \c0.data_in_7_Z0Z_2\ : std_logic;
signal \c0.data_in_6_Z0Z_2\ : std_logic;
signal \c0.rx_data_ready_g\ : std_logic;
signal \c0.d_4_45\ : std_logic;
signal \c0.d_4_37\ : std_logic;
signal \c0.d_4_29\ : std_logic;
signal \c0.d_4_21\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_5_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_5\ : std_logic;
signal \c0.m75_ns_1_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_5\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_5\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_5\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_5\ : std_logic;
signal \c0.d_4_47\ : std_logic;
signal \c0.d_4_39\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_7\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_0\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_0\ : std_logic;
signal \c0.N_164_0\ : std_logic;
signal \c0.d_4_22\ : std_logic;
signal \c0.d_4_30\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_6\ : std_logic;
signal \c0.d_4_4\ : std_logic;
signal \c0.d_4_12\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_4\ : std_logic;
signal \c0.d_4_28\ : std_logic;
signal \c0.d_4_20\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_4\ : std_logic;
signal \c0.d_4_13\ : std_logic;
signal \c0.d_4_5\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_5\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_7\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_3\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_6\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_5\ : std_logic;
signal \c0.m45_0_0_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_4\ : std_logic;
signal \c0.N_204_mux_cascade_\ : std_logic;
signal \c0.N_215_mux\ : std_logic;
signal \c0.d_4_0\ : std_logic;
signal \c0.d_4_8\ : std_logic;
signal \c0.d_4_16\ : std_logic;
signal \c0.d_4_24\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_1\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_0\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_0_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_2\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_0\ : std_logic;
signal \c0.m146_ns_1_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_0\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_0\ : std_logic;
signal \c0.d_4_32\ : std_logic;
signal \c0.N_204_mux\ : std_logic;
signal \c0.d_4_40\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_0\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \c0.tx2.un1_r_Clock_Count_cry_0\ : std_logic;
signal \c0.tx2.un1_r_Clock_Count_cry_1\ : std_logic;
signal \c0.tx2.un1_r_Clock_Count_cry_2\ : std_logic;
signal \c0.tx2.r_Clock_CountZ0Z_2\ : std_logic;
signal \c0.tx2.r_Clock_CountZ0Z_1\ : std_logic;
signal \c0.tx2.r_Clock_CountZ0Z_3\ : std_logic;
signal \c0.tx2.r_Clock_CountZ0Z_0\ : std_logic;
signal \c0.tx2.N_16_0\ : std_logic;
signal \c0.tx2.r_Clock_Count_0_sqmuxa\ : std_logic;
signal \c0.tx2.N_83_0_cascade_\ : std_logic;
signal \c0.N_90_dup_cascade_\ : std_logic;
signal \c0.tx2.i97_mux_cascade_\ : std_logic;
signal \c0.tx2.r_SM_Main_illegal_0\ : std_logic;
signal \c0.tx2.N_214_0\ : std_logic;
signal \c0.tx2.r_Clock_Count12_THRU_CO\ : std_logic;
signal \c0.tx2.N_17_0_cascade_\ : std_logic;
signal \c0.tx2.r_SM_Main_dup_4\ : std_logic;
signal \c0.tx2.r_Bit_IndexZ1Z_0\ : std_logic;
signal \c0.tx2.N_212_0_cascade_\ : std_logic;
signal \c0.tx2.r_SM_Main_dup_1\ : std_logic;
signal \c0.tx2.N_496_cascade_\ : std_logic;
signal \c0.tx2.r_SM_Main_dup_2\ : std_logic;
signal \c0.tx2.N_171_0\ : std_logic;
signal \c0.tx2.N_17_0\ : std_logic;
signal \c0.tx2.N_212_0\ : std_logic;
signal \c0.tx2.N_493\ : std_logic;
signal \c0.tx2.r_SM_Main_dup_3\ : std_logic;
signal \c0.tx2_transmitZ0\ : std_logic;
signal \c0.N_19_0\ : std_logic;
signal \c0.r_SM_Main_0\ : std_logic;
signal \c0.N_90_dup\ : std_logic;
signal \c0.tx2.N_9_1_cascade_\ : std_logic;
signal \c0.tx2.r_Bit_IndexZ0Z_2\ : std_logic;
signal \c0.tx2.N_12_0\ : std_logic;
signal \c0.tx2.N_9_1\ : std_logic;
signal \c0.tx2.r_Bit_IndexZ0Z_1\ : std_logic;
signal \c0.tx2_active\ : std_logic;
signal \c0.N_170_0\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \c0.tx2_transmit_0_sqmuxa\ : std_logic;
signal \c0.wait_for_transmissionZ0\ : std_logic;
signal \c0.i12_THRU_CO\ : std_logic;
signal \c0.data_in_frame_0__0_sqmuxa\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \PIN_1_wire\ : std_logic;
signal \PIN_2_wire\ : std_logic;
signal \PIN_3_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    LED <= \LED_wire\;
    PIN_1 <= \PIN_1_wire\;
    \PIN_2_wire\ <= PIN_2;
    PIN_3 <= \PIN_3_wire\;
    USBPU <= \USBPU_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__20078\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20080\,
            DIN => \N__20079\,
            DOUT => \N__20078\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20080\,
            PADOUT => \N__20079\,
            PADIN => \N__20078\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20069\,
            DIN => \N__20068\,
            DOUT => \N__20067\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20069\,
            PADOUT => \N__20068\,
            PADIN => \N__20067\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__9190\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20060\,
            DIN => \N__20059\,
            DOUT => \N__20058\,
            PACKAGEPIN => \PIN_1_wire\
        );

    \PIN_1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20060\,
            PADOUT => \N__20059\,
            PADIN => \N__20058\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10288\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20051\,
            DIN => \N__20050\,
            DOUT => \N__20049\,
            PACKAGEPIN => \PIN_2_wire\
        );

    \PIN_2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20051\,
            PADOUT => \N__20050\,
            PADIN => \N__20049\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_2_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20042\,
            DIN => \N__20041\,
            DOUT => \N__20040\,
            PACKAGEPIN => \PIN_3_wire\
        );

    \PIN_3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20042\,
            PADOUT => \N__20041\,
            PADIN => \N__20040\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__17404\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20033\,
            DIN => \N__20032\,
            DOUT => \N__20031\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20033\,
            PADOUT => \N__20032\,
            PADIN => \N__20031\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__4707\ : InMux
    port map (
            O => \N__20014\,
            I => \N__20008\
        );

    \I__4706\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20005\
        );

    \I__4705\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20002\
        );

    \I__4704\ : InMux
    port map (
            O => \N__20011\,
            I => \N__19999\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__19996\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__20005\,
            I => \N__19993\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20002\,
            I => \N__19990\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__19999\,
            I => \N__19983\
        );

    \I__4699\ : Span4Mux_v
    port map (
            O => \N__19996\,
            I => \N__19983\
        );

    \I__4698\ : Span4Mux_h
    port map (
            O => \N__19993\,
            I => \N__19983\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__19990\,
            I => \c0.tx2_transmitZ0\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__19983\,
            I => \c0.tx2_transmitZ0\
        );

    \I__4695\ : CEMux
    port map (
            O => \N__19978\,
            I => \N__19974\
        );

    \I__4694\ : CEMux
    port map (
            O => \N__19977\,
            I => \N__19970\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19965\
        );

    \I__4692\ : CEMux
    port map (
            O => \N__19973\,
            I => \N__19962\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19959\
        );

    \I__4690\ : CEMux
    port map (
            O => \N__19969\,
            I => \N__19956\
        );

    \I__4689\ : CEMux
    port map (
            O => \N__19968\,
            I => \N__19953\
        );

    \I__4688\ : Span4Mux_v
    port map (
            O => \N__19965\,
            I => \N__19947\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__19962\,
            I => \N__19947\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__19959\,
            I => \N__19941\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__19956\,
            I => \N__19941\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__19953\,
            I => \N__19938\
        );

    \I__4683\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19935\
        );

    \I__4682\ : Span4Mux_h
    port map (
            O => \N__19947\,
            I => \N__19932\
        );

    \I__4681\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19929\
        );

    \I__4680\ : Span4Mux_v
    port map (
            O => \N__19941\,
            I => \N__19922\
        );

    \I__4679\ : Span4Mux_h
    port map (
            O => \N__19938\,
            I => \N__19922\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__19935\,
            I => \N__19922\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__19932\,
            I => \c0.N_19_0\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__19929\,
            I => \c0.N_19_0\
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__19922\,
            I => \c0.N_19_0\
        );

    \I__4674\ : CascadeMux
    port map (
            O => \N__19915\,
            I => \N__19909\
        );

    \I__4673\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19904\
        );

    \I__4672\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19904\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__19912\,
            I => \N__19900\
        );

    \I__4670\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19895\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19892\
        );

    \I__4668\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19883\
        );

    \I__4667\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19883\
        );

    \I__4666\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19883\
        );

    \I__4665\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19883\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__19895\,
            I => \c0.r_SM_Main_0\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__19892\,
            I => \c0.r_SM_Main_0\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__19883\,
            I => \c0.r_SM_Main_0\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__19876\,
            I => \N__19872\
        );

    \I__4660\ : InMux
    port map (
            O => \N__19875\,
            I => \N__19867\
        );

    \I__4659\ : InMux
    port map (
            O => \N__19872\,
            I => \N__19862\
        );

    \I__4658\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19862\
        );

    \I__4657\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19853\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__19867\,
            I => \N__19848\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__19862\,
            I => \N__19848\
        );

    \I__4654\ : InMux
    port map (
            O => \N__19861\,
            I => \N__19841\
        );

    \I__4653\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19841\
        );

    \I__4652\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19841\
        );

    \I__4651\ : InMux
    port map (
            O => \N__19858\,
            I => \N__19834\
        );

    \I__4650\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19834\
        );

    \I__4649\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19834\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__19853\,
            I => \c0.N_90_dup\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__19848\,
            I => \c0.N_90_dup\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__19841\,
            I => \c0.N_90_dup\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__19834\,
            I => \c0.N_90_dup\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__19825\,
            I => \c0.tx2.N_9_1_cascade_\
        );

    \I__4643\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19819\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__19819\,
            I => \N__19812\
        );

    \I__4641\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19806\
        );

    \I__4640\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19806\
        );

    \I__4639\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19803\
        );

    \I__4638\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19800\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__19812\,
            I => \N__19797\
        );

    \I__4636\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19794\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__19806\,
            I => \N__19791\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__19803\,
            I => \c0.tx2.r_Bit_IndexZ0Z_2\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__19800\,
            I => \c0.tx2.r_Bit_IndexZ0Z_2\
        );

    \I__4632\ : Odrv4
    port map (
            O => \N__19797\,
            I => \c0.tx2.r_Bit_IndexZ0Z_2\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__19794\,
            I => \c0.tx2.r_Bit_IndexZ0Z_2\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__19791\,
            I => \c0.tx2.r_Bit_IndexZ0Z_2\
        );

    \I__4629\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19774\
        );

    \I__4628\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19774\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__19774\,
            I => \c0.tx2.N_12_0\
        );

    \I__4626\ : SRMux
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__4624\ : Sp12to4
    port map (
            O => \N__19765\,
            I => \N__19760\
        );

    \I__4623\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19757\
        );

    \I__4622\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19754\
        );

    \I__4621\ : Odrv12
    port map (
            O => \N__19760\,
            I => \c0.tx2.N_9_1\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__19757\,
            I => \c0.tx2.N_9_1\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__19754\,
            I => \c0.tx2.N_9_1\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19747\,
            I => \N__19742\
        );

    \I__4617\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19736\
        );

    \I__4616\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19736\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__19742\,
            I => \N__19733\
        );

    \I__4614\ : InMux
    port map (
            O => \N__19741\,
            I => \N__19730\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__19736\,
            I => \c0.tx2.r_Bit_IndexZ0Z_1\
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__19733\,
            I => \c0.tx2.r_Bit_IndexZ0Z_1\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__19730\,
            I => \c0.tx2.r_Bit_IndexZ0Z_1\
        );

    \I__4610\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19717\
        );

    \I__4609\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19714\
        );

    \I__4608\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19711\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__19720\,
            I => \N__19708\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19705\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__19714\,
            I => \N__19700\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__19711\,
            I => \N__19700\
        );

    \I__4603\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19697\
        );

    \I__4602\ : Span12Mux_v
    port map (
            O => \N__19705\,
            I => \N__19694\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__19700\,
            I => \N__19691\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__19697\,
            I => \c0.tx2_active\
        );

    \I__4599\ : Odrv12
    port map (
            O => \N__19694\,
            I => \c0.tx2_active\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__19691\,
            I => \c0.tx2_active\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19684\,
            I => \N__19681\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__19681\,
            I => \c0.N_170_0\
        );

    \I__4595\ : ClkMux
    port map (
            O => \N__19678\,
            I => \N__19375\
        );

    \I__4594\ : ClkMux
    port map (
            O => \N__19677\,
            I => \N__19375\
        );

    \I__4593\ : ClkMux
    port map (
            O => \N__19676\,
            I => \N__19375\
        );

    \I__4592\ : ClkMux
    port map (
            O => \N__19675\,
            I => \N__19375\
        );

    \I__4591\ : ClkMux
    port map (
            O => \N__19674\,
            I => \N__19375\
        );

    \I__4590\ : ClkMux
    port map (
            O => \N__19673\,
            I => \N__19375\
        );

    \I__4589\ : ClkMux
    port map (
            O => \N__19672\,
            I => \N__19375\
        );

    \I__4588\ : ClkMux
    port map (
            O => \N__19671\,
            I => \N__19375\
        );

    \I__4587\ : ClkMux
    port map (
            O => \N__19670\,
            I => \N__19375\
        );

    \I__4586\ : ClkMux
    port map (
            O => \N__19669\,
            I => \N__19375\
        );

    \I__4585\ : ClkMux
    port map (
            O => \N__19668\,
            I => \N__19375\
        );

    \I__4584\ : ClkMux
    port map (
            O => \N__19667\,
            I => \N__19375\
        );

    \I__4583\ : ClkMux
    port map (
            O => \N__19666\,
            I => \N__19375\
        );

    \I__4582\ : ClkMux
    port map (
            O => \N__19665\,
            I => \N__19375\
        );

    \I__4581\ : ClkMux
    port map (
            O => \N__19664\,
            I => \N__19375\
        );

    \I__4580\ : ClkMux
    port map (
            O => \N__19663\,
            I => \N__19375\
        );

    \I__4579\ : ClkMux
    port map (
            O => \N__19662\,
            I => \N__19375\
        );

    \I__4578\ : ClkMux
    port map (
            O => \N__19661\,
            I => \N__19375\
        );

    \I__4577\ : ClkMux
    port map (
            O => \N__19660\,
            I => \N__19375\
        );

    \I__4576\ : ClkMux
    port map (
            O => \N__19659\,
            I => \N__19375\
        );

    \I__4575\ : ClkMux
    port map (
            O => \N__19658\,
            I => \N__19375\
        );

    \I__4574\ : ClkMux
    port map (
            O => \N__19657\,
            I => \N__19375\
        );

    \I__4573\ : ClkMux
    port map (
            O => \N__19656\,
            I => \N__19375\
        );

    \I__4572\ : ClkMux
    port map (
            O => \N__19655\,
            I => \N__19375\
        );

    \I__4571\ : ClkMux
    port map (
            O => \N__19654\,
            I => \N__19375\
        );

    \I__4570\ : ClkMux
    port map (
            O => \N__19653\,
            I => \N__19375\
        );

    \I__4569\ : ClkMux
    port map (
            O => \N__19652\,
            I => \N__19375\
        );

    \I__4568\ : ClkMux
    port map (
            O => \N__19651\,
            I => \N__19375\
        );

    \I__4567\ : ClkMux
    port map (
            O => \N__19650\,
            I => \N__19375\
        );

    \I__4566\ : ClkMux
    port map (
            O => \N__19649\,
            I => \N__19375\
        );

    \I__4565\ : ClkMux
    port map (
            O => \N__19648\,
            I => \N__19375\
        );

    \I__4564\ : ClkMux
    port map (
            O => \N__19647\,
            I => \N__19375\
        );

    \I__4563\ : ClkMux
    port map (
            O => \N__19646\,
            I => \N__19375\
        );

    \I__4562\ : ClkMux
    port map (
            O => \N__19645\,
            I => \N__19375\
        );

    \I__4561\ : ClkMux
    port map (
            O => \N__19644\,
            I => \N__19375\
        );

    \I__4560\ : ClkMux
    port map (
            O => \N__19643\,
            I => \N__19375\
        );

    \I__4559\ : ClkMux
    port map (
            O => \N__19642\,
            I => \N__19375\
        );

    \I__4558\ : ClkMux
    port map (
            O => \N__19641\,
            I => \N__19375\
        );

    \I__4557\ : ClkMux
    port map (
            O => \N__19640\,
            I => \N__19375\
        );

    \I__4556\ : ClkMux
    port map (
            O => \N__19639\,
            I => \N__19375\
        );

    \I__4555\ : ClkMux
    port map (
            O => \N__19638\,
            I => \N__19375\
        );

    \I__4554\ : ClkMux
    port map (
            O => \N__19637\,
            I => \N__19375\
        );

    \I__4553\ : ClkMux
    port map (
            O => \N__19636\,
            I => \N__19375\
        );

    \I__4552\ : ClkMux
    port map (
            O => \N__19635\,
            I => \N__19375\
        );

    \I__4551\ : ClkMux
    port map (
            O => \N__19634\,
            I => \N__19375\
        );

    \I__4550\ : ClkMux
    port map (
            O => \N__19633\,
            I => \N__19375\
        );

    \I__4549\ : ClkMux
    port map (
            O => \N__19632\,
            I => \N__19375\
        );

    \I__4548\ : ClkMux
    port map (
            O => \N__19631\,
            I => \N__19375\
        );

    \I__4547\ : ClkMux
    port map (
            O => \N__19630\,
            I => \N__19375\
        );

    \I__4546\ : ClkMux
    port map (
            O => \N__19629\,
            I => \N__19375\
        );

    \I__4545\ : ClkMux
    port map (
            O => \N__19628\,
            I => \N__19375\
        );

    \I__4544\ : ClkMux
    port map (
            O => \N__19627\,
            I => \N__19375\
        );

    \I__4543\ : ClkMux
    port map (
            O => \N__19626\,
            I => \N__19375\
        );

    \I__4542\ : ClkMux
    port map (
            O => \N__19625\,
            I => \N__19375\
        );

    \I__4541\ : ClkMux
    port map (
            O => \N__19624\,
            I => \N__19375\
        );

    \I__4540\ : ClkMux
    port map (
            O => \N__19623\,
            I => \N__19375\
        );

    \I__4539\ : ClkMux
    port map (
            O => \N__19622\,
            I => \N__19375\
        );

    \I__4538\ : ClkMux
    port map (
            O => \N__19621\,
            I => \N__19375\
        );

    \I__4537\ : ClkMux
    port map (
            O => \N__19620\,
            I => \N__19375\
        );

    \I__4536\ : ClkMux
    port map (
            O => \N__19619\,
            I => \N__19375\
        );

    \I__4535\ : ClkMux
    port map (
            O => \N__19618\,
            I => \N__19375\
        );

    \I__4534\ : ClkMux
    port map (
            O => \N__19617\,
            I => \N__19375\
        );

    \I__4533\ : ClkMux
    port map (
            O => \N__19616\,
            I => \N__19375\
        );

    \I__4532\ : ClkMux
    port map (
            O => \N__19615\,
            I => \N__19375\
        );

    \I__4531\ : ClkMux
    port map (
            O => \N__19614\,
            I => \N__19375\
        );

    \I__4530\ : ClkMux
    port map (
            O => \N__19613\,
            I => \N__19375\
        );

    \I__4529\ : ClkMux
    port map (
            O => \N__19612\,
            I => \N__19375\
        );

    \I__4528\ : ClkMux
    port map (
            O => \N__19611\,
            I => \N__19375\
        );

    \I__4527\ : ClkMux
    port map (
            O => \N__19610\,
            I => \N__19375\
        );

    \I__4526\ : ClkMux
    port map (
            O => \N__19609\,
            I => \N__19375\
        );

    \I__4525\ : ClkMux
    port map (
            O => \N__19608\,
            I => \N__19375\
        );

    \I__4524\ : ClkMux
    port map (
            O => \N__19607\,
            I => \N__19375\
        );

    \I__4523\ : ClkMux
    port map (
            O => \N__19606\,
            I => \N__19375\
        );

    \I__4522\ : ClkMux
    port map (
            O => \N__19605\,
            I => \N__19375\
        );

    \I__4521\ : ClkMux
    port map (
            O => \N__19604\,
            I => \N__19375\
        );

    \I__4520\ : ClkMux
    port map (
            O => \N__19603\,
            I => \N__19375\
        );

    \I__4519\ : ClkMux
    port map (
            O => \N__19602\,
            I => \N__19375\
        );

    \I__4518\ : ClkMux
    port map (
            O => \N__19601\,
            I => \N__19375\
        );

    \I__4517\ : ClkMux
    port map (
            O => \N__19600\,
            I => \N__19375\
        );

    \I__4516\ : ClkMux
    port map (
            O => \N__19599\,
            I => \N__19375\
        );

    \I__4515\ : ClkMux
    port map (
            O => \N__19598\,
            I => \N__19375\
        );

    \I__4514\ : ClkMux
    port map (
            O => \N__19597\,
            I => \N__19375\
        );

    \I__4513\ : ClkMux
    port map (
            O => \N__19596\,
            I => \N__19375\
        );

    \I__4512\ : ClkMux
    port map (
            O => \N__19595\,
            I => \N__19375\
        );

    \I__4511\ : ClkMux
    port map (
            O => \N__19594\,
            I => \N__19375\
        );

    \I__4510\ : ClkMux
    port map (
            O => \N__19593\,
            I => \N__19375\
        );

    \I__4509\ : ClkMux
    port map (
            O => \N__19592\,
            I => \N__19375\
        );

    \I__4508\ : ClkMux
    port map (
            O => \N__19591\,
            I => \N__19375\
        );

    \I__4507\ : ClkMux
    port map (
            O => \N__19590\,
            I => \N__19375\
        );

    \I__4506\ : ClkMux
    port map (
            O => \N__19589\,
            I => \N__19375\
        );

    \I__4505\ : ClkMux
    port map (
            O => \N__19588\,
            I => \N__19375\
        );

    \I__4504\ : ClkMux
    port map (
            O => \N__19587\,
            I => \N__19375\
        );

    \I__4503\ : ClkMux
    port map (
            O => \N__19586\,
            I => \N__19375\
        );

    \I__4502\ : ClkMux
    port map (
            O => \N__19585\,
            I => \N__19375\
        );

    \I__4501\ : ClkMux
    port map (
            O => \N__19584\,
            I => \N__19375\
        );

    \I__4500\ : ClkMux
    port map (
            O => \N__19583\,
            I => \N__19375\
        );

    \I__4499\ : ClkMux
    port map (
            O => \N__19582\,
            I => \N__19375\
        );

    \I__4498\ : ClkMux
    port map (
            O => \N__19581\,
            I => \N__19375\
        );

    \I__4497\ : ClkMux
    port map (
            O => \N__19580\,
            I => \N__19375\
        );

    \I__4496\ : ClkMux
    port map (
            O => \N__19579\,
            I => \N__19375\
        );

    \I__4495\ : ClkMux
    port map (
            O => \N__19578\,
            I => \N__19375\
        );

    \I__4494\ : GlobalMux
    port map (
            O => \N__19375\,
            I => \N__19372\
        );

    \I__4493\ : gio2CtrlBuf
    port map (
            O => \N__19372\,
            I => \CLK_c_g\
        );

    \I__4492\ : SRMux
    port map (
            O => \N__19369\,
            I => \N__19366\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__19366\,
            I => \N__19362\
        );

    \I__4490\ : SRMux
    port map (
            O => \N__19365\,
            I => \N__19359\
        );

    \I__4489\ : Span4Mux_v
    port map (
            O => \N__19362\,
            I => \N__19354\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__19359\,
            I => \N__19354\
        );

    \I__4487\ : Span4Mux_h
    port map (
            O => \N__19354\,
            I => \N__19350\
        );

    \I__4486\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19347\
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__19350\,
            I => \c0.tx2_transmit_0_sqmuxa\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__19347\,
            I => \c0.tx2_transmit_0_sqmuxa\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19336\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19341\,
            I => \N__19333\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__19340\,
            I => \N__19330\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19327\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19336\,
            I => \N__19323\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__19333\,
            I => \N__19320\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19317\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__19327\,
            I => \N__19314\
        );

    \I__4475\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19311\
        );

    \I__4474\ : Span4Mux_h
    port map (
            O => \N__19323\,
            I => \N__19308\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__19320\,
            I => \N__19305\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__19317\,
            I => \N__19300\
        );

    \I__4471\ : Span4Mux_h
    port map (
            O => \N__19314\,
            I => \N__19300\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__19311\,
            I => \c0.wait_for_transmissionZ0\
        );

    \I__4469\ : Odrv4
    port map (
            O => \N__19308\,
            I => \c0.wait_for_transmissionZ0\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__19305\,
            I => \c0.wait_for_transmissionZ0\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__19300\,
            I => \c0.wait_for_transmissionZ0\
        );

    \I__4466\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19288\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19288\,
            I => \N__19284\
        );

    \I__4464\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19281\
        );

    \I__4463\ : Span12Mux_h
    port map (
            O => \N__19284\,
            I => \N__19278\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__19281\,
            I => \N__19275\
        );

    \I__4461\ : Odrv12
    port map (
            O => \N__19278\,
            I => \c0.i12_THRU_CO\
        );

    \I__4460\ : Odrv12
    port map (
            O => \N__19275\,
            I => \c0.i12_THRU_CO\
        );

    \I__4459\ : IoInMux
    port map (
            O => \N__19270\,
            I => \N__19267\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__19267\,
            I => \N__19264\
        );

    \I__4457\ : Span12Mux_s4_h
    port map (
            O => \N__19264\,
            I => \N__19261\
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__19261\,
            I => \c0.data_in_frame_0__0_sqmuxa\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__19258\,
            I => \N__19255\
        );

    \I__4454\ : InMux
    port map (
            O => \N__19255\,
            I => \N__19252\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__19252\,
            I => \c0.tx2.N_214_0\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19240\
        );

    \I__4451\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19240\
        );

    \I__4450\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19237\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19232\
        );

    \I__4448\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19232\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__19240\,
            I => \c0.tx2.r_Clock_Count12_THRU_CO\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__19237\,
            I => \c0.tx2.r_Clock_Count12_THRU_CO\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__19232\,
            I => \c0.tx2.r_Clock_Count12_THRU_CO\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__19225\,
            I => \c0.tx2.N_17_0_cascade_\
        );

    \I__4443\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19215\
        );

    \I__4442\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19212\
        );

    \I__4441\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19205\
        );

    \I__4440\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19205\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19218\,
            I => \N__19205\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__19215\,
            I => \c0.tx2.r_SM_Main_dup_4\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__19212\,
            I => \c0.tx2.r_SM_Main_dup_4\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__19205\,
            I => \c0.tx2.r_SM_Main_dup_4\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__19198\,
            I => \N__19195\
        );

    \I__4434\ : InMux
    port map (
            O => \N__19195\,
            I => \N__19186\
        );

    \I__4433\ : InMux
    port map (
            O => \N__19194\,
            I => \N__19186\
        );

    \I__4432\ : InMux
    port map (
            O => \N__19193\,
            I => \N__19183\
        );

    \I__4431\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19178\
        );

    \I__4430\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19178\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__19186\,
            I => \c0.tx2.r_Bit_IndexZ1Z_0\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__19183\,
            I => \c0.tx2.r_Bit_IndexZ1Z_0\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19178\,
            I => \c0.tx2.r_Bit_IndexZ1Z_0\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__19171\,
            I => \c0.tx2.N_212_0_cascade_\
        );

    \I__4425\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19161\
        );

    \I__4424\ : InMux
    port map (
            O => \N__19167\,
            I => \N__19158\
        );

    \I__4423\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19151\
        );

    \I__4422\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19151\
        );

    \I__4421\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19151\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__19161\,
            I => \c0.tx2.r_SM_Main_dup_1\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__19158\,
            I => \c0.tx2.r_SM_Main_dup_1\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__19151\,
            I => \c0.tx2.r_SM_Main_dup_1\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__19144\,
            I => \c0.tx2.N_496_cascade_\
        );

    \I__4416\ : CascadeMux
    port map (
            O => \N__19141\,
            I => \N__19135\
        );

    \I__4415\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19127\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19127\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19122\
        );

    \I__4412\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19122\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19115\
        );

    \I__4410\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19115\
        );

    \I__4409\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19115\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19127\,
            I => \c0.tx2.r_SM_Main_dup_2\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__19122\,
            I => \c0.tx2.r_SM_Main_dup_2\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__19115\,
            I => \c0.tx2.r_SM_Main_dup_2\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19100\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19107\,
            I => \N__19100\
        );

    \I__4403\ : InMux
    port map (
            O => \N__19106\,
            I => \N__19097\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19105\,
            I => \N__19094\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__19100\,
            I => \N__19091\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19097\,
            I => \N__19088\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__19094\,
            I => \N__19085\
        );

    \I__4398\ : Odrv12
    port map (
            O => \N__19091\,
            I => \c0.tx2.N_171_0\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__19088\,
            I => \c0.tx2.N_171_0\
        );

    \I__4396\ : Odrv4
    port map (
            O => \N__19085\,
            I => \c0.tx2.N_171_0\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19074\
        );

    \I__4394\ : InMux
    port map (
            O => \N__19077\,
            I => \N__19071\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__19074\,
            I => \c0.tx2.N_17_0\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__19071\,
            I => \c0.tx2.N_17_0\
        );

    \I__4391\ : CascadeMux
    port map (
            O => \N__19066\,
            I => \N__19063\
        );

    \I__4390\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19060\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__19060\,
            I => \c0.tx2.N_212_0\
        );

    \I__4388\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19051\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19051\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__19051\,
            I => \c0.tx2.N_493\
        );

    \I__4385\ : InMux
    port map (
            O => \N__19048\,
            I => \N__19042\
        );

    \I__4384\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19039\
        );

    \I__4383\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19036\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19033\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__19042\,
            I => \c0.tx2.r_SM_Main_dup_3\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__19039\,
            I => \c0.tx2.r_SM_Main_dup_3\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__19036\,
            I => \c0.tx2.r_SM_Main_dup_3\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__19033\,
            I => \c0.tx2.r_SM_Main_dup_3\
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__19024\,
            I => \N__19021\
        );

    \I__4376\ : InMux
    port map (
            O => \N__19021\,
            I => \N__19014\
        );

    \I__4375\ : InMux
    port map (
            O => \N__19020\,
            I => \N__19014\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19011\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__19014\,
            I => \c0.tx2.r_Clock_CountZ0Z_2\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__19011\,
            I => \c0.tx2.r_Clock_CountZ0Z_2\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__19006\,
            I => \N__19003\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19003\,
            I => \N__18996\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19002\,
            I => \N__18996\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18993\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__18996\,
            I => \c0.tx2.r_Clock_CountZ0Z_1\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__18993\,
            I => \c0.tx2.r_Clock_CountZ0Z_1\
        );

    \I__4365\ : CascadeMux
    port map (
            O => \N__18988\,
            I => \N__18984\
        );

    \I__4364\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18978\
        );

    \I__4363\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18978\
        );

    \I__4362\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18975\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__18978\,
            I => \c0.tx2.r_Clock_CountZ0Z_3\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__18975\,
            I => \c0.tx2.r_Clock_CountZ0Z_3\
        );

    \I__4359\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18963\
        );

    \I__4358\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18963\
        );

    \I__4357\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18960\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__18963\,
            I => \c0.tx2.r_Clock_CountZ0Z_0\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__18960\,
            I => \c0.tx2.r_Clock_CountZ0Z_0\
        );

    \I__4354\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18949\
        );

    \I__4353\ : InMux
    port map (
            O => \N__18954\,
            I => \N__18949\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__18949\,
            I => \N__18944\
        );

    \I__4351\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18939\
        );

    \I__4350\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18939\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__18944\,
            I => \c0.tx2.N_16_0\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__18939\,
            I => \c0.tx2.N_16_0\
        );

    \I__4347\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18930\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__18933\,
            I => \N__18927\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__18930\,
            I => \N__18924\
        );

    \I__4344\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18921\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__18924\,
            I => \c0.tx2.r_Clock_Count_0_sqmuxa\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__18921\,
            I => \c0.tx2.r_Clock_Count_0_sqmuxa\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__18916\,
            I => \c0.tx2.N_83_0_cascade_\
        );

    \I__4340\ : CascadeMux
    port map (
            O => \N__18913\,
            I => \c0.N_90_dup_cascade_\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__18910\,
            I => \c0.tx2.i97_mux_cascade_\
        );

    \I__4338\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18904\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__18904\,
            I => \c0.tx2.r_SM_Main_illegal_0\
        );

    \I__4336\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18898\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18895\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__18895\,
            I => \N__18891\
        );

    \I__4333\ : InMux
    port map (
            O => \N__18894\,
            I => \N__18888\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__18891\,
            I => \c0.d_4_0\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__18888\,
            I => \c0.d_4_0\
        );

    \I__4330\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18880\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__18880\,
            I => \N__18877\
        );

    \I__4328\ : Span4Mux_v
    port map (
            O => \N__18877\,
            I => \N__18873\
        );

    \I__4327\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18870\
        );

    \I__4326\ : Sp12to4
    port map (
            O => \N__18873\,
            I => \N__18864\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__18870\,
            I => \N__18864\
        );

    \I__4324\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18861\
        );

    \I__4323\ : Odrv12
    port map (
            O => \N__18864\,
            I => \c0.d_4_8\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__18861\,
            I => \c0.d_4_8\
        );

    \I__4321\ : InMux
    port map (
            O => \N__18856\,
            I => \N__18853\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__18853\,
            I => \N__18850\
        );

    \I__4319\ : Span4Mux_h
    port map (
            O => \N__18850\,
            I => \N__18844\
        );

    \I__4318\ : InMux
    port map (
            O => \N__18849\,
            I => \N__18839\
        );

    \I__4317\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18839\
        );

    \I__4316\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18836\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__18844\,
            I => \c0.d_4_16\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__18839\,
            I => \c0.d_4_16\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__18836\,
            I => \c0.d_4_16\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__18829\,
            I => \N__18826\
        );

    \I__4311\ : InMux
    port map (
            O => \N__18826\,
            I => \N__18823\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__18823\,
            I => \N__18820\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__18820\,
            I => \N__18815\
        );

    \I__4308\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18812\
        );

    \I__4307\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18809\
        );

    \I__4306\ : Span4Mux_h
    port map (
            O => \N__18815\,
            I => \N__18804\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__18812\,
            I => \N__18804\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__18809\,
            I => \c0.d_4_24\
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__18804\,
            I => \c0.d_4_24\
        );

    \I__4302\ : InMux
    port map (
            O => \N__18799\,
            I => \N__18792\
        );

    \I__4301\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18788\
        );

    \I__4300\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18785\
        );

    \I__4299\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18779\
        );

    \I__4298\ : InMux
    port map (
            O => \N__18795\,
            I => \N__18779\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__18792\,
            I => \N__18776\
        );

    \I__4296\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18773\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__18788\,
            I => \N__18768\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__18785\,
            I => \N__18768\
        );

    \I__4293\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18765\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__18779\,
            I => \N__18759\
        );

    \I__4291\ : Span4Mux_h
    port map (
            O => \N__18776\,
            I => \N__18754\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__18773\,
            I => \N__18754\
        );

    \I__4289\ : Span4Mux_v
    port map (
            O => \N__18768\,
            I => \N__18749\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__18765\,
            I => \N__18749\
        );

    \I__4287\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18746\
        );

    \I__4286\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18741\
        );

    \I__4285\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18741\
        );

    \I__4284\ : Odrv12
    port map (
            O => \N__18759\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__18754\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__18749\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__18746\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__18741\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4279\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18727\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__18727\,
            I => \c0.tx2_data_RNO_3Z0Z_0\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__18724\,
            I => \c0.tx2_data_RNO_4Z0Z_0_cascade_\
        );

    \I__4276\ : InMux
    port map (
            O => \N__18721\,
            I => \N__18705\
        );

    \I__4275\ : InMux
    port map (
            O => \N__18720\,
            I => \N__18700\
        );

    \I__4274\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18700\
        );

    \I__4273\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18697\
        );

    \I__4272\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18690\
        );

    \I__4271\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18690\
        );

    \I__4270\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18690\
        );

    \I__4269\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18687\
        );

    \I__4268\ : InMux
    port map (
            O => \N__18713\,
            I => \N__18684\
        );

    \I__4267\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18681\
        );

    \I__4266\ : InMux
    port map (
            O => \N__18711\,
            I => \N__18674\
        );

    \I__4265\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18674\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18674\
        );

    \I__4263\ : InMux
    port map (
            O => \N__18708\,
            I => \N__18671\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__18705\,
            I => \N__18666\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__18700\,
            I => \N__18666\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__18697\,
            I => \N__18663\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__18690\,
            I => \N__18658\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__18687\,
            I => \N__18658\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__18684\,
            I => \N__18649\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__18681\,
            I => \N__18649\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18646\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__18671\,
            I => \N__18641\
        );

    \I__4253\ : Span4Mux_v
    port map (
            O => \N__18666\,
            I => \N__18641\
        );

    \I__4252\ : Span4Mux_v
    port map (
            O => \N__18663\,
            I => \N__18636\
        );

    \I__4251\ : Span4Mux_h
    port map (
            O => \N__18658\,
            I => \N__18636\
        );

    \I__4250\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18633\
        );

    \I__4249\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18626\
        );

    \I__4248\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18626\
        );

    \I__4247\ : InMux
    port map (
            O => \N__18654\,
            I => \N__18626\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__18649\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4245\ : Odrv12
    port map (
            O => \N__18646\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__18641\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__18636\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__18633\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__18626\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4240\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18610\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__18610\,
            I => \N__18607\
        );

    \I__4238\ : Odrv12
    port map (
            O => \N__18607\,
            I => \c0.tx2_data_RNO_1Z0Z_0\
        );

    \I__4237\ : CascadeMux
    port map (
            O => \N__18604\,
            I => \c0.m146_ns_1_cascade_\
        );

    \I__4236\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18598\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__18598\,
            I => \c0.tx2.r_Tx_DataZ0Z_0\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__18595\,
            I => \N__18583\
        );

    \I__4233\ : CascadeMux
    port map (
            O => \N__18594\,
            I => \N__18579\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__18593\,
            I => \N__18573\
        );

    \I__4231\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18562\
        );

    \I__4230\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18555\
        );

    \I__4229\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18555\
        );

    \I__4228\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18555\
        );

    \I__4227\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18550\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18550\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18543\
        );

    \I__4224\ : InMux
    port map (
            O => \N__18583\,
            I => \N__18543\
        );

    \I__4223\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18543\
        );

    \I__4222\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18536\
        );

    \I__4221\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18536\
        );

    \I__4220\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18536\
        );

    \I__4219\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18533\
        );

    \I__4218\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18528\
        );

    \I__4217\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18521\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18521\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__18570\,
            I => \N__18515\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18510\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18501\
        );

    \I__4212\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18501\
        );

    \I__4211\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18501\
        );

    \I__4210\ : InMux
    port map (
            O => \N__18565\,
            I => \N__18501\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__18562\,
            I => \N__18496\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__18555\,
            I => \N__18496\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18493\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__18543\,
            I => \N__18490\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__18536\,
            I => \N__18485\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__18533\,
            I => \N__18485\
        );

    \I__4203\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18479\
        );

    \I__4202\ : InMux
    port map (
            O => \N__18531\,
            I => \N__18476\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__18528\,
            I => \N__18473\
        );

    \I__4200\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18468\
        );

    \I__4199\ : InMux
    port map (
            O => \N__18526\,
            I => \N__18468\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__18521\,
            I => \N__18465\
        );

    \I__4197\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18458\
        );

    \I__4196\ : InMux
    port map (
            O => \N__18519\,
            I => \N__18458\
        );

    \I__4195\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18458\
        );

    \I__4194\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18453\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18514\,
            I => \N__18453\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18450\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__18510\,
            I => \N__18443\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__18501\,
            I => \N__18443\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__18496\,
            I => \N__18443\
        );

    \I__4188\ : Span4Mux_h
    port map (
            O => \N__18493\,
            I => \N__18436\
        );

    \I__4187\ : Span4Mux_v
    port map (
            O => \N__18490\,
            I => \N__18436\
        );

    \I__4186\ : Span4Mux_h
    port map (
            O => \N__18485\,
            I => \N__18436\
        );

    \I__4185\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18429\
        );

    \I__4184\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18429\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18429\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__18479\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__18476\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4180\ : Odrv12
    port map (
            O => \N__18473\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__18468\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4178\ : Odrv12
    port map (
            O => \N__18465\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__18458\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__18453\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__18450\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__18443\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__18436\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__18429\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18403\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__18403\,
            I => \N__18396\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18402\,
            I => \N__18393\
        );

    \I__4168\ : InMux
    port map (
            O => \N__18401\,
            I => \N__18390\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18400\,
            I => \N__18385\
        );

    \I__4166\ : InMux
    port map (
            O => \N__18399\,
            I => \N__18385\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__18396\,
            I => \c0.d_4_32\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__18393\,
            I => \c0.d_4_32\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__18390\,
            I => \c0.d_4_32\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__18385\,
            I => \c0.d_4_32\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__18376\,
            I => \N__18366\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__18375\,
            I => \N__18362\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__18374\,
            I => \N__18358\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__18373\,
            I => \N__18349\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__18372\,
            I => \N__18344\
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__18371\,
            I => \N__18341\
        );

    \I__4155\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18334\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18334\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18366\,
            I => \N__18334\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18324\
        );

    \I__4151\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18324\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18319\
        );

    \I__4149\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18319\
        );

    \I__4148\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18312\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18312\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18312\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18309\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \N__18306\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__18352\,
            I => \N__18298\
        );

    \I__4142\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18293\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18293\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18286\
        );

    \I__4139\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18286\
        );

    \I__4138\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18286\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__18334\,
            I => \N__18283\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__18333\,
            I => \N__18279\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__18332\,
            I => \N__18275\
        );

    \I__4134\ : CascadeMux
    port map (
            O => \N__18331\,
            I => \N__18271\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__18330\,
            I => \N__18268\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__18329\,
            I => \N__18264\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__18324\,
            I => \N__18261\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__18319\,
            I => \N__18258\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__18312\,
            I => \N__18253\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__18309\,
            I => \N__18253\
        );

    \I__4127\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18248\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18248\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18237\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18237\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18237\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18237\
        );

    \I__4121\ : InMux
    port map (
            O => \N__18298\,
            I => \N__18237\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__18293\,
            I => \N__18232\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__18286\,
            I => \N__18232\
        );

    \I__4118\ : Span4Mux_h
    port map (
            O => \N__18283\,
            I => \N__18229\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18224\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18224\
        );

    \I__4115\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18215\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18215\
        );

    \I__4113\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18215\
        );

    \I__4112\ : InMux
    port map (
            O => \N__18271\,
            I => \N__18215\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18208\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18208\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18208\
        );

    \I__4108\ : Span4Mux_v
    port map (
            O => \N__18261\,
            I => \N__18199\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__18258\,
            I => \N__18199\
        );

    \I__4106\ : Span4Mux_v
    port map (
            O => \N__18253\,
            I => \N__18199\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18248\,
            I => \N__18199\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__18237\,
            I => \N__18194\
        );

    \I__4103\ : Span4Mux_h
    port map (
            O => \N__18232\,
            I => \N__18194\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__18229\,
            I => \c0.N_204_mux\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__18224\,
            I => \c0.N_204_mux\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__18215\,
            I => \c0.N_204_mux\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__18208\,
            I => \c0.N_204_mux\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__18199\,
            I => \c0.N_204_mux\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__18194\,
            I => \c0.N_204_mux\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18181\,
            I => \N__18178\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18178\,
            I => \N__18175\
        );

    \I__4094\ : Span4Mux_h
    port map (
            O => \N__18175\,
            I => \N__18170\
        );

    \I__4093\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18167\
        );

    \I__4092\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18164\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__18170\,
            I => \c0.d_4_40\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__18167\,
            I => \c0.d_4_40\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18164\,
            I => \c0.d_4_40\
        );

    \I__4088\ : InMux
    port map (
            O => \N__18157\,
            I => \N__18154\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18154\,
            I => \c0.tx2_data_RNO_0Z0Z_0\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18151\,
            I => \c0.tx2.un1_r_Clock_Count_cry_0\
        );

    \I__4085\ : InMux
    port map (
            O => \N__18148\,
            I => \c0.tx2.un1_r_Clock_Count_cry_1\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18145\,
            I => \c0.tx2.un1_r_Clock_Count_cry_2\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18142\,
            I => \N__18138\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18135\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__18138\,
            I => \N__18132\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18135\,
            I => \N__18129\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__18132\,
            I => \c0.N_164_0\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__18129\,
            I => \c0.N_164_0\
        );

    \I__4077\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18121\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__18121\,
            I => \N__18118\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__18118\,
            I => \N__18114\
        );

    \I__4074\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18111\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__18114\,
            I => \c0.d_4_22\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__18111\,
            I => \c0.d_4_22\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__18106\,
            I => \N__18103\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18100\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__18100\,
            I => \N__18097\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__18097\,
            I => \N__18091\
        );

    \I__4067\ : InMux
    port map (
            O => \N__18096\,
            I => \N__18088\
        );

    \I__4066\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18085\
        );

    \I__4065\ : InMux
    port map (
            O => \N__18094\,
            I => \N__18082\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__18091\,
            I => \c0.d_4_30\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__18088\,
            I => \c0.d_4_30\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__18085\,
            I => \c0.d_4_30\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__18082\,
            I => \c0.d_4_30\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__18073\,
            I => \N__18070\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18067\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__18067\,
            I => \N__18064\
        );

    \I__4057\ : Odrv4
    port map (
            O => \N__18064\,
            I => \c0.tx2_data_RNO_4Z0Z_6\
        );

    \I__4056\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18058\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__18058\,
            I => \N__18055\
        );

    \I__4054\ : Span12Mux_h
    port map (
            O => \N__18055\,
            I => \N__18051\
        );

    \I__4053\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18048\
        );

    \I__4052\ : Odrv12
    port map (
            O => \N__18051\,
            I => \c0.d_4_4\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__18048\,
            I => \c0.d_4_4\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18043\,
            I => \N__18040\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__18040\,
            I => \N__18037\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__18037\,
            I => \N__18031\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18036\,
            I => \N__18026\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18026\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18034\,
            I => \N__18023\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__18031\,
            I => \c0.d_4_12\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18026\,
            I => \c0.d_4_12\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__18023\,
            I => \c0.d_4_12\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__18016\,
            I => \N__18013\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18013\,
            I => \N__18010\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__18010\,
            I => \N__18007\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__18007\,
            I => \c0.tx2_data_RNO_3Z0Z_4\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__18004\,
            I => \N__18000\
        );

    \I__4036\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17997\
        );

    \I__4035\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17994\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__17997\,
            I => \N__17988\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__17994\,
            I => \N__17988\
        );

    \I__4032\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17985\
        );

    \I__4031\ : Span4Mux_v
    port map (
            O => \N__17988\,
            I => \N__17981\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__17985\,
            I => \N__17978\
        );

    \I__4029\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17975\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__17981\,
            I => \c0.d_4_28\
        );

    \I__4027\ : Odrv12
    port map (
            O => \N__17978\,
            I => \c0.d_4_28\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__17975\,
            I => \c0.d_4_28\
        );

    \I__4025\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17965\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__17965\,
            I => \N__17961\
        );

    \I__4023\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17957\
        );

    \I__4022\ : Span4Mux_h
    port map (
            O => \N__17961\,
            I => \N__17954\
        );

    \I__4021\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17951\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__17957\,
            I => \N__17948\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__17954\,
            I => \c0.d_4_20\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__17951\,
            I => \c0.d_4_20\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__17948\,
            I => \c0.d_4_20\
        );

    \I__4016\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17938\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__17938\,
            I => \N__17935\
        );

    \I__4014\ : Span4Mux_v
    port map (
            O => \N__17935\,
            I => \N__17932\
        );

    \I__4013\ : Odrv4
    port map (
            O => \N__17932\,
            I => \c0.tx2_data_RNO_4Z0Z_4\
        );

    \I__4012\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17926\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__17926\,
            I => \N__17923\
        );

    \I__4010\ : Span4Mux_h
    port map (
            O => \N__17923\,
            I => \N__17919\
        );

    \I__4009\ : InMux
    port map (
            O => \N__17922\,
            I => \N__17916\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__17919\,
            I => \c0.d_4_13\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__17916\,
            I => \c0.d_4_13\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__17911\,
            I => \N__17908\
        );

    \I__4005\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17905\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__17905\,
            I => \N__17901\
        );

    \I__4003\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17897\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__17901\,
            I => \N__17894\
        );

    \I__4001\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17891\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17888\
        );

    \I__3999\ : Odrv4
    port map (
            O => \N__17894\,
            I => \c0.d_4_5\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__17891\,
            I => \c0.d_4_5\
        );

    \I__3997\ : Odrv12
    port map (
            O => \N__17888\,
            I => \c0.d_4_5\
        );

    \I__3996\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17878\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__17878\,
            I => \c0.tx2_data_RNO_3Z0Z_5\
        );

    \I__3994\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17871\
        );

    \I__3993\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17868\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__17871\,
            I => \c0.byte_transmit_counter2Z0Z_7\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__17868\,
            I => \c0.byte_transmit_counter2Z0Z_7\
        );

    \I__3990\ : InMux
    port map (
            O => \N__17863\,
            I => \N__17859\
        );

    \I__3989\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17856\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__17859\,
            I => \c0.byte_transmit_counter2Z0Z_3\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__17856\,
            I => \c0.byte_transmit_counter2Z0Z_3\
        );

    \I__3986\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17847\
        );

    \I__3985\ : InMux
    port map (
            O => \N__17850\,
            I => \N__17844\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__17847\,
            I => \c0.byte_transmit_counter2Z0Z_6\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__17844\,
            I => \c0.byte_transmit_counter2Z0Z_6\
        );

    \I__3982\ : InMux
    port map (
            O => \N__17839\,
            I => \N__17835\
        );

    \I__3981\ : InMux
    port map (
            O => \N__17838\,
            I => \N__17832\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__17835\,
            I => \c0.byte_transmit_counter2Z0Z_5\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__17832\,
            I => \c0.byte_transmit_counter2Z0Z_5\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__17827\,
            I => \c0.m45_0_0_cascade_\
        );

    \I__3977\ : InMux
    port map (
            O => \N__17824\,
            I => \N__17820\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17817\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__17820\,
            I => \c0.byte_transmit_counter2Z0Z_4\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__17817\,
            I => \c0.byte_transmit_counter2Z0Z_4\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__17812\,
            I => \c0.N_204_mux_cascade_\
        );

    \I__3972\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17806\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__17806\,
            I => \N__17802\
        );

    \I__3970\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17799\
        );

    \I__3969\ : Span4Mux_h
    port map (
            O => \N__17802\,
            I => \N__17796\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__17799\,
            I => \c0.N_215_mux\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__17796\,
            I => \c0.N_215_mux\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__17791\,
            I => \N__17787\
        );

    \I__3965\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17784\
        );

    \I__3964\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17781\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__17784\,
            I => \N__17776\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__17781\,
            I => \N__17776\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__17776\,
            I => \N__17772\
        );

    \I__3960\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17769\
        );

    \I__3959\ : Span4Mux_h
    port map (
            O => \N__17772\,
            I => \N__17766\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__17769\,
            I => \c0.data_in_7_Z0Z_2\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__17766\,
            I => \c0.data_in_7_Z0Z_2\
        );

    \I__3956\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17758\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17754\
        );

    \I__3954\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17751\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__17754\,
            I => \N__17746\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__17751\,
            I => \N__17746\
        );

    \I__3951\ : Span4Mux_h
    port map (
            O => \N__17746\,
            I => \N__17742\
        );

    \I__3950\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17739\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__17742\,
            I => \c0.data_in_6_Z0Z_2\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__17739\,
            I => \c0.data_in_6_Z0Z_2\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__17734\,
            I => \N__17731\
        );

    \I__3946\ : InMux
    port map (
            O => \N__17731\,
            I => \N__17728\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__17728\,
            I => \N__17712\
        );

    \I__3944\ : CEMux
    port map (
            O => \N__17727\,
            I => \N__17683\
        );

    \I__3943\ : CEMux
    port map (
            O => \N__17726\,
            I => \N__17683\
        );

    \I__3942\ : CEMux
    port map (
            O => \N__17725\,
            I => \N__17683\
        );

    \I__3941\ : CEMux
    port map (
            O => \N__17724\,
            I => \N__17683\
        );

    \I__3940\ : CEMux
    port map (
            O => \N__17723\,
            I => \N__17683\
        );

    \I__3939\ : CEMux
    port map (
            O => \N__17722\,
            I => \N__17683\
        );

    \I__3938\ : CEMux
    port map (
            O => \N__17721\,
            I => \N__17683\
        );

    \I__3937\ : CEMux
    port map (
            O => \N__17720\,
            I => \N__17683\
        );

    \I__3936\ : CEMux
    port map (
            O => \N__17719\,
            I => \N__17683\
        );

    \I__3935\ : CEMux
    port map (
            O => \N__17718\,
            I => \N__17683\
        );

    \I__3934\ : CEMux
    port map (
            O => \N__17717\,
            I => \N__17683\
        );

    \I__3933\ : CEMux
    port map (
            O => \N__17716\,
            I => \N__17683\
        );

    \I__3932\ : CEMux
    port map (
            O => \N__17715\,
            I => \N__17683\
        );

    \I__3931\ : Glb2LocalMux
    port map (
            O => \N__17712\,
            I => \N__17683\
        );

    \I__3930\ : GlobalMux
    port map (
            O => \N__17683\,
            I => \N__17680\
        );

    \I__3929\ : gio2CtrlBuf
    port map (
            O => \N__17680\,
            I => \c0.rx_data_ready_g\
        );

    \I__3928\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17673\
        );

    \I__3927\ : InMux
    port map (
            O => \N__17676\,
            I => \N__17670\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__17673\,
            I => \N__17667\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__17670\,
            I => \N__17664\
        );

    \I__3924\ : Span4Mux_v
    port map (
            O => \N__17667\,
            I => \N__17659\
        );

    \I__3923\ : Span4Mux_v
    port map (
            O => \N__17664\,
            I => \N__17659\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__17659\,
            I => \c0.d_4_45\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__17656\,
            I => \N__17653\
        );

    \I__3920\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17650\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__17650\,
            I => \N__17644\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__17649\,
            I => \N__17641\
        );

    \I__3917\ : InMux
    port map (
            O => \N__17648\,
            I => \N__17636\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17636\
        );

    \I__3915\ : Span4Mux_h
    port map (
            O => \N__17644\,
            I => \N__17633\
        );

    \I__3914\ : InMux
    port map (
            O => \N__17641\,
            I => \N__17630\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__17636\,
            I => \N__17627\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__17633\,
            I => \c0.d_4_37\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__17630\,
            I => \c0.d_4_37\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__17627\,
            I => \c0.d_4_37\
        );

    \I__3909\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17613\
        );

    \I__3908\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17613\
        );

    \I__3907\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17610\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__17613\,
            I => \N__17607\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__17610\,
            I => \N__17603\
        );

    \I__3904\ : Span4Mux_v
    port map (
            O => \N__17607\,
            I => \N__17600\
        );

    \I__3903\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17597\
        );

    \I__3902\ : Odrv12
    port map (
            O => \N__17603\,
            I => \c0.d_4_29\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__17600\,
            I => \c0.d_4_29\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__17597\,
            I => \c0.d_4_29\
        );

    \I__3899\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17587\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__17587\,
            I => \N__17584\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__17584\,
            I => \N__17579\
        );

    \I__3896\ : InMux
    port map (
            O => \N__17583\,
            I => \N__17576\
        );

    \I__3895\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17573\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__17579\,
            I => \c0.d_4_21\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__17576\,
            I => \c0.d_4_21\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__17573\,
            I => \c0.d_4_21\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__17566\,
            I => \c0.tx2_data_RNO_4Z0Z_5_cascade_\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17560\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__17560\,
            I => \c0.tx2_data_RNO_0Z0Z_5\
        );

    \I__3888\ : CascadeMux
    port map (
            O => \N__17557\,
            I => \c0.m75_ns_1_cascade_\
        );

    \I__3887\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17551\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__17551\,
            I => \N__17548\
        );

    \I__3885\ : Span4Mux_h
    port map (
            O => \N__17548\,
            I => \N__17545\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__17545\,
            I => \c0.tx2.r_Tx_DataZ0Z_5\
        );

    \I__3883\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17539\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__17539\,
            I => \N__17536\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__17536\,
            I => \c0.data_in_frame_6_Z0Z_5\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__17533\,
            I => \N__17530\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17527\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__17527\,
            I => \N__17524\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__17524\,
            I => \c0.data_in_frame_7_Z0Z_5\
        );

    \I__3876\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17518\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__17518\,
            I => \c0.tx2_data_RNO_1Z0Z_5\
        );

    \I__3874\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17511\
        );

    \I__3873\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17508\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__17511\,
            I => \N__17505\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__17508\,
            I => \N__17501\
        );

    \I__3870\ : Span4Mux_v
    port map (
            O => \N__17505\,
            I => \N__17498\
        );

    \I__3869\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17495\
        );

    \I__3868\ : Span12Mux_v
    port map (
            O => \N__17501\,
            I => \N__17492\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__17498\,
            I => \c0.d_4_47\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17495\,
            I => \c0.d_4_47\
        );

    \I__3865\ : Odrv12
    port map (
            O => \N__17492\,
            I => \c0.d_4_47\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__17485\,
            I => \N__17481\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__17484\,
            I => \N__17478\
        );

    \I__3862\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17475\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17478\,
            I => \N__17472\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__17475\,
            I => \N__17469\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17466\
        );

    \I__3858\ : Span4Mux_h
    port map (
            O => \N__17469\,
            I => \N__17460\
        );

    \I__3857\ : Span4Mux_h
    port map (
            O => \N__17466\,
            I => \N__17460\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17465\,
            I => \N__17457\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__17460\,
            I => \c0.d_4_39\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17457\,
            I => \c0.d_4_39\
        );

    \I__3853\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17449\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__17449\,
            I => \N__17446\
        );

    \I__3851\ : Span4Mux_v
    port map (
            O => \N__17446\,
            I => \N__17443\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__17443\,
            I => \c0.tx2_data_RNO_0Z0Z_7\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17437\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__17437\,
            I => \N__17434\
        );

    \I__3847\ : Span4Mux_v
    port map (
            O => \N__17434\,
            I => \N__17431\
        );

    \I__3846\ : Span4Mux_h
    port map (
            O => \N__17431\,
            I => \N__17428\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__17428\,
            I => \c0.data_in_frame_6_Z0Z_0\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__17425\,
            I => \N__17422\
        );

    \I__3843\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17419\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17419\,
            I => \N__17416\
        );

    \I__3841\ : Odrv12
    port map (
            O => \N__17416\,
            I => \c0.data_in_frame_7_Z0Z_0\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__17413\,
            I => \c0.tx2.N_493_cascade_\
        );

    \I__3839\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17407\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__17407\,
            I => \c0.tx2.N_205_mux\
        );

    \I__3837\ : IoInMux
    port map (
            O => \N__17404\,
            I => \N__17401\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__17401\,
            I => \N__17398\
        );

    \I__3835\ : IoSpan4Mux
    port map (
            O => \N__17398\,
            I => \N__17395\
        );

    \I__3834\ : Span4Mux_s1_h
    port map (
            O => \N__17395\,
            I => \N__17392\
        );

    \I__3833\ : Sp12to4
    port map (
            O => \N__17392\,
            I => \N__17388\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__17391\,
            I => \N__17385\
        );

    \I__3831\ : Span12Mux_h
    port map (
            O => \N__17388\,
            I => \N__17382\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17379\
        );

    \I__3829\ : Odrv12
    port map (
            O => \N__17382\,
            I => \PIN_3_c\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__17379\,
            I => \PIN_3_c\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17371\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__17371\,
            I => \N__17366\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__17370\,
            I => \N__17363\
        );

    \I__3824\ : InMux
    port map (
            O => \N__17369\,
            I => \N__17360\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__17366\,
            I => \N__17357\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17363\,
            I => \N__17354\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__17360\,
            I => \N__17351\
        );

    \I__3820\ : Sp12to4
    port map (
            O => \N__17357\,
            I => \N__17346\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__17354\,
            I => \N__17346\
        );

    \I__3818\ : Odrv12
    port map (
            O => \N__17351\,
            I => \c0.data_in_7_Z0Z_0\
        );

    \I__3817\ : Odrv12
    port map (
            O => \N__17346\,
            I => \c0.data_in_7_Z0Z_0\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17341\,
            I => \N__17338\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__17338\,
            I => \N__17334\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17337\,
            I => \N__17330\
        );

    \I__3813\ : Span4Mux_v
    port map (
            O => \N__17334\,
            I => \N__17327\
        );

    \I__3812\ : InMux
    port map (
            O => \N__17333\,
            I => \N__17324\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17330\,
            I => \N__17321\
        );

    \I__3810\ : Sp12to4
    port map (
            O => \N__17327\,
            I => \N__17316\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__17324\,
            I => \N__17316\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__17321\,
            I => \c0.data_in_7_Z0Z_1\
        );

    \I__3807\ : Odrv12
    port map (
            O => \N__17316\,
            I => \c0.data_in_7_Z0Z_1\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17308\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17308\,
            I => \N__17305\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__17305\,
            I => \N__17302\
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__17302\,
            I => \c0.data_in_frame_7_Z0Z_1\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17296\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__17296\,
            I => \N__17293\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__17293\,
            I => \N__17288\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17285\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17291\,
            I => \N__17282\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__17288\,
            I => \c0.data_in_6_Z0Z_5\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__17285\,
            I => \c0.data_in_6_Z0Z_5\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__17282\,
            I => \c0.data_in_6_Z0Z_5\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__17275\,
            I => \N__17272\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17267\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17271\,
            I => \N__17264\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17261\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__17267\,
            I => \N__17258\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__17264\,
            I => \c0.data_in_7_Z0Z_5\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17261\,
            I => \c0.data_in_7_Z0Z_5\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__17258\,
            I => \c0.data_in_7_Z0Z_5\
        );

    \I__3786\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17248\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17248\,
            I => \N__17243\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17247\,
            I => \N__17240\
        );

    \I__3783\ : InMux
    port map (
            O => \N__17246\,
            I => \N__17237\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__17243\,
            I => \N__17234\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__17240\,
            I => \c0.data_in_7_Z0Z_6\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__17237\,
            I => \c0.data_in_7_Z0Z_6\
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__17234\,
            I => \c0.data_in_7_Z0Z_6\
        );

    \I__3778\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17224\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__17224\,
            I => \c0.data_in_frame_7_Z0Z_6\
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__17221\,
            I => \N__17218\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17218\,
            I => \N__17213\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17210\
        );

    \I__3773\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17207\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17204\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17210\,
            I => \c0.data_in_6_Z0Z_6\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__17207\,
            I => \c0.data_in_6_Z0Z_6\
        );

    \I__3769\ : Odrv12
    port map (
            O => \N__17204\,
            I => \c0.data_in_6_Z0Z_6\
        );

    \I__3768\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17194\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__17194\,
            I => \N__17191\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__17191\,
            I => \c0.data_in_frame_6_Z0Z_6\
        );

    \I__3765\ : CEMux
    port map (
            O => \N__17188\,
            I => \N__17131\
        );

    \I__3764\ : CEMux
    port map (
            O => \N__17187\,
            I => \N__17131\
        );

    \I__3763\ : CEMux
    port map (
            O => \N__17186\,
            I => \N__17131\
        );

    \I__3762\ : CEMux
    port map (
            O => \N__17185\,
            I => \N__17131\
        );

    \I__3761\ : CEMux
    port map (
            O => \N__17184\,
            I => \N__17131\
        );

    \I__3760\ : CEMux
    port map (
            O => \N__17183\,
            I => \N__17131\
        );

    \I__3759\ : CEMux
    port map (
            O => \N__17182\,
            I => \N__17131\
        );

    \I__3758\ : CEMux
    port map (
            O => \N__17181\,
            I => \N__17131\
        );

    \I__3757\ : CEMux
    port map (
            O => \N__17180\,
            I => \N__17131\
        );

    \I__3756\ : CEMux
    port map (
            O => \N__17179\,
            I => \N__17131\
        );

    \I__3755\ : CEMux
    port map (
            O => \N__17178\,
            I => \N__17131\
        );

    \I__3754\ : CEMux
    port map (
            O => \N__17177\,
            I => \N__17131\
        );

    \I__3753\ : CEMux
    port map (
            O => \N__17176\,
            I => \N__17131\
        );

    \I__3752\ : CEMux
    port map (
            O => \N__17175\,
            I => \N__17131\
        );

    \I__3751\ : CEMux
    port map (
            O => \N__17174\,
            I => \N__17131\
        );

    \I__3750\ : CEMux
    port map (
            O => \N__17173\,
            I => \N__17131\
        );

    \I__3749\ : CEMux
    port map (
            O => \N__17172\,
            I => \N__17131\
        );

    \I__3748\ : CEMux
    port map (
            O => \N__17171\,
            I => \N__17131\
        );

    \I__3747\ : CEMux
    port map (
            O => \N__17170\,
            I => \N__17131\
        );

    \I__3746\ : GlobalMux
    port map (
            O => \N__17131\,
            I => \N__17128\
        );

    \I__3745\ : gio2CtrlBuf
    port map (
            O => \N__17128\,
            I => \c0.data_in_frame_0__0_sqmuxa_g\
        );

    \I__3744\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17122\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__17122\,
            I => \c0.tx2.r_Clock_Count_i_3\
        );

    \I__3742\ : InMux
    port map (
            O => \N__17119\,
            I => \c0.tx2.r_Clock_Count12\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__17116\,
            I => \N__17109\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__17115\,
            I => \N__17106\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__17114\,
            I => \N__17100\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__17113\,
            I => \N__17097\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__17112\,
            I => \N__17094\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17109\,
            I => \N__17076\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17106\,
            I => \N__17076\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17076\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17076\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17071\
        );

    \I__3731\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17068\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17061\
        );

    \I__3729\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17061\
        );

    \I__3728\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17061\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__17092\,
            I => \N__17057\
        );

    \I__3726\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17053\
        );

    \I__3725\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17040\
        );

    \I__3724\ : InMux
    port map (
            O => \N__17089\,
            I => \N__17040\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17088\,
            I => \N__17040\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17040\
        );

    \I__3721\ : InMux
    port map (
            O => \N__17086\,
            I => \N__17040\
        );

    \I__3720\ : InMux
    port map (
            O => \N__17085\,
            I => \N__17040\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17076\,
            I => \N__17037\
        );

    \I__3718\ : InMux
    port map (
            O => \N__17075\,
            I => \N__17032\
        );

    \I__3717\ : InMux
    port map (
            O => \N__17074\,
            I => \N__17032\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__17071\,
            I => \N__17029\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__17068\,
            I => \N__17024\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__17061\,
            I => \N__17024\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17060\,
            I => \N__17021\
        );

    \I__3712\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17015\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17056\,
            I => \N__17012\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17053\,
            I => \N__17001\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__17040\,
            I => \N__17001\
        );

    \I__3708\ : Span4Mux_v
    port map (
            O => \N__17037\,
            I => \N__16996\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__17032\,
            I => \N__16996\
        );

    \I__3706\ : Span4Mux_h
    port map (
            O => \N__17029\,
            I => \N__16991\
        );

    \I__3705\ : Span4Mux_v
    port map (
            O => \N__17024\,
            I => \N__16991\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__17021\,
            I => \N__16988\
        );

    \I__3703\ : InMux
    port map (
            O => \N__17020\,
            I => \N__16981\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17019\,
            I => \N__16981\
        );

    \I__3701\ : InMux
    port map (
            O => \N__17018\,
            I => \N__16981\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17015\,
            I => \N__16976\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__17012\,
            I => \N__16976\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17011\,
            I => \N__16967\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17010\,
            I => \N__16967\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17009\,
            I => \N__16967\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17008\,
            I => \N__16967\
        );

    \I__3694\ : InMux
    port map (
            O => \N__17007\,
            I => \N__16962\
        );

    \I__3693\ : InMux
    port map (
            O => \N__17006\,
            I => \N__16962\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__17001\,
            I => \N__16952\
        );

    \I__3691\ : Span4Mux_h
    port map (
            O => \N__16996\,
            I => \N__16949\
        );

    \I__3690\ : Span4Mux_h
    port map (
            O => \N__16991\,
            I => \N__16942\
        );

    \I__3689\ : Span4Mux_h
    port map (
            O => \N__16988\,
            I => \N__16942\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__16981\,
            I => \N__16942\
        );

    \I__3687\ : Span12Mux_v
    port map (
            O => \N__16976\,
            I => \N__16935\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__16967\,
            I => \N__16935\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__16962\,
            I => \N__16935\
        );

    \I__3684\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16920\
        );

    \I__3683\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16920\
        );

    \I__3682\ : InMux
    port map (
            O => \N__16959\,
            I => \N__16920\
        );

    \I__3681\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16920\
        );

    \I__3680\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16920\
        );

    \I__3679\ : InMux
    port map (
            O => \N__16956\,
            I => \N__16920\
        );

    \I__3678\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16920\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__16952\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__16949\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__16942\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3674\ : Odrv12
    port map (
            O => \N__16935\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__16920\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3672\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16906\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__16906\,
            I => \N__16902\
        );

    \I__3670\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16899\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__16902\,
            I => \N__16896\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__16899\,
            I => \N__16893\
        );

    \I__3667\ : Span4Mux_h
    port map (
            O => \N__16896\,
            I => \N__16890\
        );

    \I__3666\ : Span4Mux_h
    port map (
            O => \N__16893\,
            I => \N__16887\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__16890\,
            I => \c0.d_2_29\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__16887\,
            I => \c0.d_2_29\
        );

    \I__3663\ : SRMux
    port map (
            O => \N__16882\,
            I => \N__16869\
        );

    \I__3662\ : SRMux
    port map (
            O => \N__16881\,
            I => \N__16866\
        );

    \I__3661\ : SRMux
    port map (
            O => \N__16880\,
            I => \N__16863\
        );

    \I__3660\ : SRMux
    port map (
            O => \N__16879\,
            I => \N__16860\
        );

    \I__3659\ : SRMux
    port map (
            O => \N__16878\,
            I => \N__16857\
        );

    \I__3658\ : SRMux
    port map (
            O => \N__16877\,
            I => \N__16854\
        );

    \I__3657\ : SRMux
    port map (
            O => \N__16876\,
            I => \N__16851\
        );

    \I__3656\ : SRMux
    port map (
            O => \N__16875\,
            I => \N__16848\
        );

    \I__3655\ : SRMux
    port map (
            O => \N__16874\,
            I => \N__16845\
        );

    \I__3654\ : SRMux
    port map (
            O => \N__16873\,
            I => \N__16842\
        );

    \I__3653\ : SRMux
    port map (
            O => \N__16872\,
            I => \N__16839\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__16869\,
            I => \N__16821\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__16866\,
            I => \N__16818\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__16863\,
            I => \N__16815\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__16860\,
            I => \N__16812\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__16857\,
            I => \N__16809\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__16854\,
            I => \N__16806\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__16851\,
            I => \N__16803\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__16848\,
            I => \N__16800\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__16845\,
            I => \N__16797\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__16842\,
            I => \N__16794\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__16839\,
            I => \N__16791\
        );

    \I__3641\ : CEMux
    port map (
            O => \N__16838\,
            I => \N__16738\
        );

    \I__3640\ : CEMux
    port map (
            O => \N__16837\,
            I => \N__16738\
        );

    \I__3639\ : CEMux
    port map (
            O => \N__16836\,
            I => \N__16738\
        );

    \I__3638\ : CEMux
    port map (
            O => \N__16835\,
            I => \N__16738\
        );

    \I__3637\ : CEMux
    port map (
            O => \N__16834\,
            I => \N__16738\
        );

    \I__3636\ : CEMux
    port map (
            O => \N__16833\,
            I => \N__16738\
        );

    \I__3635\ : CEMux
    port map (
            O => \N__16832\,
            I => \N__16738\
        );

    \I__3634\ : CEMux
    port map (
            O => \N__16831\,
            I => \N__16738\
        );

    \I__3633\ : CEMux
    port map (
            O => \N__16830\,
            I => \N__16738\
        );

    \I__3632\ : CEMux
    port map (
            O => \N__16829\,
            I => \N__16738\
        );

    \I__3631\ : CEMux
    port map (
            O => \N__16828\,
            I => \N__16738\
        );

    \I__3630\ : CEMux
    port map (
            O => \N__16827\,
            I => \N__16738\
        );

    \I__3629\ : CEMux
    port map (
            O => \N__16826\,
            I => \N__16738\
        );

    \I__3628\ : CEMux
    port map (
            O => \N__16825\,
            I => \N__16738\
        );

    \I__3627\ : CEMux
    port map (
            O => \N__16824\,
            I => \N__16738\
        );

    \I__3626\ : Glb2LocalMux
    port map (
            O => \N__16821\,
            I => \N__16738\
        );

    \I__3625\ : Glb2LocalMux
    port map (
            O => \N__16818\,
            I => \N__16738\
        );

    \I__3624\ : Glb2LocalMux
    port map (
            O => \N__16815\,
            I => \N__16738\
        );

    \I__3623\ : Glb2LocalMux
    port map (
            O => \N__16812\,
            I => \N__16738\
        );

    \I__3622\ : Glb2LocalMux
    port map (
            O => \N__16809\,
            I => \N__16738\
        );

    \I__3621\ : Glb2LocalMux
    port map (
            O => \N__16806\,
            I => \N__16738\
        );

    \I__3620\ : Glb2LocalMux
    port map (
            O => \N__16803\,
            I => \N__16738\
        );

    \I__3619\ : Glb2LocalMux
    port map (
            O => \N__16800\,
            I => \N__16738\
        );

    \I__3618\ : Glb2LocalMux
    port map (
            O => \N__16797\,
            I => \N__16738\
        );

    \I__3617\ : Glb2LocalMux
    port map (
            O => \N__16794\,
            I => \N__16738\
        );

    \I__3616\ : Glb2LocalMux
    port map (
            O => \N__16791\,
            I => \N__16738\
        );

    \I__3615\ : GlobalMux
    port map (
            O => \N__16738\,
            I => \N__16735\
        );

    \I__3614\ : gio2CtrlBuf
    port map (
            O => \N__16735\,
            I => \c0.data_out_0__1_sqmuxa_g\
        );

    \I__3613\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16729\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__16729\,
            I => \N__16726\
        );

    \I__3611\ : Span4Mux_v
    port map (
            O => \N__16726\,
            I => \N__16723\
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__16723\,
            I => \c0.tx2.r_Tx_DataZ0Z_6\
        );

    \I__3609\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16717\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__16717\,
            I => \N__16714\
        );

    \I__3607\ : Span4Mux_h
    port map (
            O => \N__16714\,
            I => \N__16711\
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__16711\,
            I => \c0.tx2.r_Tx_DataZ0Z_2\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__16708\,
            I => \c0.tx2.o_Tx_Serial_RNOZ0Z_6_cascade_\
        );

    \I__3604\ : InMux
    port map (
            O => \N__16705\,
            I => \N__16702\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__16702\,
            I => \N__16699\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__16699\,
            I => \c0.tx2.o_Tx_Serial_RNOZ0Z_5\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16696\,
            I => \N__16693\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__16693\,
            I => \c0.tx2.o_Tx_Serial_RNOZ0Z_3\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__16690\,
            I => \c0.tx2.m195_ns_1_cascade_\
        );

    \I__3598\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16684\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__16684\,
            I => \N__16681\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__16681\,
            I => \c0.tx2.o_Tx_Serial_RNOZ0Z_2\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__16678\,
            I => \c0.tx2.N_196_0_cascade_\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__16675\,
            I => \N__16671\
        );

    \I__3593\ : InMux
    port map (
            O => \N__16674\,
            I => \N__16667\
        );

    \I__3592\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16664\
        );

    \I__3591\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16661\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__16667\,
            I => \N__16656\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__16664\,
            I => \N__16656\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__16661\,
            I => \c0.d_4_1\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__16656\,
            I => \c0.d_4_1\
        );

    \I__3586\ : InMux
    port map (
            O => \N__16651\,
            I => \N__16648\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__16648\,
            I => \N__16643\
        );

    \I__3584\ : InMux
    port map (
            O => \N__16647\,
            I => \N__16638\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16638\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__16643\,
            I => \c0.d_4_9\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16638\,
            I => \c0.d_4_9\
        );

    \I__3580\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16630\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__16630\,
            I => \N__16627\
        );

    \I__3578\ : Odrv12
    port map (
            O => \N__16627\,
            I => \c0.tx2_data_RNO_3Z0Z_1\
        );

    \I__3577\ : InMux
    port map (
            O => \N__16624\,
            I => \N__16621\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__16621\,
            I => \N__16618\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__16618\,
            I => \c0.tx2.r_Tx_DataZ0Z_1\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__16615\,
            I => \N__16612\
        );

    \I__3573\ : InMux
    port map (
            O => \N__16612\,
            I => \N__16609\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__16609\,
            I => \N__16606\
        );

    \I__3571\ : Span4Mux_h
    port map (
            O => \N__16606\,
            I => \N__16603\
        );

    \I__3570\ : Span4Mux_h
    port map (
            O => \N__16603\,
            I => \N__16600\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__16600\,
            I => \c0.data_in_frame_6_Z0Z_1\
        );

    \I__3568\ : InMux
    port map (
            O => \N__16597\,
            I => \N__16594\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__16594\,
            I => \N__16591\
        );

    \I__3566\ : Odrv12
    port map (
            O => \N__16591\,
            I => \c0.tx2_data_RNO_1Z0Z_1\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16585\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__16585\,
            I => \N__16582\
        );

    \I__3563\ : Odrv12
    port map (
            O => \N__16582\,
            I => \c0.tx2.r_Tx_DataZ0Z_4\
        );

    \I__3562\ : InMux
    port map (
            O => \N__16579\,
            I => \N__16576\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__16576\,
            I => \N__16573\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__16573\,
            I => \c0.N_173_0\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16566\
        );

    \I__3558\ : InMux
    port map (
            O => \N__16569\,
            I => \N__16563\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__16566\,
            I => \c0.tx2.r_Clock_Count_i_0\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__16563\,
            I => \c0.tx2.r_Clock_Count_i_0\
        );

    \I__3555\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16555\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__16555\,
            I => \c0.tx2.r_Clock_Count_i_1\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16549\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__16549\,
            I => \c0.tx2.r_Clock_Count_i_2\
        );

    \I__3551\ : InMux
    port map (
            O => \N__16546\,
            I => \N__16539\
        );

    \I__3550\ : InMux
    port map (
            O => \N__16545\,
            I => \N__16539\
        );

    \I__3549\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16536\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__16539\,
            I => \N__16533\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__16536\,
            I => \N__16529\
        );

    \I__3546\ : Span4Mux_h
    port map (
            O => \N__16533\,
            I => \N__16526\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16532\,
            I => \N__16523\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__16529\,
            I => \c0.N_123\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__16526\,
            I => \c0.N_123\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__16523\,
            I => \c0.N_123\
        );

    \I__3541\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16512\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16509\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__16512\,
            I => \N__16506\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__16509\,
            I => \N__16502\
        );

    \I__3537\ : Span4Mux_v
    port map (
            O => \N__16506\,
            I => \N__16498\
        );

    \I__3536\ : InMux
    port map (
            O => \N__16505\,
            I => \N__16495\
        );

    \I__3535\ : Span4Mux_h
    port map (
            O => \N__16502\,
            I => \N__16492\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16489\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__16498\,
            I => \c0.d_4_15\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16495\,
            I => \c0.d_4_15\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__16492\,
            I => \c0.d_4_15\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16489\,
            I => \c0.d_4_15\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16480\,
            I => \N__16477\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__16477\,
            I => \c0.N_129\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__16474\,
            I => \N__16470\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16467\
        );

    \I__3525\ : InMux
    port map (
            O => \N__16470\,
            I => \N__16464\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__16467\,
            I => \c0.N_18\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__16464\,
            I => \c0.N_18\
        );

    \I__3522\ : InMux
    port map (
            O => \N__16459\,
            I => \c0.un1_byte_transmit_counter2_1_cry_0\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16456\,
            I => \c0.un1_byte_transmit_counter2_1_cry_1\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16453\,
            I => \c0.un1_byte_transmit_counter2_1_cry_2\
        );

    \I__3519\ : InMux
    port map (
            O => \N__16450\,
            I => \c0.un1_byte_transmit_counter2_1_cry_3\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16447\,
            I => \c0.un1_byte_transmit_counter2_1_cry_4\
        );

    \I__3517\ : InMux
    port map (
            O => \N__16444\,
            I => \c0.un1_byte_transmit_counter2_1_cry_5\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16441\,
            I => \c0.un1_byte_transmit_counter2_1_cry_6\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__16438\,
            I => \N__16431\
        );

    \I__3514\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16428\
        );

    \I__3513\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16423\
        );

    \I__3512\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16423\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16420\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16431\,
            I => \N__16417\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__16428\,
            I => \N__16414\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__16423\,
            I => \c0.d_4_38\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__16420\,
            I => \c0.d_4_38\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__16417\,
            I => \c0.d_4_38\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__16414\,
            I => \c0.d_4_38\
        );

    \I__3504\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16400\
        );

    \I__3503\ : InMux
    port map (
            O => \N__16404\,
            I => \N__16397\
        );

    \I__3502\ : InMux
    port map (
            O => \N__16403\,
            I => \N__16394\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__16400\,
            I => \N__16391\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__16397\,
            I => \c0.N_107\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__16394\,
            I => \c0.N_107\
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__16391\,
            I => \c0.N_107\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__16384\,
            I => \c0.un1_data_in_6__2_0_a2_6_a2_2_cascade_\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16378\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__16378\,
            I => \N__16375\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__16375\,
            I => \c0.un1_data_in_6__2\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__16372\,
            I => \N__16368\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__16371\,
            I => \N__16364\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16361\
        );

    \I__3490\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16358\
        );

    \I__3489\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16355\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__16361\,
            I => \N__16350\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__16358\,
            I => \N__16350\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__16355\,
            I => \N__16347\
        );

    \I__3485\ : Span4Mux_v
    port map (
            O => \N__16350\,
            I => \N__16344\
        );

    \I__3484\ : Span4Mux_v
    port map (
            O => \N__16347\,
            I => \N__16341\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__16344\,
            I => \c0.d_4_46\
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__16341\,
            I => \c0.d_4_46\
        );

    \I__3481\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16332\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16329\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__16332\,
            I => \N__16324\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__16329\,
            I => \N__16321\
        );

    \I__3477\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16318\
        );

    \I__3476\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16315\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__16324\,
            I => \c0.d_4_42\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__16321\,
            I => \c0.d_4_42\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__16318\,
            I => \c0.d_4_42\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__16315\,
            I => \c0.d_4_42\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16303\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__16303\,
            I => \N__16298\
        );

    \I__3469\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16295\
        );

    \I__3468\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16292\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__16298\,
            I => \c0.N_133\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__16295\,
            I => \c0.N_133\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__16292\,
            I => \c0.N_133\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__16285\,
            I => \c0.un1_data_in_7__2_0_a2_0_a2_5_cascade_\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16279\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__16279\,
            I => \N__16276\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__16276\,
            I => \c0.un1_data_in_7__2\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16269\
        );

    \I__3459\ : InMux
    port map (
            O => \N__16272\,
            I => \N__16265\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__16269\,
            I => \N__16262\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16259\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__16265\,
            I => \N__16256\
        );

    \I__3455\ : Span4Mux_v
    port map (
            O => \N__16262\,
            I => \N__16253\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__16259\,
            I => \c0.d_4_14\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__16256\,
            I => \c0.d_4_14\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__16253\,
            I => \c0.d_4_14\
        );

    \I__3451\ : InMux
    port map (
            O => \N__16246\,
            I => \N__16239\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16245\,
            I => \N__16236\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16244\,
            I => \N__16229\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16229\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16242\,
            I => \N__16229\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16239\,
            I => \c0.d_4_31\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16236\,
            I => \c0.d_4_31\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__16229\,
            I => \c0.d_4_31\
        );

    \I__3443\ : InMux
    port map (
            O => \N__16222\,
            I => \N__16219\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__16219\,
            I => \N__16216\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__16216\,
            I => \c0.un1_data_in_7__2_0_a2_0_a2_4\
        );

    \I__3440\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__16210\,
            I => \N__16207\
        );

    \I__3438\ : Span4Mux_v
    port map (
            O => \N__16207\,
            I => \N__16204\
        );

    \I__3437\ : Span4Mux_h
    port map (
            O => \N__16204\,
            I => \N__16201\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__16201\,
            I => \c0.un1_data_in_7__3_0_a2_0_a2_3\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16194\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16191\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__16194\,
            I => \N__16188\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16191\,
            I => \N__16185\
        );

    \I__3431\ : Span4Mux_v
    port map (
            O => \N__16188\,
            I => \N__16180\
        );

    \I__3430\ : Span4Mux_h
    port map (
            O => \N__16185\,
            I => \N__16177\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16174\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16171\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__16180\,
            I => \c0.d_4_43\
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__16177\,
            I => \c0.d_4_43\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__16174\,
            I => \c0.d_4_43\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__16171\,
            I => \c0.d_4_43\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16158\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16154\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16158\,
            I => \N__16151\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16148\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__16154\,
            I => \c0.N_128\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__16151\,
            I => \c0.N_128\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__16148\,
            I => \c0.N_128\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__16141\,
            I => \c0.un1_data_in_7__3_0_a2_0_a2_4_cascade_\
        );

    \I__3415\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16135\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__16135\,
            I => \c0.un1_data_in_7__5_0_a2_0_a2_1\
        );

    \I__3413\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16129\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16129\,
            I => \N__16126\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__16126\,
            I => \c0.m163_9\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16120\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__16120\,
            I => \N__16117\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__16117\,
            I => \N__16114\
        );

    \I__3407\ : Span4Mux_h
    port map (
            O => \N__16114\,
            I => \N__16110\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16107\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__16110\,
            I => \c0.data_in_0_Z0Z_1\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__16107\,
            I => \c0.data_in_0_Z0Z_1\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16099\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__16099\,
            I => \N__16095\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16098\,
            I => \N__16092\
        );

    \I__3400\ : Odrv12
    port map (
            O => \N__16095\,
            I => \c0.data_in_4_Z0Z_6\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16092\,
            I => \c0.data_in_4_Z0Z_6\
        );

    \I__3398\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16084\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__16084\,
            I => \N__16081\
        );

    \I__3396\ : Span4Mux_v
    port map (
            O => \N__16081\,
            I => \N__16077\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16074\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__16077\,
            I => \c0.data_in_5_Z0Z_6\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16074\,
            I => \c0.data_in_5_Z0Z_6\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16069\,
            I => \N__16065\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16068\,
            I => \N__16062\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__16065\,
            I => \N__16059\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__16062\,
            I => \N__16056\
        );

    \I__3388\ : Odrv12
    port map (
            O => \N__16059\,
            I => \c0.rx_data_6\
        );

    \I__3387\ : Odrv4
    port map (
            O => \N__16056\,
            I => \c0.rx_data_6\
        );

    \I__3386\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16047\
        );

    \I__3385\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16043\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__16047\,
            I => \N__16040\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16036\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16043\,
            I => \N__16033\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__16040\,
            I => \N__16030\
        );

    \I__3380\ : InMux
    port map (
            O => \N__16039\,
            I => \N__16027\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__16036\,
            I => \N__16024\
        );

    \I__3378\ : Odrv12
    port map (
            O => \N__16033\,
            I => \c0.d_4_26\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__16030\,
            I => \c0.d_4_26\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16027\,
            I => \c0.d_4_26\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__16024\,
            I => \c0.d_4_26\
        );

    \I__3374\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16012\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__16012\,
            I => \N__16007\
        );

    \I__3372\ : InMux
    port map (
            O => \N__16011\,
            I => \N__16004\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__16010\,
            I => \N__16001\
        );

    \I__3370\ : Span4Mux_h
    port map (
            O => \N__16007\,
            I => \N__15998\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__16004\,
            I => \N__15995\
        );

    \I__3368\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15992\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__15998\,
            I => \c0.data_in_6_Z0Z_4\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__15995\,
            I => \c0.data_in_6_Z0Z_4\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__15992\,
            I => \c0.data_in_6_Z0Z_4\
        );

    \I__3364\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15982\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__15982\,
            I => \N__15977\
        );

    \I__3362\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15974\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__15980\,
            I => \N__15971\
        );

    \I__3360\ : Span4Mux_v
    port map (
            O => \N__15977\,
            I => \N__15966\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15966\
        );

    \I__3358\ : InMux
    port map (
            O => \N__15971\,
            I => \N__15963\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__15966\,
            I => \N__15959\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__15963\,
            I => \N__15956\
        );

    \I__3355\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15953\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__15959\,
            I => \c0.d_4_41\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__15956\,
            I => \c0.d_4_41\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__15953\,
            I => \c0.d_4_41\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__15946\,
            I => \N__15943\
        );

    \I__3350\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15940\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__15940\,
            I => \c0.un1_data_in_6__4_0_a2_5_a2_1\
        );

    \I__3348\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15934\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__15934\,
            I => \N__15930\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__15933\,
            I => \N__15926\
        );

    \I__3345\ : Span4Mux_v
    port map (
            O => \N__15930\,
            I => \N__15923\
        );

    \I__3344\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15918\
        );

    \I__3343\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15918\
        );

    \I__3342\ : Span4Mux_h
    port map (
            O => \N__15923\,
            I => \N__15913\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__15918\,
            I => \N__15913\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__15913\,
            I => \c0.data_in_1_Z0Z_2\
        );

    \I__3339\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15907\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__15907\,
            I => \N__15902\
        );

    \I__3337\ : InMux
    port map (
            O => \N__15906\,
            I => \N__15897\
        );

    \I__3336\ : InMux
    port map (
            O => \N__15905\,
            I => \N__15897\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__15902\,
            I => \c0.d_4_10\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__15897\,
            I => \c0.d_4_10\
        );

    \I__3333\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15888\
        );

    \I__3332\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15885\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__15888\,
            I => \N__15882\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__15885\,
            I => \c0.N_127\
        );

    \I__3329\ : Odrv12
    port map (
            O => \N__15882\,
            I => \c0.N_127\
        );

    \I__3328\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15874\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__15874\,
            I => \N__15871\
        );

    \I__3326\ : Span12Mux_h
    port map (
            O => \N__15871\,
            I => \N__15866\
        );

    \I__3325\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15863\
        );

    \I__3324\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15860\
        );

    \I__3323\ : Odrv12
    port map (
            O => \N__15866\,
            I => \c0.data_in_1_Z0Z_1\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__15863\,
            I => \c0.data_in_1_Z0Z_1\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__15860\,
            I => \c0.data_in_1_Z0Z_1\
        );

    \I__3320\ : InMux
    port map (
            O => \N__15853\,
            I => \N__15850\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__15850\,
            I => \N__15846\
        );

    \I__3318\ : InMux
    port map (
            O => \N__15849\,
            I => \N__15843\
        );

    \I__3317\ : Span4Mux_h
    port map (
            O => \N__15846\,
            I => \N__15839\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__15843\,
            I => \N__15836\
        );

    \I__3315\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15833\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__15839\,
            I => \c0.data_in_3_Z0Z_1\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__15836\,
            I => \c0.data_in_3_Z0Z_1\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__15833\,
            I => \c0.data_in_3_Z0Z_1\
        );

    \I__3311\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15823\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__15823\,
            I => \N__15820\
        );

    \I__3309\ : Span4Mux_h
    port map (
            O => \N__15820\,
            I => \N__15815\
        );

    \I__3308\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15812\
        );

    \I__3307\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15809\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__15815\,
            I => \c0.d_4_25\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__15812\,
            I => \c0.d_4_25\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__15809\,
            I => \c0.d_4_25\
        );

    \I__3303\ : InMux
    port map (
            O => \N__15802\,
            I => \N__15799\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__15799\,
            I => \c0.data_in_frame_6_Z0Z_4\
        );

    \I__3301\ : InMux
    port map (
            O => \N__15796\,
            I => \N__15793\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__15793\,
            I => \c0.data_in_frame_7_Z0Z_4\
        );

    \I__3299\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15787\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__15787\,
            I => \c0.tx2_data_RNO_1Z0Z_4\
        );

    \I__3297\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15781\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__15781\,
            I => \c0.tx2_data_RNO_0Z0Z_4\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__15778\,
            I => \c0.m120_ns_1_cascade_\
        );

    \I__3294\ : InMux
    port map (
            O => \N__15775\,
            I => \N__15772\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__15772\,
            I => \c0.tx2_data_RNO_3Z0Z_6\
        );

    \I__3292\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15766\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__15766\,
            I => \c0.tx2_data_RNO_0Z0Z_6\
        );

    \I__3290\ : CascadeMux
    port map (
            O => \N__15763\,
            I => \c0.m90_ns_1_cascade_\
        );

    \I__3289\ : InMux
    port map (
            O => \N__15760\,
            I => \N__15757\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__15757\,
            I => \c0.tx2_data_RNO_1Z0Z_6\
        );

    \I__3287\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15751\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__15751\,
            I => \N__15747\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15750\,
            I => \N__15743\
        );

    \I__3284\ : Span4Mux_h
    port map (
            O => \N__15747\,
            I => \N__15740\
        );

    \I__3283\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15737\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__15743\,
            I => \N__15734\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__15740\,
            I => \c0.data_in_7_Z0Z_4\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__15737\,
            I => \c0.data_in_7_Z0Z_4\
        );

    \I__3279\ : Odrv12
    port map (
            O => \N__15734\,
            I => \c0.data_in_7_Z0Z_4\
        );

    \I__3278\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15724\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__15724\,
            I => \N__15721\
        );

    \I__3276\ : Span4Mux_h
    port map (
            O => \N__15721\,
            I => \N__15718\
        );

    \I__3275\ : Span4Mux_h
    port map (
            O => \N__15718\,
            I => \N__15714\
        );

    \I__3274\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15711\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__15714\,
            I => \c0.rx_data_5\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__15711\,
            I => \c0.rx_data_5\
        );

    \I__3271\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15699\
        );

    \I__3270\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15699\
        );

    \I__3269\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15696\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__15699\,
            I => \N__15693\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__15696\,
            I => \N__15690\
        );

    \I__3266\ : Span4Mux_h
    port map (
            O => \N__15693\,
            I => \N__15687\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__15690\,
            I => \c0.d_2_10\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__15687\,
            I => \c0.d_2_10\
        );

    \I__3263\ : InMux
    port map (
            O => \N__15682\,
            I => \N__15679\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__15679\,
            I => \c0.byte_transmit_counterZ0Z_6\
        );

    \I__3261\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15673\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15673\,
            I => \c0.byte_transmit_counterZ0Z_7\
        );

    \I__3259\ : InMux
    port map (
            O => \N__15670\,
            I => \N__15667\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__15667\,
            I => \c0.byte_transmit_counterZ0Z_3\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15664\,
            I => \N__15661\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__15661\,
            I => \c0.byte_transmit_counterZ0Z_4\
        );

    \I__3255\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15653\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15647\
        );

    \I__3253\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15644\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__15653\,
            I => \N__15641\
        );

    \I__3251\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15637\
        );

    \I__3250\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15634\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15650\,
            I => \N__15628\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__15647\,
            I => \N__15625\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15644\,
            I => \N__15622\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__15641\,
            I => \N__15619\
        );

    \I__3245\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15616\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__15637\,
            I => \N__15611\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15611\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15607\
        );

    \I__3241\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15604\
        );

    \I__3240\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15601\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__15628\,
            I => \N__15596\
        );

    \I__3238\ : Span4Mux_h
    port map (
            O => \N__15625\,
            I => \N__15596\
        );

    \I__3237\ : Span4Mux_h
    port map (
            O => \N__15622\,
            I => \N__15593\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__15619\,
            I => \N__15586\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__15616\,
            I => \N__15586\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__15611\,
            I => \N__15586\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15583\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__15607\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__15604\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__15601\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__15596\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__15593\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__15586\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__15583\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__15568\,
            I => \N__15562\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__15567\,
            I => \N__15559\
        );

    \I__3223\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15550\
        );

    \I__3222\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15550\
        );

    \I__3221\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15541\
        );

    \I__3220\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15541\
        );

    \I__3219\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15541\
        );

    \I__3218\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15541\
        );

    \I__3217\ : InMux
    port map (
            O => \N__15556\,
            I => \N__15523\
        );

    \I__3216\ : InMux
    port map (
            O => \N__15555\,
            I => \N__15523\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__15550\,
            I => \N__15518\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15518\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__15540\,
            I => \N__15512\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__15539\,
            I => \N__15507\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__15538\,
            I => \N__15504\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15489\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15536\,
            I => \N__15489\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15535\,
            I => \N__15489\
        );

    \I__3207\ : InMux
    port map (
            O => \N__15534\,
            I => \N__15489\
        );

    \I__3206\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15489\
        );

    \I__3205\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15482\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15531\,
            I => \N__15482\
        );

    \I__3203\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15482\
        );

    \I__3202\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15479\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15475\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__15523\,
            I => \N__15466\
        );

    \I__3199\ : Span4Mux_h
    port map (
            O => \N__15518\,
            I => \N__15466\
        );

    \I__3198\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15463\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15516\,
            I => \N__15460\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15515\,
            I => \N__15451\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15451\
        );

    \I__3194\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15451\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15510\,
            I => \N__15451\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15507\,
            I => \N__15438\
        );

    \I__3191\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15438\
        );

    \I__3190\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15438\
        );

    \I__3189\ : InMux
    port map (
            O => \N__15502\,
            I => \N__15438\
        );

    \I__3188\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15438\
        );

    \I__3187\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15438\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__15489\,
            I => \N__15435\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__15482\,
            I => \N__15430\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__15479\,
            I => \N__15430\
        );

    \I__3183\ : InMux
    port map (
            O => \N__15478\,
            I => \N__15426\
        );

    \I__3182\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15421\
        );

    \I__3181\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15421\
        );

    \I__3180\ : InMux
    port map (
            O => \N__15473\,
            I => \N__15416\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15472\,
            I => \N__15416\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15413\
        );

    \I__3177\ : Span4Mux_v
    port map (
            O => \N__15466\,
            I => \N__15410\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__15463\,
            I => \N__15397\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__15460\,
            I => \N__15397\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__15451\,
            I => \N__15397\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__15438\,
            I => \N__15397\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__15435\,
            I => \N__15397\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__15430\,
            I => \N__15397\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15394\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15426\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__15421\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__15416\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__15413\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__15410\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__15397\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__15394\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15379\,
            I => \N__15376\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__15376\,
            I => \N__15361\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15356\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15356\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15347\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15372\,
            I => \N__15347\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15347\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15370\,
            I => \N__15347\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15369\,
            I => \N__15321\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15368\,
            I => \N__15321\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15367\,
            I => \N__15321\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15366\,
            I => \N__15321\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15321\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15364\,
            I => \N__15318\
        );

    \I__3148\ : Span4Mux_v
    port map (
            O => \N__15361\,
            I => \N__15311\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15356\,
            I => \N__15311\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15347\,
            I => \N__15311\
        );

    \I__3145\ : InMux
    port map (
            O => \N__15346\,
            I => \N__15304\
        );

    \I__3144\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15304\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15344\,
            I => \N__15304\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15295\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15342\,
            I => \N__15295\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15295\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15295\
        );

    \I__3138\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15290\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15338\,
            I => \N__15290\
        );

    \I__3136\ : InMux
    port map (
            O => \N__15337\,
            I => \N__15279\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15274\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15274\
        );

    \I__3133\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15271\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15268\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15265\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__15321\,
            I => \N__15262\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15251\
        );

    \I__3128\ : Span4Mux_h
    port map (
            O => \N__15311\,
            I => \N__15251\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__15304\,
            I => \N__15251\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__15295\,
            I => \N__15251\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__15290\,
            I => \N__15251\
        );

    \I__3124\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15238\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15238\
        );

    \I__3122\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15238\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15238\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15285\,
            I => \N__15238\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15284\,
            I => \N__15238\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15233\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15233\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__15279\,
            I => \c0.N_132_mux\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__15274\,
            I => \c0.N_132_mux\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__15271\,
            I => \c0.N_132_mux\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__15268\,
            I => \c0.N_132_mux\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__15265\,
            I => \c0.N_132_mux\
        );

    \I__3111\ : Odrv12
    port map (
            O => \N__15262\,
            I => \c0.N_132_mux\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__15251\,
            I => \c0.N_132_mux\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15238\,
            I => \c0.N_132_mux\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__15233\,
            I => \c0.N_132_mux\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__15214\,
            I => \N__15206\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__15213\,
            I => \N__15203\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__15212\,
            I => \N__15200\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__15211\,
            I => \N__15194\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__15210\,
            I => \N__15191\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \N__15188\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15183\
        );

    \I__3100\ : InMux
    port map (
            O => \N__15203\,
            I => \N__15174\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15174\
        );

    \I__3098\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15174\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15174\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15171\
        );

    \I__3095\ : InMux
    port map (
            O => \N__15194\,
            I => \N__15168\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15156\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15156\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15156\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15186\,
            I => \N__15153\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__15183\,
            I => \N__15146\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__15174\,
            I => \N__15146\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__15171\,
            I => \N__15146\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15168\,
            I => \N__15143\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15140\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15137\
        );

    \I__3084\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15134\
        );

    \I__3083\ : InMux
    port map (
            O => \N__15164\,
            I => \N__15130\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15127\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15156\,
            I => \N__15120\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__15153\,
            I => \N__15120\
        );

    \I__3079\ : Span4Mux_h
    port map (
            O => \N__15146\,
            I => \N__15120\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__15143\,
            I => \N__15111\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15140\,
            I => \N__15111\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__15137\,
            I => \N__15111\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__15134\,
            I => \N__15111\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15107\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15130\,
            I => \N__15102\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__15127\,
            I => \N__15102\
        );

    \I__3071\ : Span4Mux_v
    port map (
            O => \N__15120\,
            I => \N__15099\
        );

    \I__3070\ : Span4Mux_v
    port map (
            O => \N__15111\,
            I => \N__15096\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15093\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__15107\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__3067\ : Odrv12
    port map (
            O => \N__15102\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__15099\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__15096\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__15093\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__15082\,
            I => \c0.N_5_1_cascade_\
        );

    \I__3062\ : CEMux
    port map (
            O => \N__15079\,
            I => \N__15076\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__15076\,
            I => \N__15072\
        );

    \I__3060\ : CEMux
    port map (
            O => \N__15075\,
            I => \N__15069\
        );

    \I__3059\ : Span4Mux_h
    port map (
            O => \N__15072\,
            I => \N__15064\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__15069\,
            I => \N__15064\
        );

    \I__3057\ : Span4Mux_v
    port map (
            O => \N__15064\,
            I => \N__15060\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15057\
        );

    \I__3055\ : Sp12to4
    port map (
            O => \N__15060\,
            I => \N__15052\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__15057\,
            I => \N__15052\
        );

    \I__3053\ : Span12Mux_s11_v
    port map (
            O => \N__15052\,
            I => \N__15049\
        );

    \I__3052\ : Odrv12
    port map (
            O => \N__15049\,
            I => \c0.byte_transmit_counter15\
        );

    \I__3051\ : IoInMux
    port map (
            O => \N__15046\,
            I => \N__15043\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15043\,
            I => \N__15040\
        );

    \I__3049\ : Span4Mux_s0_v
    port map (
            O => \N__15040\,
            I => \N__15037\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__15034\,
            I => \c0.data_out_0__1_sqmuxa\
        );

    \I__3046\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15027\
        );

    \I__3045\ : InMux
    port map (
            O => \N__15030\,
            I => \N__15023\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__15027\,
            I => \N__15020\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__15026\,
            I => \N__15017\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15023\,
            I => \N__15014\
        );

    \I__3041\ : Span4Mux_h
    port map (
            O => \N__15020\,
            I => \N__15011\
        );

    \I__3040\ : InMux
    port map (
            O => \N__15017\,
            I => \N__15008\
        );

    \I__3039\ : Odrv12
    port map (
            O => \N__15014\,
            I => \c0.d_2_14\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__15011\,
            I => \c0.d_2_14\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__15008\,
            I => \c0.d_2_14\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__15001\,
            I => \N__14998\
        );

    \I__3035\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14994\
        );

    \I__3034\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14990\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__14994\,
            I => \N__14987\
        );

    \I__3032\ : InMux
    port map (
            O => \N__14993\,
            I => \N__14984\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__14990\,
            I => \N__14980\
        );

    \I__3030\ : Span4Mux_h
    port map (
            O => \N__14987\,
            I => \N__14977\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14974\
        );

    \I__3028\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14971\
        );

    \I__3027\ : Span4Mux_h
    port map (
            O => \N__14980\,
            I => \N__14968\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__14977\,
            I => \c0.d_2_30\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__14974\,
            I => \c0.d_2_30\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__14971\,
            I => \c0.d_2_30\
        );

    \I__3023\ : Odrv4
    port map (
            O => \N__14968\,
            I => \c0.d_2_30\
        );

    \I__3022\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14954\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14958\,
            I => \N__14949\
        );

    \I__3020\ : InMux
    port map (
            O => \N__14957\,
            I => \N__14949\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__14954\,
            I => \N__14946\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__14949\,
            I => \N__14941\
        );

    \I__3017\ : Span4Mux_v
    port map (
            O => \N__14946\,
            I => \N__14941\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__14941\,
            I => \c0.d_2_16\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__14938\,
            I => \N__14935\
        );

    \I__3014\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14930\
        );

    \I__3013\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14927\
        );

    \I__3012\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14923\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__14930\,
            I => \N__14920\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__14927\,
            I => \N__14917\
        );

    \I__3009\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14914\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14907\
        );

    \I__3007\ : Span4Mux_v
    port map (
            O => \N__14920\,
            I => \N__14907\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__14917\,
            I => \N__14907\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__14914\,
            I => \c0.d_2_17\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__14907\,
            I => \c0.d_2_17\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__14902\,
            I => \N__14899\
        );

    \I__3002\ : InMux
    port map (
            O => \N__14899\,
            I => \N__14896\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__14896\,
            I => \N__14891\
        );

    \I__3000\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14886\
        );

    \I__2999\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14886\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__14891\,
            I => \N__14883\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__14886\,
            I => \N__14880\
        );

    \I__2996\ : Odrv4
    port map (
            O => \N__14883\,
            I => \c0.d_2_12\
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__14880\,
            I => \c0.d_2_12\
        );

    \I__2994\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14870\
        );

    \I__2993\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14867\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__14873\,
            I => \N__14863\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__14870\,
            I => \N__14860\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__14867\,
            I => \N__14857\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__14866\,
            I => \N__14854\
        );

    \I__2988\ : InMux
    port map (
            O => \N__14863\,
            I => \N__14851\
        );

    \I__2987\ : Span12Mux_h
    port map (
            O => \N__14860\,
            I => \N__14848\
        );

    \I__2986\ : Span4Mux_v
    port map (
            O => \N__14857\,
            I => \N__14845\
        );

    \I__2985\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14842\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__14851\,
            I => \N__14839\
        );

    \I__2983\ : Odrv12
    port map (
            O => \N__14848\,
            I => \c0.d_2_21\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__14845\,
            I => \c0.d_2_21\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14842\,
            I => \c0.d_2_21\
        );

    \I__2980\ : Odrv12
    port map (
            O => \N__14839\,
            I => \c0.d_2_21\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__14830\,
            I => \N__14826\
        );

    \I__2978\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14823\
        );

    \I__2977\ : InMux
    port map (
            O => \N__14826\,
            I => \N__14820\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__14823\,
            I => \N__14815\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__14820\,
            I => \N__14812\
        );

    \I__2974\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14807\
        );

    \I__2973\ : InMux
    port map (
            O => \N__14818\,
            I => \N__14807\
        );

    \I__2972\ : Span4Mux_h
    port map (
            O => \N__14815\,
            I => \N__14804\
        );

    \I__2971\ : Span4Mux_v
    port map (
            O => \N__14812\,
            I => \N__14799\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__14807\,
            I => \N__14799\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__14804\,
            I => \c0.d_2_11\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__14799\,
            I => \c0.d_2_11\
        );

    \I__2967\ : InMux
    port map (
            O => \N__14794\,
            I => \N__14790\
        );

    \I__2966\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14786\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__14790\,
            I => \N__14783\
        );

    \I__2964\ : InMux
    port map (
            O => \N__14789\,
            I => \N__14780\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__14786\,
            I => \N__14777\
        );

    \I__2962\ : Span4Mux_h
    port map (
            O => \N__14783\,
            I => \N__14772\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__14780\,
            I => \N__14769\
        );

    \I__2960\ : Span4Mux_h
    port map (
            O => \N__14777\,
            I => \N__14766\
        );

    \I__2959\ : InMux
    port map (
            O => \N__14776\,
            I => \N__14763\
        );

    \I__2958\ : InMux
    port map (
            O => \N__14775\,
            I => \N__14760\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__14772\,
            I => \c0.d_2_26\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__14769\,
            I => \c0.d_2_26\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__14766\,
            I => \c0.d_2_26\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__14763\,
            I => \c0.d_2_26\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__14760\,
            I => \c0.d_2_26\
        );

    \I__2952\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14744\
        );

    \I__2951\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14738\
        );

    \I__2950\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14738\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__14744\,
            I => \N__14735\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__14743\,
            I => \N__14732\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__14738\,
            I => \N__14729\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__14735\,
            I => \N__14726\
        );

    \I__2945\ : InMux
    port map (
            O => \N__14732\,
            I => \N__14723\
        );

    \I__2944\ : Span4Mux_h
    port map (
            O => \N__14729\,
            I => \N__14720\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__14726\,
            I => \c0.d_2_18\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__14723\,
            I => \c0.d_2_18\
        );

    \I__2941\ : Odrv4
    port map (
            O => \N__14720\,
            I => \c0.d_2_18\
        );

    \I__2940\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14710\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__14710\,
            I => \N__14706\
        );

    \I__2938\ : InMux
    port map (
            O => \N__14709\,
            I => \N__14701\
        );

    \I__2937\ : Span4Mux_v
    port map (
            O => \N__14706\,
            I => \N__14697\
        );

    \I__2936\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14694\
        );

    \I__2935\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14691\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__14701\,
            I => \N__14688\
        );

    \I__2933\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14685\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__14697\,
            I => \c0.d_4_35\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__14694\,
            I => \c0.d_4_35\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14691\,
            I => \c0.d_4_35\
        );

    \I__2929\ : Odrv12
    port map (
            O => \N__14688\,
            I => \c0.d_4_35\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__14685\,
            I => \c0.d_4_35\
        );

    \I__2927\ : InMux
    port map (
            O => \N__14674\,
            I => \N__14671\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__14671\,
            I => \N__14668\
        );

    \I__2925\ : Span4Mux_v
    port map (
            O => \N__14668\,
            I => \N__14662\
        );

    \I__2924\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14657\
        );

    \I__2923\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14657\
        );

    \I__2922\ : InMux
    port map (
            O => \N__14665\,
            I => \N__14654\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__14662\,
            I => \c0.d_4_27\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__14657\,
            I => \c0.d_4_27\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__14654\,
            I => \c0.d_4_27\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__14647\,
            I => \N__14644\
        );

    \I__2917\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14641\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__14641\,
            I => \N__14637\
        );

    \I__2915\ : InMux
    port map (
            O => \N__14640\,
            I => \N__14634\
        );

    \I__2914\ : Span4Mux_v
    port map (
            O => \N__14637\,
            I => \N__14629\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__14634\,
            I => \N__14629\
        );

    \I__2912\ : Span4Mux_v
    port map (
            O => \N__14629\,
            I => \N__14625\
        );

    \I__2911\ : InMux
    port map (
            O => \N__14628\,
            I => \N__14622\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__14625\,
            I => \c0.d_4_19\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__14622\,
            I => \c0.d_4_19\
        );

    \I__2908\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14614\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14614\,
            I => \N__14608\
        );

    \I__2906\ : InMux
    port map (
            O => \N__14613\,
            I => \N__14603\
        );

    \I__2905\ : InMux
    port map (
            O => \N__14612\,
            I => \N__14603\
        );

    \I__2904\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14600\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__14608\,
            I => \c0.d_4_3\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__14603\,
            I => \c0.d_4_3\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__14600\,
            I => \c0.d_4_3\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__14593\,
            I => \N__14590\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14587\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14583\
        );

    \I__2897\ : InMux
    port map (
            O => \N__14586\,
            I => \N__14580\
        );

    \I__2896\ : Span4Mux_v
    port map (
            O => \N__14583\,
            I => \N__14574\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__14580\,
            I => \N__14574\
        );

    \I__2894\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14571\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__14574\,
            I => \c0.d_4_11\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__14571\,
            I => \c0.d_4_11\
        );

    \I__2891\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14563\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__14563\,
            I => \c0.tx2_data_RNO_4Z0Z_3\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__14560\,
            I => \c0.tx2_data_RNO_3Z0Z_3_cascade_\
        );

    \I__2888\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14554\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__14554\,
            I => \c0.tx2_data_RNO_0Z0Z_3\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__14551\,
            I => \c0.m105_ns_1_cascade_\
        );

    \I__2885\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14545\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__14545\,
            I => \N__14542\
        );

    \I__2883\ : Span4Mux_h
    port map (
            O => \N__14542\,
            I => \N__14539\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__14539\,
            I => \c0.tx2_data_RNO_1Z0Z_3\
        );

    \I__2881\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14533\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__14533\,
            I => \c0.tx2.r_Tx_DataZ0Z_3\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__14530\,
            I => \N__14527\
        );

    \I__2878\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14524\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__2876\ : Span4Mux_v
    port map (
            O => \N__14521\,
            I => \N__14518\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__14518\,
            I => \c0.tx2_data_RNO_1Z0Z_7\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14512\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__14512\,
            I => \c0.m60_0_ns_1\
        );

    \I__2872\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14506\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__14506\,
            I => \c0.tx2.r_Tx_DataZ0Z_7\
        );

    \I__2870\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14499\
        );

    \I__2869\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14494\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__14499\,
            I => \N__14491\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14488\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14485\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__14494\,
            I => \N__14482\
        );

    \I__2864\ : Span12Mux_v
    port map (
            O => \N__14491\,
            I => \N__14475\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14475\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__14485\,
            I => \N__14475\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__14482\,
            I => \c0.d_2_6\
        );

    \I__2860\ : Odrv12
    port map (
            O => \N__14475\,
            I => \c0.d_2_6\
        );

    \I__2859\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14467\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__14467\,
            I => \N__14461\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14456\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14456\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__14464\,
            I => \N__14453\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__14461\,
            I => \N__14448\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__14456\,
            I => \N__14448\
        );

    \I__2852\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14445\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__14448\,
            I => \N__14442\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__14445\,
            I => \c0.d_2_22\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__14442\,
            I => \c0.d_2_22\
        );

    \I__2848\ : InMux
    port map (
            O => \N__14437\,
            I => \N__14434\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__14434\,
            I => \N__14431\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__14431\,
            I => \N__14427\
        );

    \I__2845\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14424\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__14427\,
            I => \c0.data_in_0_Z0Z_2\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14424\,
            I => \c0.data_in_0_Z0Z_2\
        );

    \I__2842\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14416\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__14416\,
            I => \N__14413\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__14413\,
            I => \N__14410\
        );

    \I__2839\ : Span4Mux_v
    port map (
            O => \N__14410\,
            I => \N__14406\
        );

    \I__2838\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14403\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__14406\,
            I => \c0.data_in_4_Z0Z_0\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__14403\,
            I => \c0.data_in_4_Z0Z_0\
        );

    \I__2835\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14395\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__14395\,
            I => \N__14391\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__14394\,
            I => \N__14387\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__14391\,
            I => \N__14384\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14390\,
            I => \N__14379\
        );

    \I__2830\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14379\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__14384\,
            I => \c0.d_4_23\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__14379\,
            I => \c0.d_4_23\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__14374\,
            I => \N__14371\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14368\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14368\,
            I => \c0.tx2_data_RNO_4Z0Z_7\
        );

    \I__2824\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14362\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__14362\,
            I => \N__14357\
        );

    \I__2822\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14352\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14352\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__14357\,
            I => \c0.d_4_2\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__14352\,
            I => \c0.d_4_2\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14344\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__14344\,
            I => \N__14341\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__14341\,
            I => \c0.tx2_data_RNO_4Z0Z_2\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__14338\,
            I => \c0.tx2_data_RNO_3Z0Z_2_cascade_\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14332\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14332\,
            I => \N__14329\
        );

    \I__2812\ : Span4Mux_h
    port map (
            O => \N__14329\,
            I => \N__14326\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__14326\,
            I => \c0.m131_ns_1\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14323\,
            I => \N__14320\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__14320\,
            I => \N__14317\
        );

    \I__2808\ : Span4Mux_v
    port map (
            O => \N__14317\,
            I => \N__14314\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__14314\,
            I => \c0.tx_data_RNO_1Z0Z_6\
        );

    \I__2806\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14308\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14308\,
            I => \c0.tx_data_RNO_0Z0Z_6\
        );

    \I__2804\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14302\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__14302\,
            I => \c0.tx_data_1_0_i_ns_1_6\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14296\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__14296\,
            I => \N__14293\
        );

    \I__2800\ : Span4Mux_v
    port map (
            O => \N__14293\,
            I => \N__14290\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__14290\,
            I => \c0.tx.r_Tx_DataZ0Z_6\
        );

    \I__2798\ : CEMux
    port map (
            O => \N__14287\,
            I => \N__14284\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14280\
        );

    \I__2796\ : CEMux
    port map (
            O => \N__14283\,
            I => \N__14276\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__14280\,
            I => \N__14273\
        );

    \I__2794\ : CEMux
    port map (
            O => \N__14279\,
            I => \N__14270\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14276\,
            I => \N__14267\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__14273\,
            I => \N__14262\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14270\,
            I => \N__14262\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__14267\,
            I => \N__14259\
        );

    \I__2789\ : Span4Mux_h
    port map (
            O => \N__14262\,
            I => \N__14256\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__14259\,
            I => \c0.tx.N_398_i\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__14256\,
            I => \c0.tx.N_398_i\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__14251\,
            I => \N__14248\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14241\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14238\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__14246\,
            I => \N__14234\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14245\,
            I => \N__14228\
        );

    \I__2781\ : InMux
    port map (
            O => \N__14244\,
            I => \N__14228\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14222\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__14238\,
            I => \N__14222\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__14237\,
            I => \N__14218\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14212\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14212\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__14228\,
            I => \N__14209\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14227\,
            I => \N__14206\
        );

    \I__2773\ : Span12Mux_h
    port map (
            O => \N__14222\,
            I => \N__14203\
        );

    \I__2772\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14196\
        );

    \I__2771\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14196\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14196\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__14212\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__14209\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__14206\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__2766\ : Odrv12
    port map (
            O => \N__14203\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__14196\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14181\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14170\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__14181\,
            I => \N__14167\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14180\,
            I => \N__14164\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14161\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14158\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14153\
        );

    \I__2757\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14153\
        );

    \I__2756\ : InMux
    port map (
            O => \N__14175\,
            I => \N__14150\
        );

    \I__2755\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14145\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14145\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__14170\,
            I => \N__14140\
        );

    \I__2752\ : Span12Mux_h
    port map (
            O => \N__14167\,
            I => \N__14140\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14164\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__14161\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__14158\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__14153\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14150\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__14145\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__2745\ : Odrv12
    port map (
            O => \N__14140\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__2744\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14121\
        );

    \I__2743\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14118\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__14121\,
            I => \N__14113\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__14118\,
            I => \N__14106\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14100\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14097\
        );

    \I__2738\ : Span4Mux_v
    port map (
            O => \N__14113\,
            I => \N__14094\
        );

    \I__2737\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14091\
        );

    \I__2736\ : InMux
    port map (
            O => \N__14111\,
            I => \N__14086\
        );

    \I__2735\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14086\
        );

    \I__2734\ : InMux
    port map (
            O => \N__14109\,
            I => \N__14083\
        );

    \I__2733\ : Span12Mux_v
    port map (
            O => \N__14106\,
            I => \N__14080\
        );

    \I__2732\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14073\
        );

    \I__2731\ : InMux
    port map (
            O => \N__14104\,
            I => \N__14073\
        );

    \I__2730\ : InMux
    port map (
            O => \N__14103\,
            I => \N__14073\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__14100\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__14097\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__14094\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__14091\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__14086\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__14083\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__2723\ : Odrv12
    port map (
            O => \N__14080\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14073\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__2721\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14053\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__14053\,
            I => \N__14050\
        );

    \I__2719\ : Span4Mux_h
    port map (
            O => \N__14050\,
            I => \N__14046\
        );

    \I__2718\ : InMux
    port map (
            O => \N__14049\,
            I => \N__14043\
        );

    \I__2717\ : Span4Mux_h
    port map (
            O => \N__14046\,
            I => \N__14040\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__14043\,
            I => \N__14037\
        );

    \I__2715\ : Odrv4
    port map (
            O => \N__14040\,
            I => \c0.rx.N_335\
        );

    \I__2714\ : Odrv12
    port map (
            O => \N__14037\,
            I => \c0.rx.N_335\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14029\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__14029\,
            I => \c0.N_121\
        );

    \I__2711\ : InMux
    port map (
            O => \N__14026\,
            I => \N__14023\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__14023\,
            I => \c0.m163_4\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14020\,
            I => \N__14017\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__14017\,
            I => \N__14014\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__14014\,
            I => \c0.un1_data_in_7__1_0_a2_24_a2_7\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14008\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__14008\,
            I => \N__14005\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__14005\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_6\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__14002\,
            I => \c0.m163_8_cascade_\
        );

    \I__2702\ : InMux
    port map (
            O => \N__13999\,
            I => \N__13996\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__13996\,
            I => \c0.un1_data_in_7__1_3\
        );

    \I__2700\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13990\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__13990\,
            I => \c0.m163_10\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__13987\,
            I => \c0.m163_1_cascade_\
        );

    \I__2697\ : InMux
    port map (
            O => \N__13984\,
            I => \N__13981\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__13981\,
            I => \c0.un1_data_in_7__0\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__13978\,
            I => \c0.N_164_0_cascade_\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__13975\,
            I => \c0.N_173_0_cascade_\
        );

    \I__2693\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13969\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__13969\,
            I => \N__13966\
        );

    \I__2691\ : Span4Mux_h
    port map (
            O => \N__13966\,
            I => \N__13961\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__13965\,
            I => \N__13958\
        );

    \I__2689\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13955\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__13961\,
            I => \N__13952\
        );

    \I__2687\ : InMux
    port map (
            O => \N__13958\,
            I => \N__13949\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__13955\,
            I => \c0.data_in_3_Z0Z_7\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__13952\,
            I => \c0.data_in_3_Z0Z_7\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__13949\,
            I => \c0.data_in_3_Z0Z_7\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13942\,
            I => \N__13939\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__13939\,
            I => \c0.d_4_RNIB3JJZ0Z_2\
        );

    \I__2681\ : InMux
    port map (
            O => \N__13936\,
            I => \N__13931\
        );

    \I__2680\ : InMux
    port map (
            O => \N__13935\,
            I => \N__13928\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__13934\,
            I => \N__13924\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__13931\,
            I => \N__13921\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__13928\,
            I => \N__13918\
        );

    \I__2676\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13915\
        );

    \I__2675\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13912\
        );

    \I__2674\ : Odrv4
    port map (
            O => \N__13921\,
            I => \c0.d_4_44\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__13918\,
            I => \c0.d_4_44\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__13915\,
            I => \c0.d_4_44\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__13912\,
            I => \c0.d_4_44\
        );

    \I__2670\ : InMux
    port map (
            O => \N__13903\,
            I => \N__13897\
        );

    \I__2669\ : InMux
    port map (
            O => \N__13902\,
            I => \N__13890\
        );

    \I__2668\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13890\
        );

    \I__2667\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13890\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__13897\,
            I => \c0.d_4_36\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__13890\,
            I => \c0.d_4_36\
        );

    \I__2664\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13878\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13884\,
            I => \N__13878\
        );

    \I__2662\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13875\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__13878\,
            I => \c0.N_104\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__13875\,
            I => \c0.N_104\
        );

    \I__2659\ : InMux
    port map (
            O => \N__13870\,
            I => \N__13867\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__13867\,
            I => \N__13864\
        );

    \I__2657\ : Span4Mux_h
    port map (
            O => \N__13864\,
            I => \N__13861\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__13861\,
            I => \c0.un1_data_in_6__3_0_a2_5_a2_2\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__13858\,
            I => \c0.un1_data_in_6__5_cascade_\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13855\,
            I => \N__13852\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__13852\,
            I => \c0.un1_data_in_6__6\
        );

    \I__2652\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13846\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__13846\,
            I => \c0.un1_data_in_6__1_0_a2_4_a2_2\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__13843\,
            I => \c0.m163_2_cascade_\
        );

    \I__2649\ : InMux
    port map (
            O => \N__13840\,
            I => \N__13837\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__13837\,
            I => \N__13834\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__13834\,
            I => \N__13830\
        );

    \I__2646\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13827\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__13830\,
            I => \c0.N_126\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__13827\,
            I => \c0.N_126\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__13822\,
            I => \c0.m163_7_cascade_\
        );

    \I__2642\ : InMux
    port map (
            O => \N__13819\,
            I => \N__13816\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__13816\,
            I => \N__13813\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__13813\,
            I => \c0.m163_0\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__13810\,
            I => \N__13807\
        );

    \I__2638\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13804\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__13804\,
            I => \c0.un1_data_in_6__5_0_a2_5_a2_2\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13798\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__13798\,
            I => \N__13794\
        );

    \I__2634\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13790\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__13794\,
            I => \N__13787\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13784\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__13790\,
            I => \c0.N_120\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__13787\,
            I => \c0.N_120\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__13784\,
            I => \c0.N_120\
        );

    \I__2628\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13774\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__13774\,
            I => \N__13770\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13767\
        );

    \I__2625\ : Span4Mux_h
    port map (
            O => \N__13770\,
            I => \N__13763\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__13767\,
            I => \N__13760\
        );

    \I__2623\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13757\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__13763\,
            I => \c0.data_in_1_Z0Z_4\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__13760\,
            I => \c0.data_in_1_Z0Z_4\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__13757\,
            I => \c0.data_in_1_Z0Z_4\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__13750\,
            I => \N__13745\
        );

    \I__2618\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13740\
        );

    \I__2617\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13740\
        );

    \I__2616\ : InMux
    port map (
            O => \N__13745\,
            I => \N__13737\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__13740\,
            I => \c0.d_4_6\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__13737\,
            I => \c0.d_4_6\
        );

    \I__2613\ : InMux
    port map (
            O => \N__13732\,
            I => \N__13729\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__13729\,
            I => \N__13726\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__13726\,
            I => \c0.N_109\
        );

    \I__2610\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13720\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__13720\,
            I => \N__13717\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__13717\,
            I => \N__13713\
        );

    \I__2607\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13710\
        );

    \I__2606\ : Span4Mux_h
    port map (
            O => \N__13713\,
            I => \N__13704\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__13710\,
            I => \N__13704\
        );

    \I__2604\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13701\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__13704\,
            I => \c0.data_in_1_Z0Z_6\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__13701\,
            I => \c0.data_in_1_Z0Z_6\
        );

    \I__2601\ : InMux
    port map (
            O => \N__13696\,
            I => \N__13693\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__13693\,
            I => \N__13690\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__13690\,
            I => \N__13685\
        );

    \I__2598\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13680\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13688\,
            I => \N__13680\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__13685\,
            I => \c0.d_4_7\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__13680\,
            I => \c0.d_4_7\
        );

    \I__2594\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13672\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__13672\,
            I => \N__13669\
        );

    \I__2592\ : Span4Mux_v
    port map (
            O => \N__13669\,
            I => \N__13666\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__13666\,
            I => \c0.tx2_data_RNO_3Z0Z_7\
        );

    \I__2590\ : InMux
    port map (
            O => \N__13663\,
            I => \N__13660\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__13660\,
            I => \N__13656\
        );

    \I__2588\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13653\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__13656\,
            I => \N__13650\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__13653\,
            I => \N__13647\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__13650\,
            I => \c0.data_in_4_Z0Z_4\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__13647\,
            I => \c0.data_in_4_Z0Z_4\
        );

    \I__2583\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13637\
        );

    \I__2582\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13634\
        );

    \I__2581\ : InMux
    port map (
            O => \N__13640\,
            I => \N__13631\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__13637\,
            I => \N__13628\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__13634\,
            I => \c0.data_in_6_Z0Z_1\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__13631\,
            I => \c0.data_in_6_Z0Z_1\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__13628\,
            I => \c0.data_in_6_Z0Z_1\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__13621\,
            I => \c0.N_34_cascade_\
        );

    \I__2575\ : InMux
    port map (
            O => \N__13618\,
            I => \N__13614\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__13617\,
            I => \N__13610\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__13614\,
            I => \N__13607\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13604\
        );

    \I__2571\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13601\
        );

    \I__2570\ : Odrv12
    port map (
            O => \N__13607\,
            I => \c0.data_in_2_Z0Z_6\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__13604\,
            I => \c0.data_in_2_Z0Z_6\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__13601\,
            I => \c0.data_in_2_Z0Z_6\
        );

    \I__2567\ : InMux
    port map (
            O => \N__13594\,
            I => \N__13591\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__13591\,
            I => \c0.byte_transmit_counterZ0Z_5\
        );

    \I__2565\ : InMux
    port map (
            O => \N__13588\,
            I => \N__13585\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__13585\,
            I => \N__13580\
        );

    \I__2563\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13577\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__13583\,
            I => \N__13574\
        );

    \I__2561\ : Span4Mux_v
    port map (
            O => \N__13580\,
            I => \N__13571\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__13577\,
            I => \N__13568\
        );

    \I__2559\ : InMux
    port map (
            O => \N__13574\,
            I => \N__13565\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__13571\,
            I => \c0.data_in_6_Z0Z_7\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__13568\,
            I => \c0.data_in_6_Z0Z_7\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__13565\,
            I => \c0.data_in_6_Z0Z_7\
        );

    \I__2555\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13555\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__13555\,
            I => \c0.data_in_frame_6_Z0Z_7\
        );

    \I__2553\ : InMux
    port map (
            O => \N__13552\,
            I => \N__13549\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__13549\,
            I => \N__13545\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13542\
        );

    \I__2550\ : Span4Mux_h
    port map (
            O => \N__13545\,
            I => \N__13536\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__13542\,
            I => \N__13536\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__13541\,
            I => \N__13533\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__13536\,
            I => \N__13530\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13527\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__13530\,
            I => \c0.data_in_7_Z0Z_7\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__13527\,
            I => \c0.data_in_7_Z0Z_7\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__13522\,
            I => \N__13519\
        );

    \I__2542\ : InMux
    port map (
            O => \N__13519\,
            I => \N__13516\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__13516\,
            I => \c0.data_in_frame_7_Z0Z_7\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13510\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__13510\,
            I => \N__13507\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__13507\,
            I => \N__13503\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__13506\,
            I => \N__13500\
        );

    \I__2536\ : Span4Mux_v
    port map (
            O => \N__13503\,
            I => \N__13497\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13500\,
            I => \N__13494\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__13497\,
            I => \c0.data_in_0_Z0Z_6\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__13494\,
            I => \c0.data_in_0_Z0Z_6\
        );

    \I__2532\ : InMux
    port map (
            O => \N__13489\,
            I => \N__13486\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__13486\,
            I => \N__13481\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13485\,
            I => \N__13478\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13484\,
            I => \N__13475\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__13481\,
            I => \N__13472\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__13478\,
            I => \N__13467\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13475\,
            I => \N__13467\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__13472\,
            I => \N__13464\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__13467\,
            I => \c0.d_2_9\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__13464\,
            I => \c0.d_2_9\
        );

    \I__2522\ : InMux
    port map (
            O => \N__13459\,
            I => \N__13456\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__13456\,
            I => \c0.tx_data_RNO_3Z0Z_1\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__13453\,
            I => \N__13449\
        );

    \I__2519\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13445\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13442\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__13448\,
            I => \N__13438\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__13445\,
            I => \N__13433\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__13442\,
            I => \N__13433\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13441\,
            I => \N__13428\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13438\,
            I => \N__13428\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__13433\,
            I => \c0.d_2_2\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__13428\,
            I => \c0.d_2_2\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__13423\,
            I => \c0.tx_data_RNO_3Z0Z_2_cascade_\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13420\,
            I => \N__13417\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__13417\,
            I => \c0.tx_data_RNO_4Z0Z_2\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13411\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13411\,
            I => \c0.tx_data_1_0_i_ns_1_2\
        );

    \I__2505\ : InMux
    port map (
            O => \N__13408\,
            I => \N__13405\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__13405\,
            I => \N__13401\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13404\,
            I => \N__13396\
        );

    \I__2502\ : Span4Mux_v
    port map (
            O => \N__13401\,
            I => \N__13392\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13400\,
            I => \N__13389\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13399\,
            I => \N__13386\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__13396\,
            I => \N__13383\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13395\,
            I => \N__13380\
        );

    \I__2497\ : Span4Mux_h
    port map (
            O => \N__13392\,
            I => \N__13375\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__13389\,
            I => \N__13375\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__13386\,
            I => \c0.d_2_39\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__13383\,
            I => \c0.d_2_39\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__13380\,
            I => \c0.d_2_39\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__13375\,
            I => \c0.d_2_39\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__13366\,
            I => \N__13362\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13365\,
            I => \N__13358\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13362\,
            I => \N__13355\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__13361\,
            I => \N__13352\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__13358\,
            I => \N__13347\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__13355\,
            I => \N__13347\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13352\,
            I => \N__13344\
        );

    \I__2484\ : Odrv12
    port map (
            O => \N__13347\,
            I => \c0.d_2_47\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__13344\,
            I => \c0.d_2_47\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13336\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13336\,
            I => \N__13333\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__13333\,
            I => \c0.tx_data_RNO_0Z0Z_7\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13330\,
            I => \N__13324\
        );

    \I__2478\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13321\
        );

    \I__2477\ : InMux
    port map (
            O => \N__13328\,
            I => \N__13316\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13327\,
            I => \N__13316\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__13324\,
            I => \N__13313\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__13321\,
            I => \N__13308\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__13316\,
            I => \N__13308\
        );

    \I__2472\ : Odrv4
    port map (
            O => \N__13313\,
            I => \c0.d_2_36\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__13308\,
            I => \c0.d_2_36\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__13303\,
            I => \N__13300\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13297\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13297\,
            I => \N__13294\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__13294\,
            I => \N__13290\
        );

    \I__2466\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13287\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__13290\,
            I => \c0.d_2_44\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__13287\,
            I => \c0.d_2_44\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13282\,
            I => \N__13279\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__13279\,
            I => \N__13276\
        );

    \I__2461\ : Span4Mux_h
    port map (
            O => \N__13276\,
            I => \N__13273\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__13273\,
            I => \c0.tx_data_RNO_0Z0Z_4\
        );

    \I__2459\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13267\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__13267\,
            I => \N__13264\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__13264\,
            I => \c0.data_out_6_Z0Z_1\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__13261\,
            I => \N__13258\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13255\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__13255\,
            I => \N__13252\
        );

    \I__2453\ : Span4Mux_v
    port map (
            O => \N__13252\,
            I => \N__13249\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__13249\,
            I => \c0.data_out_7_Z0Z_1\
        );

    \I__2451\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13243\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__13243\,
            I => \N__13240\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__13240\,
            I => \c0.tx_data_RNO_1Z0Z_1\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__13237\,
            I => \c0.m2_e_1_cascade_\
        );

    \I__2447\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__13231\,
            I => \c0.data_out_7_Z0Z_3\
        );

    \I__2445\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13225\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__13225\,
            I => \N__13222\
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__13222\,
            I => \c0.data_out_6_Z0Z_3\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__13219\,
            I => \c0.N_132_mux_cascade_\
        );

    \I__2441\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13213\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13213\,
            I => \N__13210\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__13210\,
            I => \N__13207\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__13207\,
            I => \c0.tx_data_RNO_1Z0Z_3\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13204\,
            I => \N__13201\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__13201\,
            I => \c0.tx_data_RNO_4Z0Z_5\
        );

    \I__2435\ : InMux
    port map (
            O => \N__13198\,
            I => \N__13195\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__13195\,
            I => \N__13192\
        );

    \I__2433\ : Span4Mux_h
    port map (
            O => \N__13192\,
            I => \N__13189\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__13189\,
            I => \c0.tx_data_RNO_1Z0Z_0\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13186\,
            I => \N__13183\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__13183\,
            I => \c0.tx_data_RNO_0Z0Z_0\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13180\,
            I => \N__13177\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__13177\,
            I => \c0.tx_data_1_0_i_ns_1_0\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13171\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__13171\,
            I => \N__13168\
        );

    \I__2425\ : Span4Mux_h
    port map (
            O => \N__13168\,
            I => \N__13165\
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__13165\,
            I => \c0.tx.r_Tx_DataZ0Z_0\
        );

    \I__2423\ : InMux
    port map (
            O => \N__13162\,
            I => \N__13159\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13159\,
            I => \c0.tx_data_RNO_0Z0Z_2\
        );

    \I__2421\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13153\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__13153\,
            I => \N__13150\
        );

    \I__2419\ : Span4Mux_h
    port map (
            O => \N__13150\,
            I => \N__13147\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__13147\,
            I => \c0.tx.r_Tx_DataZ0Z_2\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__13144\,
            I => \N__13141\
        );

    \I__2416\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13137\
        );

    \I__2415\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13132\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__13137\,
            I => \N__13129\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13136\,
            I => \N__13124\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13135\,
            I => \N__13124\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__13132\,
            I => \N__13121\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__13129\,
            I => \N__13118\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__13124\,
            I => \N__13115\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__13121\,
            I => \c0.d_2_25\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__13118\,
            I => \c0.d_2_25\
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__13115\,
            I => \c0.d_2_25\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__13108\,
            I => \c0.tx_data_RNO_4Z0Z_1_cascade_\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13105\,
            I => \N__13102\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13102\,
            I => \c0.tx_data_RNO_0Z0Z_1\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__13099\,
            I => \c0.tx_data_1_0_i_ns_1_1_cascade_\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13096\,
            I => \N__13093\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__13093\,
            I => \N__13090\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__13090\,
            I => \N__13087\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__13087\,
            I => \c0.tx.r_Tx_DataZ0Z_1\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13084\,
            I => \N__13081\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__13081\,
            I => \N__13078\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__13078\,
            I => \N__13075\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__13075\,
            I => \c0.data_out_7_Z0Z_2\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13072\,
            I => \N__13069\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__13069\,
            I => \N__13066\
        );

    \I__2391\ : Span4Mux_v
    port map (
            O => \N__13066\,
            I => \N__13063\
        );

    \I__2390\ : Odrv4
    port map (
            O => \N__13063\,
            I => \c0.data_out_6_Z0Z_2\
        );

    \I__2389\ : InMux
    port map (
            O => \N__13060\,
            I => \N__13057\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__13057\,
            I => \c0.tx_data_RNO_1Z0Z_2\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13054\,
            I => \N__13051\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__13051\,
            I => \N__13046\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13050\,
            I => \N__13043\
        );

    \I__2384\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13040\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__13046\,
            I => \N__13032\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13043\,
            I => \N__13032\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__13040\,
            I => \N__13032\
        );

    \I__2380\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13029\
        );

    \I__2379\ : Span4Mux_h
    port map (
            O => \N__13032\,
            I => \N__13026\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__13029\,
            I => \c0.d_2_1\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__13026\,
            I => \c0.d_2_1\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__13021\,
            I => \N__13017\
        );

    \I__2375\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13014\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13017\,
            I => \N__13010\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13014\,
            I => \N__13006\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13013\,
            I => \N__13003\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__13010\,
            I => \N__13000\
        );

    \I__2370\ : InMux
    port map (
            O => \N__13009\,
            I => \N__12997\
        );

    \I__2369\ : Span4Mux_h
    port map (
            O => \N__13006\,
            I => \N__12988\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__13003\,
            I => \N__12988\
        );

    \I__2367\ : Span4Mux_h
    port map (
            O => \N__13000\,
            I => \N__12988\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__12997\,
            I => \N__12988\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__12988\,
            I => \c0.d_2_37\
        );

    \I__2364\ : InMux
    port map (
            O => \N__12985\,
            I => \N__12981\
        );

    \I__2363\ : InMux
    port map (
            O => \N__12984\,
            I => \N__12978\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__12981\,
            I => \N__12975\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__12978\,
            I => \N__12972\
        );

    \I__2360\ : Span4Mux_v
    port map (
            O => \N__12975\,
            I => \N__12969\
        );

    \I__2359\ : Span4Mux_v
    port map (
            O => \N__12972\,
            I => \N__12966\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__12969\,
            I => \c0.d_2_45\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__12966\,
            I => \c0.d_2_45\
        );

    \I__2356\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12958\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__12958\,
            I => \c0.tx_data_RNO_0Z0Z_5\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__12955\,
            I => \c0.tx_data_RNO_3Z0Z_6_cascade_\
        );

    \I__2353\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12949\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__12949\,
            I => \c0.tx_data_RNO_4Z0Z_6\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__12946\,
            I => \N__12943\
        );

    \I__2350\ : InMux
    port map (
            O => \N__12943\,
            I => \N__12938\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__12942\,
            I => \N__12935\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__12941\,
            I => \N__12930\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__12938\,
            I => \N__12927\
        );

    \I__2346\ : InMux
    port map (
            O => \N__12935\,
            I => \N__12924\
        );

    \I__2345\ : InMux
    port map (
            O => \N__12934\,
            I => \N__12921\
        );

    \I__2344\ : InMux
    port map (
            O => \N__12933\,
            I => \N__12916\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12930\,
            I => \N__12916\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__12927\,
            I => \N__12913\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__12924\,
            I => \N__12908\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__12921\,
            I => \N__12908\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__12916\,
            I => \N__12905\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__12913\,
            I => \N__12902\
        );

    \I__2337\ : Span4Mux_v
    port map (
            O => \N__12908\,
            I => \N__12899\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__12905\,
            I => \N__12896\
        );

    \I__2335\ : Span4Mux_h
    port map (
            O => \N__12902\,
            I => \N__12893\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__12899\,
            I => \c0.d_2_42\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__12896\,
            I => \c0.d_2_42\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__12893\,
            I => \c0.d_2_42\
        );

    \I__2331\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12883\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__12883\,
            I => \c0.nextCRC16_3_3_1\
        );

    \I__2329\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12875\
        );

    \I__2328\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12870\
        );

    \I__2327\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12870\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__12875\,
            I => \N__12865\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__12870\,
            I => \N__12865\
        );

    \I__2324\ : Span4Mux_h
    port map (
            O => \N__12865\,
            I => \N__12861\
        );

    \I__2323\ : InMux
    port map (
            O => \N__12864\,
            I => \N__12858\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__12861\,
            I => \c0.d_2_4\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__12858\,
            I => \c0.d_2_4\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__12853\,
            I => \c0.nextCRC16_3_3_1_cascade_\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__12850\,
            I => \N__12847\
        );

    \I__2318\ : InMux
    port map (
            O => \N__12847\,
            I => \N__12844\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__12844\,
            I => \N__12841\
        );

    \I__2316\ : Span4Mux_h
    port map (
            O => \N__12841\,
            I => \N__12838\
        );

    \I__2315\ : Span4Mux_h
    port map (
            O => \N__12838\,
            I => \N__12835\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__12835\,
            I => \c0.nextCRC16_3_0_a2_1_1\
        );

    \I__2313\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12829\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__12829\,
            I => \N__12824\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12821\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12818\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__12824\,
            I => \c0.d_2_28\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__12821\,
            I => \c0.d_2_28\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__12818\,
            I => \c0.d_2_28\
        );

    \I__2306\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12807\
        );

    \I__2305\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12804\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__12807\,
            I => \N__12800\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__12804\,
            I => \N__12797\
        );

    \I__2302\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12794\
        );

    \I__2301\ : Span4Mux_h
    port map (
            O => \N__12800\,
            I => \N__12791\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__12797\,
            I => \N__12786\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__12794\,
            I => \N__12786\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__12791\,
            I => \N__12783\
        );

    \I__2297\ : Span4Mux_h
    port map (
            O => \N__12786\,
            I => \N__12780\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__12783\,
            I => \c0.d_2_5\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__12780\,
            I => \c0.d_2_5\
        );

    \I__2294\ : InMux
    port map (
            O => \N__12775\,
            I => \N__12771\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__12774\,
            I => \N__12768\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__12771\,
            I => \N__12764\
        );

    \I__2291\ : InMux
    port map (
            O => \N__12768\,
            I => \N__12759\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12767\,
            I => \N__12759\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__12764\,
            I => \c0.d_2_13\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__12759\,
            I => \c0.d_2_13\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__12754\,
            I => \c0.tx_data_RNO_3Z0Z_5_cascade_\
        );

    \I__2286\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12748\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__12748\,
            I => \c0.tx_data_1_0_i_ns_1_5\
        );

    \I__2284\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12742\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__12742\,
            I => \N__12739\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__12739\,
            I => \N__12735\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12732\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__12735\,
            I => \c0.N_108\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__12732\,
            I => \c0.N_108\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__12727\,
            I => \c0.un1_data_in_7__6_0_a2_5_a2_2_cascade_\
        );

    \I__2277\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12721\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__12721\,
            I => \c0.un1_data_in_7__4_0_a2_0_a2_4\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12718\,
            I => \N__12715\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__12715\,
            I => \N__12712\
        );

    \I__2273\ : Span4Mux_h
    port map (
            O => \N__12712\,
            I => \N__12708\
        );

    \I__2272\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12705\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__12708\,
            I => \c0.data_in_0_Z0Z_3\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__12705\,
            I => \c0.data_in_0_Z0Z_3\
        );

    \I__2269\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12697\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__12697\,
            I => \N__12694\
        );

    \I__2267\ : Span4Mux_h
    port map (
            O => \N__12694\,
            I => \N__12690\
        );

    \I__2266\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12687\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__12690\,
            I => \c0.data_in_0_Z0Z_5\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__12687\,
            I => \c0.data_in_0_Z0Z_5\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12682\,
            I => \N__12679\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__12679\,
            I => \N__12676\
        );

    \I__2261\ : Span4Mux_v
    port map (
            O => \N__12676\,
            I => \N__12671\
        );

    \I__2260\ : InMux
    port map (
            O => \N__12675\,
            I => \N__12666\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12674\,
            I => \N__12666\
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__12671\,
            I => \c0.data_in_2_Z0Z_2\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__12666\,
            I => \c0.data_in_2_Z0Z_2\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__12661\,
            I => \N__12658\
        );

    \I__2255\ : InMux
    port map (
            O => \N__12658\,
            I => \N__12653\
        );

    \I__2254\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12648\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12648\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__12653\,
            I => \c0.d_4_18\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__12648\,
            I => \c0.d_4_18\
        );

    \I__2250\ : InMux
    port map (
            O => \N__12643\,
            I => \N__12638\
        );

    \I__2249\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12632\
        );

    \I__2248\ : InMux
    port map (
            O => \N__12641\,
            I => \N__12632\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12638\,
            I => \N__12629\
        );

    \I__2246\ : InMux
    port map (
            O => \N__12637\,
            I => \N__12626\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__12632\,
            I => \N__12623\
        );

    \I__2244\ : Span4Mux_h
    port map (
            O => \N__12629\,
            I => \N__12618\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__12626\,
            I => \N__12618\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__12623\,
            I => \c0.d_2_38\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__12618\,
            I => \c0.d_2_38\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__12613\,
            I => \N__12610\
        );

    \I__2239\ : InMux
    port map (
            O => \N__12610\,
            I => \N__12607\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__12607\,
            I => \N__12603\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12599\
        );

    \I__2236\ : Span4Mux_h
    port map (
            O => \N__12603\,
            I => \N__12596\
        );

    \I__2235\ : InMux
    port map (
            O => \N__12602\,
            I => \N__12593\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__12599\,
            I => \c0.d_2_46\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__12596\,
            I => \c0.d_2_46\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__12593\,
            I => \c0.d_2_46\
        );

    \I__2231\ : InMux
    port map (
            O => \N__12586\,
            I => \N__12583\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__12583\,
            I => \N__12580\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__12580\,
            I => \N__12577\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__12577\,
            I => \c0.data_out_6_Z0Z_7\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__12574\,
            I => \N__12571\
        );

    \I__2226\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12568\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__12568\,
            I => \N__12565\
        );

    \I__2224\ : Span12Mux_h
    port map (
            O => \N__12565\,
            I => \N__12562\
        );

    \I__2223\ : Odrv12
    port map (
            O => \N__12562\,
            I => \c0.data_out_7_Z0Z_7\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12556\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__12556\,
            I => \c0.tx_data_RNO_1Z0Z_7\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__12553\,
            I => \c0.un1_data_in_7__1_0_a2_24_a2_3_cascade_\
        );

    \I__2219\ : InMux
    port map (
            O => \N__12550\,
            I => \N__12547\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__12547\,
            I => \c0.un1_data_in_7__1_0_a2_24_a2_4\
        );

    \I__2217\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12541\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__12541\,
            I => \N__12538\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__12538\,
            I => \N__12534\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12531\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__12534\,
            I => \c0.data_in_5_Z0Z_4\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12531\,
            I => \c0.data_in_5_Z0Z_4\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12526\,
            I => \N__12523\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__12523\,
            I => \N__12520\
        );

    \I__2209\ : Span4Mux_h
    port map (
            O => \N__12520\,
            I => \N__12516\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12519\,
            I => \N__12513\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__12516\,
            I => \c0.data_in_5_Z0Z_2\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__12513\,
            I => \c0.data_in_5_Z0Z_2\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12508\,
            I => \N__12505\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12505\,
            I => \N__12501\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__12504\,
            I => \N__12497\
        );

    \I__2202\ : Span4Mux_v
    port map (
            O => \N__12501\,
            I => \N__12494\
        );

    \I__2201\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12491\
        );

    \I__2200\ : InMux
    port map (
            O => \N__12497\,
            I => \N__12488\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__12494\,
            I => \c0.data_in_2_Z0Z_0\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__12491\,
            I => \c0.data_in_2_Z0Z_0\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__12488\,
            I => \c0.data_in_2_Z0Z_0\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__12481\,
            I => \N__12476\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12473\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12469\
        );

    \I__2193\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12466\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12473\,
            I => \N__12463\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12472\,
            I => \N__12460\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12469\,
            I => \N__12455\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12466\,
            I => \N__12455\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__12463\,
            I => \c0.d_4_33\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__12460\,
            I => \c0.d_4_33\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__12455\,
            I => \c0.d_4_33\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__12448\,
            I => \c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12442\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__12442\,
            I => \N__12439\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__12439\,
            I => \c0.N_124\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__12436\,
            I => \c0.N_124_cascade_\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__12433\,
            I => \c0.un1_data_in_7__0_0_a2_1_a2_5_cascade_\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__12430\,
            I => \c0.N_121_cascade_\
        );

    \I__2178\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12423\
        );

    \I__2177\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12420\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__12423\,
            I => \N__12417\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__12420\,
            I => \c0.N_125\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__12417\,
            I => \c0.N_125\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__12412\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_4_3_cascade_\
        );

    \I__2172\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12406\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12406\,
            I => \c0.N_136\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__12403\,
            I => \c0.N_136_cascade_\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__12400\,
            I => \N__12397\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12394\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__12394\,
            I => \N__12391\
        );

    \I__2166\ : Odrv12
    port map (
            O => \N__12391\,
            I => \c0.un1_data_in_7__0_0_a2_1_a2_2\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__12388\,
            I => \N__12383\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12380\
        );

    \I__2163\ : InMux
    port map (
            O => \N__12386\,
            I => \N__12377\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12383\,
            I => \N__12374\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__12380\,
            I => \N__12371\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__12377\,
            I => \N__12366\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12374\,
            I => \N__12366\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__12371\,
            I => \c0.data_in_3_Z0Z_3\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__12366\,
            I => \c0.data_in_3_Z0Z_3\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__12361\,
            I => \c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_\
        );

    \I__2155\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12354\
        );

    \I__2154\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12351\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__12354\,
            I => \N__12348\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__12351\,
            I => \N__12344\
        );

    \I__2151\ : Span4Mux_h
    port map (
            O => \N__12348\,
            I => \N__12341\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12338\
        );

    \I__2149\ : Odrv12
    port map (
            O => \N__12344\,
            I => \c0.data_in_3_Z0Z_4\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__12341\,
            I => \c0.data_in_3_Z0Z_4\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__12338\,
            I => \c0.data_in_3_Z0Z_4\
        );

    \I__2146\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12328\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__12328\,
            I => \N__12325\
        );

    \I__2144\ : Span4Mux_h
    port map (
            O => \N__12325\,
            I => \N__12320\
        );

    \I__2143\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12315\
        );

    \I__2142\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12315\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__12320\,
            I => \c0.data_in_1_Z0Z_5\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__12315\,
            I => \c0.data_in_1_Z0Z_5\
        );

    \I__2139\ : InMux
    port map (
            O => \N__12310\,
            I => \N__12307\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__12307\,
            I => \N__12302\
        );

    \I__2137\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12297\
        );

    \I__2136\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12297\
        );

    \I__2135\ : Odrv12
    port map (
            O => \N__12302\,
            I => \c0.data_in_3_Z0Z_2\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__12297\,
            I => \c0.data_in_3_Z0Z_2\
        );

    \I__2133\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12289\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__12289\,
            I => \N__12285\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12288\,
            I => \N__12282\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__12285\,
            I => \c0.data_in_5_Z0Z_1\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12282\,
            I => \c0.data_in_5_Z0Z_1\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12274\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__12274\,
            I => \N__12271\
        );

    \I__2126\ : Span4Mux_h
    port map (
            O => \N__12271\,
            I => \N__12267\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12270\,
            I => \N__12264\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__12267\,
            I => \c0.data_in_5_Z0Z_0\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__12264\,
            I => \c0.data_in_5_Z0Z_0\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12259\,
            I => \N__12255\
        );

    \I__2121\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12252\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__12255\,
            I => \N__12246\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12252\,
            I => \N__12246\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12251\,
            I => \N__12243\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__12246\,
            I => \c0.N_132\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__12243\,
            I => \c0.N_132\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12235\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12235\,
            I => \N__12232\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__12232\,
            I => \N__12229\
        );

    \I__2112\ : Span4Mux_h
    port map (
            O => \N__12229\,
            I => \N__12225\
        );

    \I__2111\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12222\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__12225\,
            I => \c0.rx_data_4\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12222\,
            I => \c0.rx_data_4\
        );

    \I__2108\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12214\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__12214\,
            I => \N__12211\
        );

    \I__2106\ : Span12Mux_v
    port map (
            O => \N__12211\,
            I => \N__12207\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12210\,
            I => \N__12204\
        );

    \I__2104\ : Odrv12
    port map (
            O => \N__12207\,
            I => \c0.rx_data_2\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__12204\,
            I => \c0.rx_data_2\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12195\
        );

    \I__2101\ : InMux
    port map (
            O => \N__12198\,
            I => \N__12190\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__12195\,
            I => \N__12187\
        );

    \I__2099\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12184\
        );

    \I__2098\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12181\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__12190\,
            I => \N__12178\
        );

    \I__2096\ : Odrv12
    port map (
            O => \N__12187\,
            I => \c0.d_4_34\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__12184\,
            I => \c0.d_4_34\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__12181\,
            I => \c0.d_4_34\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__12178\,
            I => \c0.d_4_34\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__12169\,
            I => \c0.un1_data_in_7__7_0_a2_0_a2_2_cascade_\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12163\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__12163\,
            I => \N__12160\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__12160\,
            I => \c0.un1_data_in_6__0_0_a2_5_a2_2\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__12157\,
            I => \c0.un1_data_in_7__7_i_cascade_\
        );

    \I__2087\ : InMux
    port map (
            O => \N__12154\,
            I => \N__12151\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__12151\,
            I => \N__12147\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12144\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__12147\,
            I => \c0.data_in_5_Z0Z_7\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__12144\,
            I => \c0.data_in_5_Z0Z_7\
        );

    \I__2082\ : InMux
    port map (
            O => \N__12139\,
            I => \N__12135\
        );

    \I__2081\ : InMux
    port map (
            O => \N__12138\,
            I => \N__12132\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__12135\,
            I => \N__12129\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__12132\,
            I => \N__12126\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__12129\,
            I => \c0.data_in_4_Z0Z_3\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__12126\,
            I => \c0.data_in_4_Z0Z_3\
        );

    \I__2076\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12115\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12115\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__12115\,
            I => \N__12110\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12107\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12104\
        );

    \I__2071\ : Span4Mux_h
    port map (
            O => \N__12110\,
            I => \N__12101\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__12107\,
            I => \N__12098\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__12104\,
            I => \c0.d_2_32\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__12101\,
            I => \c0.d_2_32\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__12098\,
            I => \c0.d_2_32\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__12091\,
            I => \N__12087\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__12090\,
            I => \N__12083\
        );

    \I__2064\ : InMux
    port map (
            O => \N__12087\,
            I => \N__12079\
        );

    \I__2063\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12074\
        );

    \I__2062\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12074\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__12082\,
            I => \N__12071\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__12079\,
            I => \N__12068\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__12074\,
            I => \N__12065\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12062\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__12068\,
            I => \N__12059\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__12065\,
            I => \N__12056\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__12062\,
            I => \c0.d_2_24\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__12059\,
            I => \c0.d_2_24\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__12056\,
            I => \c0.d_2_24\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12046\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12046\,
            I => \c0.nextCRC16_3_3_12\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__12043\,
            I => \c0.nextCRC16_3_4_12_cascade_\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12037\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__12037\,
            I => \N__12032\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12036\,
            I => \N__12029\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12035\,
            I => \N__12026\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__12032\,
            I => \N__12019\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__12029\,
            I => \N__12019\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__12026\,
            I => \N__12019\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__12019\,
            I => \N__12016\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__12016\,
            I => \c0.d_2_41\
        );

    \I__2040\ : InMux
    port map (
            O => \N__12013\,
            I => \N__12010\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__12010\,
            I => \N__12007\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__12007\,
            I => \N__12004\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__12004\,
            I => \c0.N_94\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__12001\,
            I => \c0.N_94_cascade_\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__11998\,
            I => \N__11993\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__11997\,
            I => \N__11989\
        );

    \I__2033\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11986\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11983\
        );

    \I__2031\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11980\
        );

    \I__2030\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11977\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__11986\,
            I => \N__11974\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__11983\,
            I => \N__11969\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__11980\,
            I => \N__11969\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__11977\,
            I => \N__11964\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__11974\,
            I => \N__11964\
        );

    \I__2024\ : Odrv12
    port map (
            O => \N__11969\,
            I => \c0.d_2_23\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__11964\,
            I => \c0.d_2_23\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__11959\,
            I => \N__11956\
        );

    \I__2021\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11951\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__11955\,
            I => \N__11948\
        );

    \I__2019\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11944\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__11951\,
            I => \N__11941\
        );

    \I__2017\ : InMux
    port map (
            O => \N__11948\,
            I => \N__11935\
        );

    \I__2016\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11935\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__11944\,
            I => \N__11930\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__11941\,
            I => \N__11930\
        );

    \I__2013\ : InMux
    port map (
            O => \N__11940\,
            I => \N__11927\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__11935\,
            I => \N__11924\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__11930\,
            I => \c0.d_2_40\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__11927\,
            I => \c0.d_2_40\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__11924\,
            I => \c0.d_2_40\
        );

    \I__2008\ : InMux
    port map (
            O => \N__11917\,
            I => \N__11914\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__11914\,
            I => \c0.nextCRC16_3_0_a2_1_11\
        );

    \I__2006\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11908\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__11908\,
            I => \c0.data_out_6_Z0Z_4\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__11905\,
            I => \N__11902\
        );

    \I__2003\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11899\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__11899\,
            I => \N__11896\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__11896\,
            I => \N__11893\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__11893\,
            I => \c0.data_out_7_Z0Z_4\
        );

    \I__1999\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11887\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__11887\,
            I => \N__11884\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__11884\,
            I => \N__11881\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__11881\,
            I => \c0.tx_data_RNO_1Z0Z_4\
        );

    \I__1995\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11874\
        );

    \I__1994\ : InMux
    port map (
            O => \N__11877\,
            I => \N__11871\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__11874\,
            I => \c0.data_in_5_Z0Z_5\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__11871\,
            I => \c0.data_in_5_Z0Z_5\
        );

    \I__1991\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11863\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__11863\,
            I => \N__11859\
        );

    \I__1989\ : InMux
    port map (
            O => \N__11862\,
            I => \N__11856\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__11859\,
            I => \N__11851\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__11856\,
            I => \N__11851\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__11851\,
            I => \N__11848\
        );

    \I__1985\ : Span4Mux_h
    port map (
            O => \N__11848\,
            I => \N__11845\
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__11845\,
            I => \c0.d_2_8\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__11842\,
            I => \N__11839\
        );

    \I__1982\ : InMux
    port map (
            O => \N__11839\,
            I => \N__11836\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__11836\,
            I => \N__11832\
        );

    \I__1980\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11828\
        );

    \I__1979\ : Span4Mux_h
    port map (
            O => \N__11832\,
            I => \N__11825\
        );

    \I__1978\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11821\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__11828\,
            I => \N__11816\
        );

    \I__1976\ : Span4Mux_h
    port map (
            O => \N__11825\,
            I => \N__11816\
        );

    \I__1975\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11813\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__11821\,
            I => \c0.d_2_0\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__11816\,
            I => \c0.d_2_0\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__11813\,
            I => \c0.d_2_0\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__11806\,
            I => \c0.tx_data_RNO_3Z0Z_0_cascade_\
        );

    \I__1970\ : InMux
    port map (
            O => \N__11803\,
            I => \N__11800\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__11800\,
            I => \c0.tx_data_RNO_4Z0Z_0\
        );

    \I__1968\ : InMux
    port map (
            O => \N__11797\,
            I => \N__11791\
        );

    \I__1967\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11791\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__11791\,
            I => \N__11787\
        );

    \I__1965\ : InMux
    port map (
            O => \N__11790\,
            I => \N__11784\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__11787\,
            I => \c0.d_2_33\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__11784\,
            I => \c0.d_2_33\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__11779\,
            I => \N__11775\
        );

    \I__1961\ : InMux
    port map (
            O => \N__11778\,
            I => \N__11772\
        );

    \I__1960\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11769\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__11772\,
            I => \N__11766\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11763\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__11766\,
            I => \N__11757\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__11763\,
            I => \N__11757\
        );

    \I__1955\ : InMux
    port map (
            O => \N__11762\,
            I => \N__11754\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__11757\,
            I => \c0.d_2_34\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__11754\,
            I => \c0.d_2_34\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__11749\,
            I => \N__11745\
        );

    \I__1951\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11742\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11737\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__11742\,
            I => \N__11734\
        );

    \I__1948\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11731\
        );

    \I__1947\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11728\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__11737\,
            I => \N__11725\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__11734\,
            I => \N__11718\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__11731\,
            I => \N__11718\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__11728\,
            I => \N__11718\
        );

    \I__1942\ : Odrv12
    port map (
            O => \N__11725\,
            I => \c0.d_2_15\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__11718\,
            I => \c0.d_2_15\
        );

    \I__1940\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11707\
        );

    \I__1939\ : InMux
    port map (
            O => \N__11712\,
            I => \N__11704\
        );

    \I__1938\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11699\
        );

    \I__1937\ : InMux
    port map (
            O => \N__11710\,
            I => \N__11699\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__11707\,
            I => \N__11696\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11704\,
            I => \N__11693\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__11699\,
            I => \N__11690\
        );

    \I__1933\ : Span4Mux_h
    port map (
            O => \N__11696\,
            I => \N__11687\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__11693\,
            I => \N__11684\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__11690\,
            I => \N__11681\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__11687\,
            I => \c0.d_2_43\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__11684\,
            I => \c0.d_2_43\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__11681\,
            I => \c0.d_2_43\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__11674\,
            I => \c0.un105_newcrc_0_a2_0_cascade_\
        );

    \I__1926\ : InMux
    port map (
            O => \N__11671\,
            I => \N__11668\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__11668\,
            I => \N__11663\
        );

    \I__1924\ : InMux
    port map (
            O => \N__11667\,
            I => \N__11660\
        );

    \I__1923\ : InMux
    port map (
            O => \N__11666\,
            I => \N__11657\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__11663\,
            I => \c0.N_100\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__11660\,
            I => \c0.N_100\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__11657\,
            I => \c0.N_100\
        );

    \I__1919\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11646\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11642\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__11646\,
            I => \N__11639\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11635\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__11642\,
            I => \N__11630\
        );

    \I__1914\ : Span4Mux_h
    port map (
            O => \N__11639\,
            I => \N__11630\
        );

    \I__1913\ : InMux
    port map (
            O => \N__11638\,
            I => \N__11627\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__11635\,
            I => \c0.d_2_31\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__11630\,
            I => \c0.d_2_31\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__11627\,
            I => \c0.d_2_31\
        );

    \I__1909\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11617\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__11617\,
            I => \c0.un105_newcrc_0_a2_3\
        );

    \I__1907\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11611\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__11611\,
            I => \c0.tx_data_RNO_1Z0Z_5\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__11608\,
            I => \N__11605\
        );

    \I__1904\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11602\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__11602\,
            I => \c0.tx.r_Tx_DataZ0Z_5\
        );

    \I__1902\ : InMux
    port map (
            O => \N__11599\,
            I => \N__11595\
        );

    \I__1901\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11592\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__11595\,
            I => \N__11589\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__11592\,
            I => \N__11585\
        );

    \I__1898\ : Span4Mux_v
    port map (
            O => \N__11589\,
            I => \N__11582\
        );

    \I__1897\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11579\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__11585\,
            I => \c0.N_24_0\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__11582\,
            I => \c0.N_24_0\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__11579\,
            I => \c0.N_24_0\
        );

    \I__1893\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11569\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__11566\,
            I => \c0.un144_newcrc_2\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__11563\,
            I => \c0.un144_newcrc_5_cascade_\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__11560\,
            I => \N__11557\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11557\,
            I => \N__11554\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11554\,
            I => \c0.data_out_7_Z0Z_6\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11551\,
            I => \N__11548\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11548\,
            I => \c0.N_81\
        );

    \I__1884\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11542\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__11542\,
            I => \c0.data_out_6_Z0Z_6\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__11539\,
            I => \c0.tx_data_RNO_3Z0Z_4_cascade_\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11533\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11533\,
            I => \c0.tx_data_1_0_i_ns_1_4\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__11530\,
            I => \N__11526\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__11529\,
            I => \N__11523\
        );

    \I__1877\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11518\
        );

    \I__1876\ : InMux
    port map (
            O => \N__11523\,
            I => \N__11518\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__11518\,
            I => \N__11514\
        );

    \I__1874\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11510\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__11514\,
            I => \N__11507\
        );

    \I__1872\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11504\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__11510\,
            I => \c0.d_2_20\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__11507\,
            I => \c0.d_2_20\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__11504\,
            I => \c0.d_2_20\
        );

    \I__1868\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11494\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__11494\,
            I => \c0.tx_data_RNO_4Z0Z_4\
        );

    \I__1866\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11488\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__11488\,
            I => \c0.N_95\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__11485\,
            I => \c0.tx2_data_RNO_0Z0Z_2_cascade_\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11479\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__11479\,
            I => \N__11476\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__11476\,
            I => \N__11473\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__11473\,
            I => \c0.data_in_frame_6_Z0Z_2\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__11470\,
            I => \N__11467\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11467\,
            I => \N__11464\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__11464\,
            I => \N__11461\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__11461\,
            I => \c0.data_in_frame_7_Z0Z_2\
        );

    \I__1855\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11455\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__11455\,
            I => \c0.tx2_data_RNO_1Z0Z_2\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11449\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__11449\,
            I => \c0.tx_data_RNO_0Z0Z_3\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11446\,
            I => \N__11443\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__11443\,
            I => \c0.tx_data_1_0_i_ns_1_3\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11437\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__11434\,
            I => \c0.tx.r_Tx_DataZ0Z_3\
        );

    \I__1846\ : InMux
    port map (
            O => \N__11431\,
            I => \N__11428\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11428\,
            I => \N__11424\
        );

    \I__1844\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11421\
        );

    \I__1843\ : Odrv12
    port map (
            O => \N__11424\,
            I => \c0.d_2_7\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__11421\,
            I => \c0.d_2_7\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__11416\,
            I => \c0.tx_data_RNO_3Z0Z_7_cascade_\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11410\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__11410\,
            I => \c0.tx_data_RNO_4Z0Z_7\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__11407\,
            I => \c0.tx_data_1_0_i_ns_1_7_cascade_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11404\,
            I => \N__11401\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__11401\,
            I => \c0.tx.r_Tx_DataZ0Z_7\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__11398\,
            I => \N__11395\
        );

    \I__1834\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11392\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__11392\,
            I => \N__11389\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__11389\,
            I => \c0.tx.r_Tx_DataZ0Z_4\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11386\,
            I => \N__11382\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__11385\,
            I => \N__11378\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__11382\,
            I => \N__11375\
        );

    \I__1828\ : InMux
    port map (
            O => \N__11381\,
            I => \N__11372\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11369\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__11375\,
            I => \c0.data_in_7_Z0Z_3\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__11372\,
            I => \c0.data_in_7_Z0Z_3\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__11369\,
            I => \c0.data_in_7_Z0Z_3\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11357\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11354\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11351\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__11357\,
            I => \c0.data_in_2_Z0Z_1\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11354\,
            I => \c0.data_in_2_Z0Z_1\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__11351\,
            I => \c0.data_in_2_Z0Z_1\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11344\,
            I => \N__11341\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11341\,
            I => \N__11338\
        );

    \I__1815\ : Span4Mux_h
    port map (
            O => \N__11338\,
            I => \N__11333\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11337\,
            I => \N__11328\
        );

    \I__1813\ : InMux
    port map (
            O => \N__11336\,
            I => \N__11328\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__11333\,
            I => \c0.data_in_3_Z0Z_6\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__11328\,
            I => \c0.data_in_3_Z0Z_6\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__11323\,
            I => \N__11320\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11317\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__11317\,
            I => \N__11314\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__11314\,
            I => \c0.data_in_frame_7_Z0Z_3\
        );

    \I__1806\ : InMux
    port map (
            O => \N__11311\,
            I => \N__11307\
        );

    \I__1805\ : InMux
    port map (
            O => \N__11310\,
            I => \N__11304\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__11307\,
            I => \N__11298\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__11304\,
            I => \N__11298\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11303\,
            I => \N__11295\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__11298\,
            I => \c0.data_in_6_Z0Z_3\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__11295\,
            I => \c0.data_in_6_Z0Z_3\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11290\,
            I => \N__11287\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__11287\,
            I => \c0.data_in_frame_6_Z0Z_3\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__11284\,
            I => \N__11278\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11273\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11282\,
            I => \N__11273\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11268\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11268\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__11273\,
            I => \c0.d_4_17\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__11268\,
            I => \c0.d_4_17\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__11263\,
            I => \N__11260\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11260\,
            I => \N__11257\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11257\,
            I => \c0.tx2_data_RNO_4Z0Z_1\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__11254\,
            I => \c0.m161_ns_1_cascade_\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11248\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11248\,
            I => \c0.tx2_data_RNO_0Z0Z_1\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11242\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__11242\,
            I => \N__11238\
        );

    \I__1782\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11235\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__11238\,
            I => \c0.data_in_4_Z0Z_7\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11235\,
            I => \c0.data_in_4_Z0Z_7\
        );

    \I__1779\ : InMux
    port map (
            O => \N__11230\,
            I => \N__11227\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11227\,
            I => \N__11223\
        );

    \I__1777\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11220\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__11223\,
            I => \c0.data_in_5_Z0Z_3\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__11220\,
            I => \c0.data_in_5_Z0Z_3\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__11215\,
            I => \c0.N_108_cascade_\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__11212\,
            I => \c0.N_122_cascade_\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__11209\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_2_cascade_\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__11206\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_4_cascade_\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11203\,
            I => \N__11200\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__11200\,
            I => \N__11197\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__11197\,
            I => \N__11192\
        );

    \I__1767\ : InMux
    port map (
            O => \N__11196\,
            I => \N__11187\
        );

    \I__1766\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11187\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__11192\,
            I => \c0.data_in_2_Z0Z_4\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__11187\,
            I => \c0.data_in_2_Z0Z_4\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11182\,
            I => \N__11178\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11175\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__11178\,
            I => \c0.data_in_4_Z0Z_2\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__11175\,
            I => \c0.data_in_4_Z0Z_2\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11167\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__11167\,
            I => \N__11163\
        );

    \I__1757\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11160\
        );

    \I__1756\ : Span4Mux_h
    port map (
            O => \N__11163\,
            I => \N__11157\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__11160\,
            I => \N__11154\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__11157\,
            I => \c0.data_in_4_Z0Z_5\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__11154\,
            I => \c0.data_in_4_Z0Z_5\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11146\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__11146\,
            I => \N__11143\
        );

    \I__1750\ : Span4Mux_h
    port map (
            O => \N__11143\,
            I => \N__11139\
        );

    \I__1749\ : InMux
    port map (
            O => \N__11142\,
            I => \N__11136\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__11139\,
            I => \c0.data_in_0_Z0Z_0\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__11136\,
            I => \c0.data_in_0_Z0Z_0\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11128\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__11128\,
            I => \N__11124\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11127\,
            I => \N__11120\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__11124\,
            I => \N__11117\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11114\
        );

    \I__1741\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11111\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__11117\,
            I => \c0.data_in_1_Z0Z_3\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__11114\,
            I => \c0.data_in_1_Z0Z_3\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__11111\,
            I => \c0.data_in_1_Z0Z_3\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11101\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11101\,
            I => \N__11096\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11093\
        );

    \I__1734\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11090\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__11096\,
            I => \c0.data_in_1_Z0Z_7\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__11093\,
            I => \c0.data_in_1_Z0Z_7\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__11090\,
            I => \c0.data_in_1_Z0Z_7\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11080\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__11080\,
            I => \N__11076\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11079\,
            I => \N__11073\
        );

    \I__1727\ : Span4Mux_h
    port map (
            O => \N__11076\,
            I => \N__11069\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__11073\,
            I => \N__11066\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11072\,
            I => \N__11063\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__11069\,
            I => \c0.data_in_3_Z0Z_0\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__11066\,
            I => \c0.data_in_3_Z0Z_0\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11063\,
            I => \c0.data_in_3_Z0Z_0\
        );

    \I__1721\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11053\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__11053\,
            I => \N__11050\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__11050\,
            I => \N__11045\
        );

    \I__1718\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11042\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11039\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__11045\,
            I => \c0.data_in_3_Z0Z_5\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__11042\,
            I => \c0.data_in_3_Z0Z_5\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__11039\,
            I => \c0.data_in_3_Z0Z_5\
        );

    \I__1713\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11028\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11031\,
            I => \N__11025\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__11028\,
            I => \c0.data_in_4_Z0Z_1\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__11025\,
            I => \c0.data_in_4_Z0Z_1\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11020\,
            I => \N__11017\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11017\,
            I => \N__11014\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__11014\,
            I => \N__11009\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11013\,
            I => \N__11006\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11012\,
            I => \N__11003\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__11009\,
            I => \c0.data_in_2_Z0Z_5\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__11006\,
            I => \c0.data_in_2_Z0Z_5\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11003\,
            I => \c0.data_in_2_Z0Z_5\
        );

    \I__1701\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10993\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__10993\,
            I => \N__10988\
        );

    \I__1699\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10985\
        );

    \I__1698\ : InMux
    port map (
            O => \N__10991\,
            I => \N__10982\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__10988\,
            I => \c0.data_in_2_Z0Z_3\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__10985\,
            I => \c0.data_in_2_Z0Z_3\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__10982\,
            I => \c0.data_in_2_Z0Z_3\
        );

    \I__1694\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10972\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__10972\,
            I => \N__10969\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__10969\,
            I => \N__10965\
        );

    \I__1691\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10962\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__10965\,
            I => \c0.data_in_0_Z0Z_7\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__10962\,
            I => \c0.data_in_0_Z0Z_7\
        );

    \I__1688\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10953\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__10956\,
            I => \N__10949\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__10953\,
            I => \N__10946\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10943\
        );

    \I__1684\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10940\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__10946\,
            I => \c0.data_in_2_Z0Z_7\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__10943\,
            I => \c0.data_in_2_Z0Z_7\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__10940\,
            I => \c0.data_in_2_Z0Z_7\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__10933\,
            I => \N__10928\
        );

    \I__1679\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10925\
        );

    \I__1678\ : InMux
    port map (
            O => \N__10931\,
            I => \N__10922\
        );

    \I__1677\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10919\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__10925\,
            I => \c0.data_in_6_Z0Z_0\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__10922\,
            I => \c0.data_in_6_Z0Z_0\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__10919\,
            I => \c0.data_in_6_Z0Z_0\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__10912\,
            I => \c0.N_75_cascade_\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__10909\,
            I => \N__10906\
        );

    \I__1671\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10903\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__10903\,
            I => \c0.N_93\
        );

    \I__1669\ : InMux
    port map (
            O => \N__10900\,
            I => \N__10897\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__10897\,
            I => \N__10891\
        );

    \I__1667\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10888\
        );

    \I__1666\ : InMux
    port map (
            O => \N__10895\,
            I => \N__10885\
        );

    \I__1665\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10882\
        );

    \I__1664\ : Span4Mux_h
    port map (
            O => \N__10891\,
            I => \N__10875\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__10888\,
            I => \N__10875\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__10885\,
            I => \N__10875\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__10882\,
            I => \c0.d_2_35\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__10875\,
            I => \c0.d_2_35\
        );

    \I__1659\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10867\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__10867\,
            I => \N__10863\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__10866\,
            I => \N__10860\
        );

    \I__1656\ : Span12Mux_v
    port map (
            O => \N__10863\,
            I => \N__10857\
        );

    \I__1655\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10854\
        );

    \I__1654\ : Odrv12
    port map (
            O => \N__10857\,
            I => \c0.rx_data_7\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__10854\,
            I => \c0.rx_data_7\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__10849\,
            I => \c0.N_105_cascade_\
        );

    \I__1651\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10843\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10843\,
            I => \N__10840\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__10840\,
            I => \c0.data_out_6_Z0Z_5\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__10837\,
            I => \c0.nextCRC16_3_0_a2_1_15_cascade_\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10834\,
            I => \N__10830\
        );

    \I__1646\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10827\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__10830\,
            I => \c0.N_99\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__10827\,
            I => \c0.N_99\
        );

    \I__1643\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10819\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__10819\,
            I => \c0.nextCRC16_3_0_a2_5_15\
        );

    \I__1641\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10813\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__10813\,
            I => \c0.nextCRC16_3_0_a2_2_15\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__10810\,
            I => \c0.N_95_cascade_\
        );

    \I__1638\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10804\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__10804\,
            I => \N__10799\
        );

    \I__1636\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10794\
        );

    \I__1635\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10794\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__10799\,
            I => \c0.N_85\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__10794\,
            I => \c0.N_85\
        );

    \I__1632\ : InMux
    port map (
            O => \N__10789\,
            I => \N__10783\
        );

    \I__1631\ : InMux
    port map (
            O => \N__10788\,
            I => \N__10783\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__10783\,
            I => \c0.nextCRC16_3_2_1\
        );

    \I__1629\ : InMux
    port map (
            O => \N__10780\,
            I => \N__10777\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__10777\,
            I => \N__10773\
        );

    \I__1627\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10770\
        );

    \I__1626\ : Odrv12
    port map (
            O => \N__10773\,
            I => \c0.d_2_3\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__10770\,
            I => \c0.d_2_3\
        );

    \I__1624\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10762\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__10762\,
            I => \N__10758\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10755\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__10758\,
            I => \c0.N_75\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__10755\,
            I => \c0.N_75\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__10750\,
            I => \c0.nextCRC16_3_0_a2_1_2_cascade_\
        );

    \I__1618\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10744\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__10744\,
            I => \N__10741\
        );

    \I__1616\ : Span4Mux_h
    port map (
            O => \N__10741\,
            I => \N__10737\
        );

    \I__1615\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10734\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__10737\,
            I => \c0.dataZ0Z_6\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__10734\,
            I => \c0.dataZ0Z_6\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__10729\,
            I => \c0.N_99_cascade_\
        );

    \I__1611\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10723\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__10723\,
            I => \c0.nextCRC16_3_0_a2_0_0\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__10720\,
            I => \c0.nextCRC16_3_0_a2_3_0_cascade_\
        );

    \I__1608\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10714\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__10714\,
            I => \c0.nextCRC16_3_0_a2_4_0\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__10711\,
            I => \N__10707\
        );

    \I__1605\ : InMux
    port map (
            O => \N__10710\,
            I => \N__10704\
        );

    \I__1604\ : InMux
    port map (
            O => \N__10707\,
            I => \N__10701\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__10704\,
            I => \N__10698\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__1601\ : Span4Mux_h
    port map (
            O => \N__10698\,
            I => \N__10692\
        );

    \I__1600\ : Span4Mux_h
    port map (
            O => \N__10695\,
            I => \N__10689\
        );

    \I__1599\ : Span4Mux_h
    port map (
            O => \N__10692\,
            I => \N__10686\
        );

    \I__1598\ : Span4Mux_h
    port map (
            O => \N__10689\,
            I => \N__10683\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__10686\,
            I => \c0.d_2_27\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__10683\,
            I => \c0.d_2_27\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__10678\,
            I => \c0.N_81_cascade_\
        );

    \I__1594\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10669\
        );

    \I__1593\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10669\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__10669\,
            I => \c0.N_105\
        );

    \I__1591\ : SRMux
    port map (
            O => \N__10666\,
            I => \N__10663\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__10663\,
            I => \N__10660\
        );

    \I__1589\ : Span4Mux_h
    port map (
            O => \N__10660\,
            I => \N__10657\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__10657\,
            I => \c0.tx.N_390_i\
        );

    \I__1587\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10642\
        );

    \I__1586\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10642\
        );

    \I__1585\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10635\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10635\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10635\
        );

    \I__1582\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10628\
        );

    \I__1581\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10628\
        );

    \I__1580\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10628\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__10642\,
            I => \N__10623\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__10635\,
            I => \N__10623\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__10628\,
            I => \c0.tx.r_SM_Main_dup_2\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__10623\,
            I => \c0.tx.r_SM_Main_dup_2\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__10618\,
            I => \N__10615\
        );

    \I__1574\ : InMux
    port map (
            O => \N__10615\,
            I => \N__10612\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__10612\,
            I => \N__10609\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__10609\,
            I => \c0.tx.r_SM_Main_recr_i_0_a2_0_2_0_1_3\
        );

    \I__1571\ : InMux
    port map (
            O => \N__10606\,
            I => \N__10596\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10605\,
            I => \N__10593\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10584\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10603\,
            I => \N__10584\
        );

    \I__1567\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10584\
        );

    \I__1566\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10584\
        );

    \I__1565\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10579\
        );

    \I__1564\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10579\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__10596\,
            I => \c0.tx.r_Bit_IndexZ0Z_1\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10593\,
            I => \c0.tx.r_Bit_IndexZ0Z_1\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__10584\,
            I => \c0.tx.r_Bit_IndexZ0Z_1\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__10579\,
            I => \c0.tx.r_Bit_IndexZ0Z_1\
        );

    \I__1559\ : InMux
    port map (
            O => \N__10570\,
            I => \N__10563\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10569\,
            I => \N__10556\
        );

    \I__1557\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10556\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10567\,
            I => \N__10556\
        );

    \I__1555\ : InMux
    port map (
            O => \N__10566\,
            I => \N__10553\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__10563\,
            I => \c0.tx.r_Bit_IndexZ0Z_2\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__10556\,
            I => \c0.tx.r_Bit_IndexZ0Z_2\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__10553\,
            I => \c0.tx.r_Bit_IndexZ0Z_2\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__10546\,
            I => \N__10543\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10540\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__10540\,
            I => \N__10534\
        );

    \I__1548\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10531\
        );

    \I__1547\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10524\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10537\,
            I => \N__10524\
        );

    \I__1545\ : Span4Mux_h
    port map (
            O => \N__10534\,
            I => \N__10521\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__10531\,
            I => \N__10518\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10513\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10513\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__10524\,
            I => \c0.tx.r_SM_Main_dup_1\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__10521\,
            I => \c0.tx.r_SM_Main_dup_1\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__10518\,
            I => \c0.tx.r_SM_Main_dup_1\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__10513\,
            I => \c0.tx.r_SM_Main_dup_1\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__10504\,
            I => \N__10499\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__10503\,
            I => \N__10495\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10502\,
            I => \N__10487\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10487\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10487\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10481\
        );

    \I__1531\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10481\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__10487\,
            I => \N__10478\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10475\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__10481\,
            I => \c0.tx.r_Bit_IndexZ0Z_0\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__10478\,
            I => \c0.tx.r_Bit_IndexZ0Z_0\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__10475\,
            I => \c0.tx.r_Bit_IndexZ0Z_0\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10465\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10462\
        );

    \I__1523\ : Odrv4
    port map (
            O => \N__10462\,
            I => \c0.tx.r_SM_Main_recr_i_i_a2_0_1_2\
        );

    \I__1522\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10456\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__10456\,
            I => \c0.data_out_7_Z0Z_5\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__10453\,
            I => \c0.tx_data_RNO_3Z0Z_3_cascade_\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10450\,
            I => \N__10447\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10441\
        );

    \I__1517\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10441\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__10441\,
            I => \N__10437\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10434\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__10437\,
            I => \N__10429\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__10434\,
            I => \N__10429\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__10429\,
            I => \c0.d_2_19\
        );

    \I__1511\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10423\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__10423\,
            I => \c0.tx_data_RNO_4Z0Z_3\
        );

    \I__1509\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10417\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__10417\,
            I => \N__10414\
        );

    \I__1507\ : Span4Mux_h
    port map (
            O => \N__10414\,
            I => \N__10410\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10407\
        );

    \I__1505\ : Odrv4
    port map (
            O => \N__10410\,
            I => \c0.rx_data_0\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__10407\,
            I => \c0.rx_data_0\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__10402\,
            I => \c0.tx.o_Tx_Serial_2_3_i_m2_ns_1_cascade_\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10394\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10391\
        );

    \I__1500\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10388\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10394\,
            I => \c0.tx.N_90_ip_RNI1U1EZ0\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10391\,
            I => \c0.tx.N_90_ip_RNI1U1EZ0\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__10388\,
            I => \c0.tx.N_90_ip_RNI1U1EZ0\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__10381\,
            I => \c0.tx.o_Tx_Serial_2_6_i_m2_ns_1_cascade_\
        );

    \I__1495\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10375\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__10375\,
            I => \c0.tx.o_Tx_Serial_RNO_3_0\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__10372\,
            I => \c0.tx.o_Tx_Serial_RNO_2_0_cascade_\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__10369\,
            I => \N__10364\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__10368\,
            I => \N__10361\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__10367\,
            I => \N__10357\
        );

    \I__1489\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10347\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10347\
        );

    \I__1487\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10347\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10347\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10344\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__10347\,
            I => \N__10341\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__10344\,
            I => \N__10338\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__10341\,
            I => \N__10335\
        );

    \I__1481\ : Span4Mux_h
    port map (
            O => \N__10338\,
            I => \N__10332\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__10335\,
            I => \c0.tx.r_SM_Main_RNI522EZ0Z_4\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__10332\,
            I => \c0.tx.r_SM_Main_RNI522EZ0Z_4\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__10327\,
            I => \c0.tx.o_Tx_Serial_RNOZ0Z_1_cascade_\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10320\
        );

    \I__1476\ : InMux
    port map (
            O => \N__10323\,
            I => \N__10313\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__10320\,
            I => \N__10310\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10307\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10304\
        );

    \I__1472\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10299\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10299\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__10313\,
            I => \c0.tx.r_SM_Main_dup_3\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__10310\,
            I => \c0.tx.r_SM_Main_dup_3\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__10307\,
            I => \c0.tx.r_SM_Main_dup_3\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10304\,
            I => \c0.tx.r_SM_Main_dup_3\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__10299\,
            I => \c0.tx.r_SM_Main_dup_3\
        );

    \I__1465\ : IoInMux
    port map (
            O => \N__10288\,
            I => \N__10285\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__10285\,
            I => \N__10282\
        );

    \I__1463\ : IoSpan4Mux
    port map (
            O => \N__10282\,
            I => \N__10279\
        );

    \I__1462\ : IoSpan4Mux
    port map (
            O => \N__10279\,
            I => \N__10276\
        );

    \I__1461\ : Span4Mux_s3_h
    port map (
            O => \N__10276\,
            I => \N__10273\
        );

    \I__1460\ : Span4Mux_h
    port map (
            O => \N__10273\,
            I => \N__10269\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10266\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__10269\,
            I => \PIN_1_c\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__10266\,
            I => \PIN_1_c\
        );

    \I__1456\ : InMux
    port map (
            O => \N__10261\,
            I => \N__10258\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__10258\,
            I => \N__10255\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__10255\,
            I => \N__10251\
        );

    \I__1453\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10248\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__10251\,
            I => \c0.data_in_0_Z0Z_4\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10248\,
            I => \c0.data_in_0_Z0Z_4\
        );

    \I__1450\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10238\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10235\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10232\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__10238\,
            I => \c0.data_in_1_Z0Z_0\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__10235\,
            I => \c0.data_in_1_Z0Z_0\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__10232\,
            I => \c0.data_in_1_Z0Z_0\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10222\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__10222\,
            I => \N__10219\
        );

    \I__1442\ : Span12Mux_v
    port map (
            O => \N__10219\,
            I => \N__10215\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10218\,
            I => \N__10212\
        );

    \I__1440\ : Odrv12
    port map (
            O => \N__10215\,
            I => \c0.rx_data_3\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__10212\,
            I => \c0.rx_data_3\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10204\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__10204\,
            I => \N__10200\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__10203\,
            I => \N__10197\
        );

    \I__1435\ : Span12Mux_v
    port map (
            O => \N__10200\,
            I => \N__10194\
        );

    \I__1434\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10191\
        );

    \I__1433\ : Odrv12
    port map (
            O => \N__10194\,
            I => \c0.rx_data_1\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10191\,
            I => \c0.rx_data_1\
        );

    \I__1431\ : InMux
    port map (
            O => \N__10186\,
            I => \N__10182\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10179\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10182\,
            I => \c0.dataZ0Z_0\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__10179\,
            I => \c0.dataZ0Z_0\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10170\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10167\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__10170\,
            I => \c0.dataZ0Z_14\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__10167\,
            I => \c0.dataZ0Z_14\
        );

    \I__1423\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10158\
        );

    \I__1422\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10155\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__10158\,
            I => \c0.dataZ0Z_11\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10155\,
            I => \c0.dataZ0Z_11\
        );

    \I__1419\ : InMux
    port map (
            O => \N__10150\,
            I => \N__10146\
        );

    \I__1418\ : InMux
    port map (
            O => \N__10149\,
            I => \N__10143\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__10146\,
            I => \c0.dataZ0Z_2\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__10143\,
            I => \c0.dataZ0Z_2\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10134\
        );

    \I__1414\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10131\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__10134\,
            I => \c0.dataZ0Z_15\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__10131\,
            I => \c0.dataZ0Z_15\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10122\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10119\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__10122\,
            I => \c0.dataZ0Z_4\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__10119\,
            I => \c0.dataZ0Z_4\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10110\
        );

    \I__1406\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10107\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__10110\,
            I => \c0.dataZ0Z_8\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__10107\,
            I => \c0.dataZ0Z_8\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10099\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__10099\,
            I => \c0.nextCRC16_3_0_a2_6_0_15\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__10096\,
            I => \c0.nextCRC16_3_9_cascade_\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__10093\,
            I => \c0.N_106_cascade_\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10087\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__10087\,
            I => \N__10084\
        );

    \I__1397\ : Span12Mux_v
    port map (
            O => \N__10084\,
            I => \N__10080\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10077\
        );

    \I__1395\ : Odrv12
    port map (
            O => \N__10080\,
            I => \c0.N_92\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__10077\,
            I => \c0.N_92\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10066\
        );

    \I__1392\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10066\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__10066\,
            I => \c0.N_106\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10063\,
            I => \N__10060\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10057\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__10057\,
            I => \c0.data_out_7_Z0Z_0\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__10054\,
            I => \N__10051\
        );

    \I__1386\ : InMux
    port map (
            O => \N__10051\,
            I => \N__10048\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__10048\,
            I => \N__10045\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__10045\,
            I => \c0.nextCRC16_3_0_a2_0_10\
        );

    \I__1383\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10039\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__10039\,
            I => \N__10035\
        );

    \I__1381\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10032\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__10035\,
            I => \c0.dataZ0Z_12\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__10032\,
            I => \c0.dataZ0Z_12\
        );

    \I__1378\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10024\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10024\,
            I => \N__10019\
        );

    \I__1376\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10016\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10013\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__10019\,
            I => \c0.N_77\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__10016\,
            I => \c0.N_77\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__10013\,
            I => \c0.N_77\
        );

    \I__1371\ : InMux
    port map (
            O => \N__10006\,
            I => \N__10002\
        );

    \I__1370\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9999\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__10002\,
            I => \N__9993\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__9999\,
            I => \N__9993\
        );

    \I__1367\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9990\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__9993\,
            I => \c0.N_76\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__9990\,
            I => \c0.N_76\
        );

    \I__1364\ : InMux
    port map (
            O => \N__9985\,
            I => \N__9981\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__9984\,
            I => \N__9976\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__9981\,
            I => \N__9973\
        );

    \I__1361\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9970\
        );

    \I__1360\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9965\
        );

    \I__1359\ : InMux
    port map (
            O => \N__9976\,
            I => \N__9965\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__9973\,
            I => \c0.tx.r_SM_Main_dup_4\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__9970\,
            I => \c0.tx.r_SM_Main_dup_4\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__9965\,
            I => \c0.tx.r_SM_Main_dup_4\
        );

    \I__1355\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9954\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__9957\,
            I => \N__9951\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__9954\,
            I => \N__9948\
        );

    \I__1352\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9944\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__9948\,
            I => \N__9941\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__9947\,
            I => \N__9937\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__9944\,
            I => \N__9933\
        );

    \I__1348\ : Span4Mux_h
    port map (
            O => \N__9941\,
            I => \N__9930\
        );

    \I__1347\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9927\
        );

    \I__1346\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9922\
        );

    \I__1345\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9922\
        );

    \I__1344\ : Odrv4
    port map (
            O => \N__9933\,
            I => \c0.tx_transmitZ0\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__9930\,
            I => \c0.tx_transmitZ0\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__9927\,
            I => \c0.tx_transmitZ0\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__9922\,
            I => \c0.tx_transmitZ0\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__9913\,
            I => \N__9910\
        );

    \I__1339\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9907\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__9907\,
            I => \c0.tx.r_SM_Main_RNO_0Z0Z_0\
        );

    \I__1337\ : InMux
    port map (
            O => \N__9904\,
            I => \N__9898\
        );

    \I__1336\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9891\
        );

    \I__1335\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9891\
        );

    \I__1334\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9891\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__9898\,
            I => \c0.tx.N_171_0\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__9891\,
            I => \c0.tx.N_171_0\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__9886\,
            I => \c0.tx.r_SM_Main_RNO_0Z0Z_2_cascade_\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__9883\,
            I => \N__9880\
        );

    \I__1329\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9873\
        );

    \I__1328\ : InMux
    port map (
            O => \N__9879\,
            I => \N__9864\
        );

    \I__1327\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9864\
        );

    \I__1326\ : InMux
    port map (
            O => \N__9877\,
            I => \N__9864\
        );

    \I__1325\ : InMux
    port map (
            O => \N__9876\,
            I => \N__9864\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__9873\,
            I => \N__9858\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9858\
        );

    \I__1322\ : InMux
    port map (
            O => \N__9863\,
            I => \N__9849\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__9858\,
            I => \N__9846\
        );

    \I__1320\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9841\
        );

    \I__1319\ : InMux
    port map (
            O => \N__9856\,
            I => \N__9841\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9832\
        );

    \I__1317\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9832\
        );

    \I__1316\ : InMux
    port map (
            O => \N__9853\,
            I => \N__9832\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9852\,
            I => \N__9832\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__9849\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__9846\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__9841\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__9832\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__9823\,
            I => \N__9811\
        );

    \I__1309\ : InMux
    port map (
            O => \N__9822\,
            I => \N__9808\
        );

    \I__1308\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9803\
        );

    \I__1307\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9803\
        );

    \I__1306\ : InMux
    port map (
            O => \N__9819\,
            I => \N__9796\
        );

    \I__1305\ : InMux
    port map (
            O => \N__9818\,
            I => \N__9796\
        );

    \I__1304\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9796\
        );

    \I__1303\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9787\
        );

    \I__1302\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9787\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9814\,
            I => \N__9787\
        );

    \I__1300\ : InMux
    port map (
            O => \N__9811\,
            I => \N__9787\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__9808\,
            I => \c0.tx.N_90_dup\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__9803\,
            I => \c0.tx.N_90_dup\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__9796\,
            I => \c0.tx.N_90_dup\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__9787\,
            I => \c0.tx.N_90_dup\
        );

    \I__1295\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9775\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__9775\,
            I => \N__9772\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__9772\,
            I => \N__9763\
        );

    \I__1292\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9760\
        );

    \I__1291\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9757\
        );

    \I__1290\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9748\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9748\
        );

    \I__1288\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9748\
        );

    \I__1287\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9748\
        );

    \I__1286\ : Sp12to4
    port map (
            O => \N__9763\,
            I => \N__9741\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__9760\,
            I => \N__9741\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__9757\,
            I => \N__9741\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__9748\,
            I => \c0.tx.r_Clock_Count12_THRU_CO\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__9741\,
            I => \c0.tx.r_Clock_Count12_THRU_CO\
        );

    \I__1281\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9729\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9729\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9726\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__9729\,
            I => \c0.tx.r_SM_Main_RNIVDI71Z0Z_2\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__9726\,
            I => \c0.tx.r_SM_Main_RNIVDI71Z0Z_2\
        );

    \I__1276\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9718\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__9718\,
            I => \c0.i12_4_and\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__9715\,
            I => \c0.tx.r_Bit_Index_RNO_0Z0Z_2_cascade_\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__9712\,
            I => \c0.tx.r_Tx_Active_1_sqmuxa_cascade_\
        );

    \I__1272\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9706\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__9706\,
            I => \c0.tx.N_90_ip_RNIVJLQZ0\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9694\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9694\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9694\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__9694\,
            I => \c0.tx_active\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__9691\,
            I => \c0.tx.N_90_ip_RNI1U1EZ0_cascade_\
        );

    \I__1265\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9685\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9685\,
            I => \c0.i12_5_and\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9679\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__9679\,
            I => \c0.i12_6_and\
        );

    \I__1261\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9673\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9673\,
            I => \c0.i12_2_and\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9670\,
            I => \c0.data_cry_10\
        );

    \I__1258\ : InMux
    port map (
            O => \N__9667\,
            I => \c0.data_cry_11\
        );

    \I__1257\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__9661\,
            I => \N__9657\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9654\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__9657\,
            I => \c0.dataZ0Z_13\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__9654\,
            I => \c0.dataZ0Z_13\
        );

    \I__1252\ : InMux
    port map (
            O => \N__9649\,
            I => \c0.data_cry_12\
        );

    \I__1251\ : InMux
    port map (
            O => \N__9646\,
            I => \c0.data_cry_13\
        );

    \I__1250\ : InMux
    port map (
            O => \N__9643\,
            I => \c0.data_cry_14\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9637\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__9637\,
            I => \c0.i12_3_and\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9634\,
            I => \c0.data_cry_1\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9628\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__9628\,
            I => \N__9624\
        );

    \I__1244\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9621\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__9624\,
            I => \c0.dataZ0Z_3\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__9621\,
            I => \c0.dataZ0Z_3\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9616\,
            I => \c0.data_cry_2\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9613\,
            I => \c0.data_cry_3\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9607\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__9607\,
            I => \N__9603\
        );

    \I__1237\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9600\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__9603\,
            I => \c0.dataZ0Z_5\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__9600\,
            I => \c0.dataZ0Z_5\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9595\,
            I => \c0.data_cry_4\
        );

    \I__1233\ : InMux
    port map (
            O => \N__9592\,
            I => \c0.data_cry_5\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9585\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9582\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__9585\,
            I => \c0.dataZ0Z_7\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__9582\,
            I => \c0.dataZ0Z_7\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9577\,
            I => \c0.data_cry_6\
        );

    \I__1227\ : InMux
    port map (
            O => \N__9574\,
            I => \bfn_9_28_0_\
        );

    \I__1226\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9568\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__9568\,
            I => \N__9564\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9561\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__9564\,
            I => \c0.dataZ0Z_9\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__9561\,
            I => \c0.dataZ0Z_9\
        );

    \I__1221\ : InMux
    port map (
            O => \N__9556\,
            I => \c0.data_cry_8\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9550\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__9550\,
            I => \N__9546\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9543\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__9546\,
            I => \c0.dataZ0Z_10\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__9543\,
            I => \c0.dataZ0Z_10\
        );

    \I__1215\ : InMux
    port map (
            O => \N__9538\,
            I => \c0.data_cry_9\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9535\,
            I => \bfn_9_27_0_\
        );

    \I__1213\ : InMux
    port map (
            O => \N__9532\,
            I => \N__9528\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9531\,
            I => \N__9525\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__9528\,
            I => \c0.dataZ0Z_1\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__9525\,
            I => \c0.dataZ0Z_1\
        );

    \I__1209\ : InMux
    port map (
            O => \N__9520\,
            I => \c0.data_cry_0\
        );

    \I__1208\ : InMux
    port map (
            O => \N__9517\,
            I => \N__9514\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__9514\,
            I => \N__9511\
        );

    \I__1206\ : Odrv12
    port map (
            O => \N__9511\,
            I => \c0.tx.r_Clock_Count_RNO_0Z0Z_2\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9508\,
            I => \c0.tx.un1_r_Clock_Count_cry_1\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9505\,
            I => \c0.tx.un1_r_Clock_Count_cry_2\
        );

    \I__1203\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9499\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9496\
        );

    \I__1201\ : Odrv12
    port map (
            O => \N__9496\,
            I => \c0.tx.r_Clock_Count_RNO_0Z0Z_3\
        );

    \I__1200\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9489\
        );

    \I__1199\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9486\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__9489\,
            I => \N__9480\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__9486\,
            I => \N__9480\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9477\
        );

    \I__1195\ : Odrv12
    port map (
            O => \N__9480\,
            I => \c0.tx.r_Clock_CountZ0Z_2\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__9477\,
            I => \c0.tx.r_Clock_CountZ0Z_2\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9468\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9465\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__9468\,
            I => \N__9459\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9459\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9464\,
            I => \N__9456\
        );

    \I__1188\ : Odrv12
    port map (
            O => \N__9459\,
            I => \c0.tx.r_Clock_CountZ0Z_1\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9456\,
            I => \c0.tx.r_Clock_CountZ0Z_1\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__9451\,
            I => \N__9447\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9442\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9447\,
            I => \N__9442\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__9442\,
            I => \N__9439\
        );

    \I__1182\ : Span4Mux_h
    port map (
            O => \N__9439\,
            I => \N__9435\
        );

    \I__1181\ : InMux
    port map (
            O => \N__9438\,
            I => \N__9432\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__9435\,
            I => \c0.tx.r_Clock_CountZ0Z_3\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__9432\,
            I => \c0.tx.r_Clock_CountZ0Z_3\
        );

    \I__1178\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9421\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9421\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9421\,
            I => \N__9417\
        );

    \I__1175\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9414\
        );

    \I__1174\ : Odrv12
    port map (
            O => \N__9417\,
            I => \c0.tx.r_Clock_CountZ0Z_0\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__9414\,
            I => \c0.tx.r_Clock_CountZ0Z_0\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9406\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__9406\,
            I => \N__9403\
        );

    \I__1170\ : Span4Mux_h
    port map (
            O => \N__9403\,
            I => \N__9400\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__9400\,
            I => \c0.tx.r_SM_Main_RNO_0Z0Z_1\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__9397\,
            I => \c0.tx.N_171_0_cascade_\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__9394\,
            I => \c0.nextCRC16_3_0_a2_1_8_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9388\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__9388\,
            I => \c0.data_out_6_Z0Z_0\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__9385\,
            I => \N__9382\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9379\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__9379\,
            I => \N__9376\
        );

    \I__1161\ : Span12Mux_v
    port map (
            O => \N__9376\,
            I => \N__9373\
        );

    \I__1160\ : Odrv12
    port map (
            O => \N__9373\,
            I => \c0.N_71\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__9370\,
            I => \c0.tx.N_90_ip_RNIVJLQZ0_cascade_\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9364\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__9364\,
            I => \c0.tx.r_SM_Main_illegal_0\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__9361\,
            I => \c0.tx.N_90_dup_cascade_\
        );

    \I__1155\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9355\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__9355\,
            I => \c0.tx.N_83_0\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9348\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__9351\,
            I => \N__9345\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9348\,
            I => \N__9342\
        );

    \I__1150\ : InMux
    port map (
            O => \N__9345\,
            I => \N__9339\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__9342\,
            I => \c0.tx.r_Clock_Count_0_sqmuxa\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__9339\,
            I => \c0.tx.r_Clock_Count_0_sqmuxa\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9331\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9331\,
            I => \N__9328\
        );

    \I__1145\ : Span4Mux_h
    port map (
            O => \N__9328\,
            I => \N__9325\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__9325\,
            I => \c0.tx.r_Clock_Count_RNO_0Z0Z_0\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9319\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9319\,
            I => \N__9316\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__9316\,
            I => \N__9313\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__9313\,
            I => \c0.tx.r_Clock_Count_RNO_0Z0Z_1\
        );

    \I__1139\ : InMux
    port map (
            O => \N__9310\,
            I => \c0.tx.un1_r_Clock_Count_cry_0\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9307\,
            I => \N__9304\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9304\,
            I => \c0.i12_1_and\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9298\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__9298\,
            I => \N__9295\
        );

    \I__1134\ : Span4Mux_v
    port map (
            O => \N__9295\,
            I => \N__9291\
        );

    \I__1133\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9288\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__9291\,
            I => \blink_counterZ0Z_21\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9288\,
            I => \blink_counterZ0Z_21\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9277\
        );

    \I__1129\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9277\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__9277\,
            I => \N__9274\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__9274\,
            I => \N__9270\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9267\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__9270\,
            I => \blink_counterZ0Z_22\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9267\,
            I => \blink_counterZ0Z_22\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__9262\,
            I => \N__9259\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9253\
        );

    \I__1121\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9253\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__9253\,
            I => \N__9250\
        );

    \I__1119\ : Span4Mux_v
    port map (
            O => \N__9250\,
            I => \N__9246\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9243\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__9246\,
            I => \blink_counterZ0Z_24\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__9243\,
            I => \blink_counterZ0Z_24\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__9235\,
            I => \N_12\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9226\
        );

    \I__1112\ : InMux
    port map (
            O => \N__9231\,
            I => \N__9226\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__1110\ : Span4Mux_v
    port map (
            O => \N__9223\,
            I => \N__9219\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9216\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__9219\,
            I => \blink_counterZ0Z_25\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9216\,
            I => \blink_counterZ0Z_25\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__9211\,
            I => \N_8_0_cascade_\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9205\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__9205\,
            I => \N__9202\
        );

    \I__1103\ : Span4Mux_h
    port map (
            O => \N__9202\,
            I => \N__9198\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9201\,
            I => \N__9195\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__9198\,
            I => \blink_counterZ0Z_23\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__9195\,
            I => \blink_counterZ0Z_23\
        );

    \I__1099\ : IoInMux
    port map (
            O => \N__9190\,
            I => \N__9187\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__1097\ : Span4Mux_s1_h
    port map (
            O => \N__9184\,
            I => \N__9181\
        );

    \I__1096\ : Sp12to4
    port map (
            O => \N__9181\,
            I => \N__9178\
        );

    \I__1095\ : Span12Mux_s11_v
    port map (
            O => \N__9178\,
            I => \N__9175\
        );

    \I__1094\ : Odrv12
    port map (
            O => \N__9175\,
            I => \LED_c\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__9172\,
            I => \N__9169\
        );

    \I__1092\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9166\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9166\,
            I => \c0.i12_7_and\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9163\,
            I => \bfn_9_20_0_\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9157\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9157\,
            I => \c0.i12_0_and\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__9154\,
            I => \N__9151\
        );

    \I__1086\ : InMux
    port map (
            O => \N__9151\,
            I => \N__9148\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__9148\,
            I => \c0.rx.r_SM_Main_ns_0_i_a2_1_0_2\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9137\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9132\
        );

    \I__1082\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9132\
        );

    \I__1081\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9125\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9125\
        );

    \I__1079\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9125\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__9137\,
            I => \c0.rx.r_SM_Main_dup_1\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__9132\,
            I => \c0.rx.r_SM_Main_dup_1\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__9125\,
            I => \c0.rx.r_SM_Main_dup_1\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__9118\,
            I => \c0.rx.un1_r_Rx_DV7_i_0_cascade_\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9112\,
            I => \N__9109\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__9106\,
            I => \c0.rx.r_Rx_DV_RNOZ0Z_0\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9097\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9097\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__9097\,
            I => \N__9088\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9081\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9081\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9081\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9074\
        );

    \I__1063\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9074\
        );

    \I__1062\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9074\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__9088\,
            I => \c0.rx.r_SM_Main_dup_2\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__9081\,
            I => \c0.rx.r_SM_Main_dup_2\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__9074\,
            I => \c0.rx.r_SM_Main_dup_2\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9064\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__9064\,
            I => \c0.rx.r_SM_Main_ns_0_i_0_0_2\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9061\,
            I => \N__9057\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9060\,
            I => \N__9054\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9039\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9054\,
            I => \N__9039\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9036\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9033\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9028\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9028\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9049\,
            I => \N__9025\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9022\
        );

    \I__1046\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9019\
        );

    \I__1045\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9016\
        );

    \I__1044\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9013\
        );

    \I__1043\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9010\
        );

    \I__1042\ : Span4Mux_v
    port map (
            O => \N__9039\,
            I => \N__9005\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__9036\,
            I => \N__9005\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__9033\,
            I => \N__8990\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__9028\,
            I => \N__8990\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9025\,
            I => \N__8990\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9022\,
            I => \N__8990\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__9019\,
            I => \N__8990\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__9016\,
            I => \N__8990\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9013\,
            I => \N__8990\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__8987\
        );

    \I__1032\ : Span4Mux_h
    port map (
            O => \N__9005\,
            I => \N__8984\
        );

    \I__1031\ : Span4Mux_v
    port map (
            O => \N__8990\,
            I => \N__8981\
        );

    \I__1030\ : Span4Mux_h
    port map (
            O => \N__8987\,
            I => \N__8976\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__8984\,
            I => \N__8976\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__8981\,
            I => \c0.rx.r_Rx_DataZ0\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__8976\,
            I => \c0.rx.r_Rx_DataZ0\
        );

    \I__1026\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8966\
        );

    \I__1025\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8963\
        );

    \I__1024\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8960\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8957\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__8963\,
            I => \c0.rx.N_383\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__8960\,
            I => \c0.rx.N_383\
        );

    \I__1020\ : Odrv4
    port map (
            O => \N__8957\,
            I => \c0.rx.N_383\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8947\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__8947\,
            I => \N__8940\
        );

    \I__1017\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8937\
        );

    \I__1016\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8930\
        );

    \I__1015\ : InMux
    port map (
            O => \N__8944\,
            I => \N__8930\
        );

    \I__1014\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8930\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__8940\,
            I => \c0.rx.N_321\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__8937\,
            I => \c0.rx.N_321\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__8930\,
            I => \c0.rx.N_321\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__8923\,
            I => \c0.rx.r_Clock_Count_8_f0_0_a2_0_0_2_cascade_\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__8920\,
            I => \N__8916\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__8919\,
            I => \N__8913\
        );

    \I__1007\ : InMux
    port map (
            O => \N__8916\,
            I => \N__8909\
        );

    \I__1006\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8906\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8903\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__8909\,
            I => \N__8898\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__8906\,
            I => \N__8898\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__8903\,
            I => \N__8893\
        );

    \I__1001\ : Span4Mux_h
    port map (
            O => \N__8898\,
            I => \N__8893\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__8893\,
            I => \c0.rx.N_371\
        );

    \I__999\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8887\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__8887\,
            I => \N__8878\
        );

    \I__997\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8869\
        );

    \I__996\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8869\
        );

    \I__995\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8869\
        );

    \I__994\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8869\
        );

    \I__993\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8866\
        );

    \I__992\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8863\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__8878\,
            I => \c0.rx.N_332\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__8869\,
            I => \c0.rx.N_332\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__8866\,
            I => \c0.rx.N_332\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__8863\,
            I => \c0.rx.N_332\
        );

    \I__987\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8851\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__8851\,
            I => \N__8844\
        );

    \I__985\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8841\
        );

    \I__984\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8838\
        );

    \I__983\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8835\
        );

    \I__982\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8826\
        );

    \I__981\ : Span4Mux_v
    port map (
            O => \N__8844\,
            I => \N__8821\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__8841\,
            I => \N__8821\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__8838\,
            I => \N__8818\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__8835\,
            I => \N__8815\
        );

    \I__977\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8810\
        );

    \I__976\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8810\
        );

    \I__975\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8801\
        );

    \I__974\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8801\
        );

    \I__973\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8801\
        );

    \I__972\ : InMux
    port map (
            O => \N__8829\,
            I => \N__8801\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__8826\,
            I => \c0.rx.r_SM_Main_RNI58REZ0Z_0\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__8821\,
            I => \c0.rx.r_SM_Main_RNI58REZ0Z_0\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__8818\,
            I => \c0.rx.r_SM_Main_RNI58REZ0Z_0\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__8815\,
            I => \c0.rx.r_SM_Main_RNI58REZ0Z_0\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__8810\,
            I => \c0.rx.r_SM_Main_RNI58REZ0Z_0\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__8801\,
            I => \c0.rx.r_SM_Main_RNI58REZ0Z_0\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__8788\,
            I => \N__8783\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__8787\,
            I => \N__8780\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__8786\,
            I => \N__8776\
        );

    \I__962\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8770\
        );

    \I__961\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8770\
        );

    \I__960\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8767\
        );

    \I__959\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8764\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__8775\,
            I => \N__8761\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8754\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__8767\,
            I => \N__8754\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__8764\,
            I => \N__8754\
        );

    \I__954\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8751\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__8754\,
            I => \c0.rx.N_361\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__8751\,
            I => \c0.rx.N_361\
        );

    \I__951\ : InMux
    port map (
            O => \N__8746\,
            I => \N__8743\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__8743\,
            I => \N__8740\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__8740\,
            I => \c0.rx.r_Clock_Count_RNO_0_0_3\
        );

    \I__948\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8731\
        );

    \I__947\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8728\
        );

    \I__946\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8723\
        );

    \I__945\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8723\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__8731\,
            I => \N__8720\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__8728\,
            I => \N__8715\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__8723\,
            I => \N__8715\
        );

    \I__941\ : Odrv12
    port map (
            O => \N__8720\,
            I => \c0.rx.r_Clock_CountZ1Z_3\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__8715\,
            I => \c0.rx.r_Clock_CountZ1Z_3\
        );

    \I__939\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8700\
        );

    \I__938\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8700\
        );

    \I__937\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8697\
        );

    \I__936\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8690\
        );

    \I__935\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8690\
        );

    \I__934\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8690\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__8700\,
            I => \N__8687\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__8697\,
            I => \N__8682\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8690\,
            I => \N__8682\
        );

    \I__930\ : Odrv4
    port map (
            O => \N__8687\,
            I => \c0.rx.N_386\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__8682\,
            I => \c0.rx.N_386\
        );

    \I__928\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8669\
        );

    \I__927\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8662\
        );

    \I__926\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8662\
        );

    \I__925\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8662\
        );

    \I__924\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8657\
        );

    \I__923\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8657\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__8669\,
            I => \c0.rx.r_SM_Main_dup_3\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__8662\,
            I => \c0.rx.r_SM_Main_dup_3\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__8657\,
            I => \c0.rx.r_SM_Main_dup_3\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__8650\,
            I => \N__8641\
        );

    \I__918\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8636\
        );

    \I__917\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8636\
        );

    \I__916\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8627\
        );

    \I__915\ : InMux
    port map (
            O => \N__8646\,
            I => \N__8627\
        );

    \I__914\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8620\
        );

    \I__913\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8620\
        );

    \I__912\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8617\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8614\
        );

    \I__910\ : InMux
    port map (
            O => \N__8635\,
            I => \N__8607\
        );

    \I__909\ : InMux
    port map (
            O => \N__8634\,
            I => \N__8607\
        );

    \I__908\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8607\
        );

    \I__907\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8604\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8601\
        );

    \I__905\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8596\
        );

    \I__904\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8596\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__8620\,
            I => \c0.rx.N_98_dup\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__8617\,
            I => \c0.rx.N_98_dup\
        );

    \I__901\ : Odrv12
    port map (
            O => \N__8614\,
            I => \c0.rx.N_98_dup\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8607\,
            I => \c0.rx.N_98_dup\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__8604\,
            I => \c0.rx.N_98_dup\
        );

    \I__898\ : Odrv4
    port map (
            O => \N__8601\,
            I => \c0.rx.N_98_dup\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8596\,
            I => \c0.rx.N_98_dup\
        );

    \I__896\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8576\
        );

    \I__895\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8571\
        );

    \I__894\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8571\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8576\,
            I => \N__8561\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__8571\,
            I => \N__8561\
        );

    \I__891\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8556\
        );

    \I__890\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8556\
        );

    \I__889\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8553\
        );

    \I__888\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8548\
        );

    \I__887\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8548\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__8561\,
            I => \N__8545\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8542\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__8553\,
            I => \c0.rx.r_SM_Main_dup_4\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__8548\,
            I => \c0.rx.r_SM_Main_dup_4\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__8545\,
            I => \c0.rx.r_SM_Main_dup_4\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__8542\,
            I => \c0.rx.r_SM_Main_dup_4\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__8533\,
            I => \c0.rx.N_138r_0_i_1_cascade_\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__8530\,
            I => \N__8527\
        );

    \I__878\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8521\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__8526\,
            I => \N__8516\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__8525\,
            I => \N__8513\
        );

    \I__875\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8509\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8506\
        );

    \I__873\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8501\
        );

    \I__872\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8501\
        );

    \I__871\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8494\
        );

    \I__870\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8494\
        );

    \I__869\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8494\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__8509\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__8506\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__8501\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__8494\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__8485\,
            I => \c0.rx.N_91_0_cascade_\
        );

    \I__863\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8479\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__8479\,
            I => \c0.rx.r_SM_Main_illegal_0\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__8476\,
            I => \c0.rx.r_SM_Main_ns_0_i_a2_0_3_cascade_\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__8473\,
            I => \c0.rx.N_320_cascade_\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__8470\,
            I => \c0.rx.r_Clock_Count_8_f0_0_o2_0_2_cascade_\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__8467\,
            I => \N__8463\
        );

    \I__857\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8460\
        );

    \I__856\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8457\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__8460\,
            I => \c0.rx.un1_r_Clock_Count_2_sqmuxa_0_i\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__8457\,
            I => \c0.rx.un1_r_Clock_Count_2_sqmuxa_0_i\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__8452\,
            I => \N__8449\
        );

    \I__852\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8446\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__8446\,
            I => \c0.rx.r_Clock_Count_8_f0_0_o2_0_2\
        );

    \I__850\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8440\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__8440\,
            I => \c0.rx.r_Clock_Count_RNO_0_0_2\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__8437\,
            I => \c0.rx.N_332_cascade_\
        );

    \I__847\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8430\
        );

    \I__846\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8427\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8430\,
            I => \c0.rx.r_Clock_CountZ1Z_2\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__8427\,
            I => \c0.rx.r_Clock_CountZ1Z_2\
        );

    \I__843\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8418\
        );

    \I__842\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8415\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8418\,
            I => \c0.rx.r_Clock_CountZ1Z_6\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__8415\,
            I => \c0.rx.r_Clock_CountZ1Z_6\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__8410\,
            I => \N__8406\
        );

    \I__838\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8403\
        );

    \I__837\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8400\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8403\,
            I => \c0.rx.r_Clock_CountZ0Z_7\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__8400\,
            I => \c0.rx.r_Clock_CountZ0Z_7\
        );

    \I__834\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8391\
        );

    \I__833\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8388\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8391\,
            I => \c0.rx.r_Clock_CountZ1Z_4\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8388\,
            I => \c0.rx.r_Clock_CountZ1Z_4\
        );

    \I__830\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8380\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8380\,
            I => \c0.rx.r_Clock_Count_RNO_0Z0Z_5\
        );

    \I__828\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8373\
        );

    \I__827\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8370\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__8373\,
            I => \c0.rx.r_Clock_CountZ1Z_5\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__8370\,
            I => \c0.rx.r_Clock_CountZ1Z_5\
        );

    \I__824\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8361\
        );

    \I__823\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8358\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__8361\,
            I => \c0.rx.N_320\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__8358\,
            I => \c0.rx.N_320\
        );

    \I__820\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8348\
        );

    \I__819\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8343\
        );

    \I__818\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8343\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__8348\,
            I => \c0.rx.N_317\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__8343\,
            I => \c0.rx.N_317\
        );

    \I__815\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8335\,
            I => \c0.rx.N_337\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__8332\,
            I => \c0.rx.N_383_cascade_\
        );

    \I__812\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8326\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8326\,
            I => \c0.rx.r_Clock_Count_RNO_0_0_1\
        );

    \I__810\ : InMux
    port map (
            O => \N__8323\,
            I => \c0.rx.un1_r_Clock_Count_5_cry_0\
        );

    \I__809\ : InMux
    port map (
            O => \N__8320\,
            I => \c0.rx.un1_r_Clock_Count_5_cry_1\
        );

    \I__808\ : InMux
    port map (
            O => \N__8317\,
            I => \c0.rx.un1_r_Clock_Count_5_cry_2\
        );

    \I__807\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8311\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8311\,
            I => \c0.rx.r_Clock_Count_RNO_0Z0Z_4\
        );

    \I__805\ : InMux
    port map (
            O => \N__8308\,
            I => \c0.rx.un1_r_Clock_Count_5_cry_3\
        );

    \I__804\ : InMux
    port map (
            O => \N__8305\,
            I => \c0.rx.un1_r_Clock_Count_5_cry_4\
        );

    \I__803\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8299\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__8299\,
            I => \c0.rx.r_Clock_Count_RNO_0Z0Z_6\
        );

    \I__801\ : InMux
    port map (
            O => \N__8296\,
            I => \c0.rx.un1_r_Clock_Count_5_cry_5\
        );

    \I__800\ : InMux
    port map (
            O => \N__8293\,
            I => \c0.rx.un1_r_Clock_Count_5_cry_6\
        );

    \I__799\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__8287\,
            I => \c0.rx.r_Clock_Count_RNO_0Z0Z_7\
        );

    \I__797\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8280\
        );

    \I__796\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8277\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8280\,
            I => \c0.rx.r_Clock_CountZ1Z_1\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__8277\,
            I => \c0.rx.r_Clock_CountZ1Z_1\
        );

    \I__793\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8268\
        );

    \I__792\ : InMux
    port map (
            O => \N__8271\,
            I => \N__8265\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8268\,
            I => \c0.rx.r_Clock_CountZ1Z_0\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__8265\,
            I => \c0.rx.r_Clock_CountZ1Z_0\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__8260\,
            I => \c0.rx.r_Rx_Bytece_0_5_cascade_\
        );

    \I__788\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8252\
        );

    \I__787\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8249\
        );

    \I__786\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8246\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8252\,
            I => \c0.rx.N_388\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__8249\,
            I => \c0.rx.N_388\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__8246\,
            I => \c0.rx.N_388\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__8239\,
            I => \c0.rx.r_Rx_Bytece_0_6_cascade_\
        );

    \I__781\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8227\
        );

    \I__780\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8224\
        );

    \I__779\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8221\
        );

    \I__778\ : InMux
    port map (
            O => \N__8233\,
            I => \N__8216\
        );

    \I__777\ : InMux
    port map (
            O => \N__8232\,
            I => \N__8216\
        );

    \I__776\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8211\
        );

    \I__775\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8211\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8227\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8224\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8221\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__8216\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__8211\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__769\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__8197\,
            I => \c0.rx.r_Rx_Bytece_0_0\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__8194\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa_cascade_\
        );

    \I__766\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8188\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__8188\,
            I => \c0.rx.r_Clock_Count_RNO_0_0_0\
        );

    \I__764\ : InMux
    port map (
            O => \N__8185\,
            I => blink_counter_cry_20
        );

    \I__763\ : InMux
    port map (
            O => \N__8182\,
            I => blink_counter_cry_21
        );

    \I__762\ : InMux
    port map (
            O => \N__8179\,
            I => blink_counter_cry_22
        );

    \I__761\ : InMux
    port map (
            O => \N__8176\,
            I => \bfn_6_24_0_\
        );

    \I__760\ : InMux
    port map (
            O => \N__8173\,
            I => blink_counter_cry_24
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__8170\,
            I => \c0.rx.r_Rx_Bytece_0_2_cascade_\
        );

    \I__758\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__8164\,
            I => \c0.rx.N_325\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__8161\,
            I => \c0.rx.N_325_cascade_\
        );

    \I__755\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8155\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__8155\,
            I => \blink_counterZ0Z_13\
        );

    \I__753\ : InMux
    port map (
            O => \N__8152\,
            I => blink_counter_cry_12
        );

    \I__752\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8146\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8146\,
            I => \blink_counterZ0Z_14\
        );

    \I__750\ : InMux
    port map (
            O => \N__8143\,
            I => blink_counter_cry_13
        );

    \I__749\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8137\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__8137\,
            I => \blink_counterZ0Z_15\
        );

    \I__747\ : InMux
    port map (
            O => \N__8134\,
            I => blink_counter_cry_14
        );

    \I__746\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8128\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8128\,
            I => \blink_counterZ0Z_16\
        );

    \I__744\ : InMux
    port map (
            O => \N__8125\,
            I => \bfn_6_23_0_\
        );

    \I__743\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8119\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__8119\,
            I => \blink_counterZ0Z_17\
        );

    \I__741\ : InMux
    port map (
            O => \N__8116\,
            I => blink_counter_cry_16
        );

    \I__740\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8110\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__8110\,
            I => \blink_counterZ0Z_18\
        );

    \I__738\ : InMux
    port map (
            O => \N__8107\,
            I => blink_counter_cry_17
        );

    \I__737\ : InMux
    port map (
            O => \N__8104\,
            I => \N__8101\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__8101\,
            I => \blink_counterZ0Z_19\
        );

    \I__735\ : InMux
    port map (
            O => \N__8098\,
            I => blink_counter_cry_18
        );

    \I__734\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8092\,
            I => \blink_counterZ0Z_20\
        );

    \I__732\ : InMux
    port map (
            O => \N__8089\,
            I => blink_counter_cry_19
        );

    \I__731\ : InMux
    port map (
            O => \N__8086\,
            I => \N__8083\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__8083\,
            I => \blink_counterZ0Z_4\
        );

    \I__729\ : InMux
    port map (
            O => \N__8080\,
            I => blink_counter_cry_3
        );

    \I__728\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8074\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__8074\,
            I => \blink_counterZ0Z_5\
        );

    \I__726\ : InMux
    port map (
            O => \N__8071\,
            I => blink_counter_cry_4
        );

    \I__725\ : InMux
    port map (
            O => \N__8068\,
            I => \N__8065\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__8065\,
            I => \blink_counterZ0Z_6\
        );

    \I__723\ : InMux
    port map (
            O => \N__8062\,
            I => blink_counter_cry_5
        );

    \I__722\ : InMux
    port map (
            O => \N__8059\,
            I => \N__8056\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__8056\,
            I => \blink_counterZ0Z_7\
        );

    \I__720\ : InMux
    port map (
            O => \N__8053\,
            I => blink_counter_cry_6
        );

    \I__719\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8047\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__8047\,
            I => \blink_counterZ0Z_8\
        );

    \I__717\ : InMux
    port map (
            O => \N__8044\,
            I => \bfn_6_22_0_\
        );

    \I__716\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8038\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__8038\,
            I => \blink_counterZ0Z_9\
        );

    \I__714\ : InMux
    port map (
            O => \N__8035\,
            I => blink_counter_cry_8
        );

    \I__713\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8029\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__8029\,
            I => \blink_counterZ0Z_10\
        );

    \I__711\ : InMux
    port map (
            O => \N__8026\,
            I => blink_counter_cry_9
        );

    \I__710\ : InMux
    port map (
            O => \N__8023\,
            I => \N__8020\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__8020\,
            I => \blink_counterZ0Z_11\
        );

    \I__708\ : InMux
    port map (
            O => \N__8017\,
            I => blink_counter_cry_10
        );

    \I__707\ : InMux
    port map (
            O => \N__8014\,
            I => \N__8011\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__8011\,
            I => \blink_counterZ0Z_12\
        );

    \I__705\ : InMux
    port map (
            O => \N__8008\,
            I => blink_counter_cry_11
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__8005\,
            I => \c0.rx.r_SM_Main_RNI58REZ0Z_0_cascade_\
        );

    \I__703\ : IoInMux
    port map (
            O => \N__8002\,
            I => \N__7999\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7996\
        );

    \I__701\ : Span4Mux_s1_h
    port map (
            O => \N__7996\,
            I => \N__7993\
        );

    \I__700\ : Span4Mux_h
    port map (
            O => \N__7993\,
            I => \N__7990\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__7990\,
            I => \c0.rx.rx_data_ready\
        );

    \I__698\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7984\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__7984\,
            I => \blink_counterZ0Z_0\
        );

    \I__696\ : InMux
    port map (
            O => \N__7981\,
            I => \bfn_6_21_0_\
        );

    \I__695\ : InMux
    port map (
            O => \N__7978\,
            I => \N__7975\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__7975\,
            I => \blink_counterZ0Z_1\
        );

    \I__693\ : InMux
    port map (
            O => \N__7972\,
            I => blink_counter_cry_0
        );

    \I__692\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7966\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__7966\,
            I => \blink_counterZ0Z_2\
        );

    \I__690\ : InMux
    port map (
            O => \N__7963\,
            I => blink_counter_cry_1
        );

    \I__689\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7957\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__7957\,
            I => \blink_counterZ0Z_3\
        );

    \I__687\ : InMux
    port map (
            O => \N__7954\,
            I => blink_counter_cry_2
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__7951\,
            I => \c0.rx.N_336_cascade_\
        );

    \I__685\ : InMux
    port map (
            O => \N__7948\,
            I => \N__7945\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__7945\,
            I => \c0.rx.r_Rx_Bytece_0_1\
        );

    \I__683\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7938\
        );

    \I__682\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7938\,
            I => \c0.tx.r_Clock_Count_i_0\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__7935\,
            I => \c0.tx.r_Clock_Count_i_0\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__7930\,
            I => \c0.rx.r_Rx_Bytece_0_4_cascade_\
        );

    \I__678\ : InMux
    port map (
            O => \N__7927\,
            I => \N__7924\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__7924\,
            I => \N__7921\
        );

    \I__676\ : Span4Mux_v
    port map (
            O => \N__7921\,
            I => \N__7918\
        );

    \I__675\ : Span4Mux_v
    port map (
            O => \N__7918\,
            I => \N__7915\
        );

    \I__674\ : Span4Mux_v
    port map (
            O => \N__7915\,
            I => \N__7912\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__7912\,
            I => \PIN_2_c\
        );

    \I__672\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__7906\,
            I => \N__7903\
        );

    \I__670\ : Span4Mux_h
    port map (
            O => \N__7903\,
            I => \N__7900\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__7900\,
            I => \c0.rx.r_Rx_Data_RZ0\
        );

    \I__668\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7894\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__7894\,
            I => \c0.tx.r_Clock_Count_i_1\
        );

    \I__666\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7888\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__7888\,
            I => \c0.tx.r_Clock_Count_i_2\
        );

    \I__664\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7882\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__7882\,
            I => \c0.tx.r_Clock_Count_i_3\
        );

    \I__662\ : InMux
    port map (
            O => \N__7879\,
            I => \c0.tx.r_Clock_Count12\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_5_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_22_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.i12\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.data_cry_7\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_6_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => blink_counter_cry_7,
            carryinitout => \bfn_6_22_0_\
        );

    \IN_MUX_bfv_6_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => blink_counter_cry_15,
            carryinitout => \bfn_6_23_0_\
        );

    \IN_MUX_bfv_6_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => blink_counter_cry_23,
            carryinitout => \bfn_6_24_0_\
        );

    \c0.rx.r_Rx_DV_RNID002\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8002\,
            GLOBALBUFFEROUTPUT => \c0.rx_data_ready_g\
        );

    \c0.byte_transmit_counter_RNI4QES5_0_2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__15046\,
            GLOBALBUFFEROUTPUT => \c0.data_out_0__1_sqmuxa_g\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19270\,
            GLOBALBUFFEROUTPUT => \c0.data_in_frame_0__0_sqmuxa_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_R_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7927\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.r_Rx_Data_RZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7909\,
            lcout => \c0.rx.r_Rx_DataZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_0_c_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7941\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_22_0_\,
            carryout => \c0.tx.r_Clock_Count12_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9464\,
            in1 => \N__7897\,
            in2 => \N__17115\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx.r_Clock_Count_i_1\,
            ltout => OPEN,
            carryin => \c0.tx.r_Clock_Count12_cry_0\,
            carryout => \c0.tx.r_Clock_Count12_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7891\,
            in2 => \N__17092\,
            in3 => \N__9485\,
            lcout => \c0.tx.r_Clock_Count_i_2\,
            ltout => OPEN,
            carryin => \c0.tx.r_Clock_Count12_cry_1\,
            carryout => \c0.tx.r_Clock_Count12_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7885\,
            in2 => \N__17116\,
            in3 => \N__9438\,
            lcout => \c0.tx.r_Clock_Count_i_3\,
            ltout => OPEN,
            carryin => \c0.tx.r_Clock_Count12_cry_2\,
            carryout => \c0.tx.r_Clock_Count12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7879\,
            lcout => \c0.tx.r_Clock_Count12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__0_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17104\,
            lcout => \c0.d_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19587\,
            ce => 'H',
            sr => \N__16882\
        );

    \c0.data_out_3__3_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19587\,
            ce => 'H',
            sr => \N__16882\
        );

    \c0.tx.r_SM_Main_RNO_0_1_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__9958\,
            in1 => \N__9876\,
            in2 => \_gnd_net_\,
            in3 => \N__10539\,
            lcout => \c0.tx.r_SM_Main_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_0_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__9877\,
            in1 => \N__9334\,
            in2 => \N__10368\,
            in3 => \N__9768\,
            lcout => \c0.tx.r_Clock_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__17056\,
            in1 => \N__9420\,
            in2 => \_gnd_net_\,
            in3 => \N__7942\,
            lcout => \c0.tx.r_Clock_Count_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_1_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__9878\,
            in1 => \N__9322\,
            in2 => \N__10369\,
            in3 => \N__9769\,
            lcout => \c0.tx.r_Clock_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_2_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__9766\,
            in1 => \N__10360\,
            in2 => \N__9883\,
            in3 => \N__9517\,
            lcout => \c0.tx.r_Clock_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_3_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__9879\,
            in1 => \N__9767\,
            in2 => \N__10367\,
            in3 => \N__9502\,
            lcout => \c0.tx.r_Clock_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_4_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14233\,
            in1 => \N__14112\,
            in2 => \_gnd_net_\,
            in3 => \N__14178\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_Bytece_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_4_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__9046\,
            in1 => \N__12228\,
            in2 => \N__7930\,
            in3 => \N__8235\,
            lcout => \c0.rx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_1_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__14117\,
            in1 => \N__8256\,
            in2 => \N__14246\,
            in3 => \N__8849\,
            lcout => \c0.rx.r_Bit_IndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_0_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__14116\,
            in1 => \N__8255\,
            in2 => \_gnd_net_\,
            in3 => \N__8848\,
            lcout => \c0.rx.r_Bit_IndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_3_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14173\,
            in2 => \_gnd_net_\,
            in3 => \N__8167\,
            lcout => OPEN,
            ltout => \c0.rx.N_336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_3_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__10218\,
            in1 => \N__9048\,
            in2 => \N__7951\,
            in3 => \N__8236\,
            lcout => \c0.rx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_1_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14227\,
            in1 => \N__14174\,
            in2 => \_gnd_net_\,
            in3 => \N__14109\,
            lcout => \c0.rx.r_Rx_Bytece_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_6_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8886\,
            in1 => \N__8832\,
            in2 => \N__8788\,
            in3 => \N__8302\,
            lcout => \c0.rx.r_Clock_CountZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_1_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__8830\,
            in1 => \N__8884\,
            in2 => \N__8919\,
            in3 => \N__8329\,
            lcout => \c0.rx.r_Clock_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_1_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__7948\,
            in1 => \N__9044\,
            in2 => \N__10203\,
            in3 => \N__8234\,
            lcout => \c0.rx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_4_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8885\,
            in1 => \N__8831\,
            in2 => \N__8787\,
            in3 => \N__8314\,
            lcout => \c0.rx.r_Clock_CountZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_0_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__8883\,
            in1 => \N__8829\,
            in2 => \N__8920\,
            in3 => \N__8191\,
            lcout => \c0.rx.r_Clock_CountZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNO_0_1_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__8520\,
            in1 => \N__9045\,
            in2 => \_gnd_net_\,
            in3 => \N__9145\,
            lcout => \c0.rx.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNI58RE_0_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8632\,
            in2 => \_gnd_net_\,
            in3 => \N__8519\,
            lcout => \c0.rx.r_SM_Main_RNI58REZ0Z_0\,
            ltout => \c0.rx.r_SM_Main_RNI58REZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_7_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8779\,
            in1 => \N__8882\,
            in2 => \N__8005\,
            in3 => \N__8290\,
            lcout => \c0.rx.r_Clock_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010100010"
        )
    port map (
            in0 => \N__8847\,
            in1 => \N__9115\,
            in2 => \N__17734\,
            in3 => \N__8581\,
            lcout => \c0.rx.rx_data_ready\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_0_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7987\,
            in2 => \_gnd_net_\,
            in3 => \N__7981\,
            lcout => \blink_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => blink_counter_cry_0,
            clk => \N__19588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7978\,
            in2 => \_gnd_net_\,
            in3 => \N__7972\,
            lcout => \blink_counterZ0Z_1\,
            ltout => OPEN,
            carryin => blink_counter_cry_0,
            carryout => blink_counter_cry_1,
            clk => \N__19588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7969\,
            in2 => \_gnd_net_\,
            in3 => \N__7963\,
            lcout => \blink_counterZ0Z_2\,
            ltout => OPEN,
            carryin => blink_counter_cry_1,
            carryout => blink_counter_cry_2,
            clk => \N__19588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_3_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7960\,
            in2 => \_gnd_net_\,
            in3 => \N__7954\,
            lcout => \blink_counterZ0Z_3\,
            ltout => OPEN,
            carryin => blink_counter_cry_2,
            carryout => blink_counter_cry_3,
            clk => \N__19588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_4_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8086\,
            in2 => \_gnd_net_\,
            in3 => \N__8080\,
            lcout => \blink_counterZ0Z_4\,
            ltout => OPEN,
            carryin => blink_counter_cry_3,
            carryout => blink_counter_cry_4,
            clk => \N__19588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_5_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8077\,
            in2 => \_gnd_net_\,
            in3 => \N__8071\,
            lcout => \blink_counterZ0Z_5\,
            ltout => OPEN,
            carryin => blink_counter_cry_4,
            carryout => blink_counter_cry_5,
            clk => \N__19588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_6_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8068\,
            in2 => \_gnd_net_\,
            in3 => \N__8062\,
            lcout => \blink_counterZ0Z_6\,
            ltout => OPEN,
            carryin => blink_counter_cry_5,
            carryout => blink_counter_cry_6,
            clk => \N__19588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_7_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8059\,
            in2 => \_gnd_net_\,
            in3 => \N__8053\,
            lcout => \blink_counterZ0Z_7\,
            ltout => OPEN,
            carryin => blink_counter_cry_6,
            carryout => blink_counter_cry_7,
            clk => \N__19588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_8_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8050\,
            in2 => \_gnd_net_\,
            in3 => \N__8044\,
            lcout => \blink_counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_6_22_0_\,
            carryout => blink_counter_cry_8,
            clk => \N__19595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_9_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8041\,
            in2 => \_gnd_net_\,
            in3 => \N__8035\,
            lcout => \blink_counterZ0Z_9\,
            ltout => OPEN,
            carryin => blink_counter_cry_8,
            carryout => blink_counter_cry_9,
            clk => \N__19595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_10_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8032\,
            in2 => \_gnd_net_\,
            in3 => \N__8026\,
            lcout => \blink_counterZ0Z_10\,
            ltout => OPEN,
            carryin => blink_counter_cry_9,
            carryout => blink_counter_cry_10,
            clk => \N__19595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_11_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8023\,
            in2 => \_gnd_net_\,
            in3 => \N__8017\,
            lcout => \blink_counterZ0Z_11\,
            ltout => OPEN,
            carryin => blink_counter_cry_10,
            carryout => blink_counter_cry_11,
            clk => \N__19595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_12_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8014\,
            in2 => \_gnd_net_\,
            in3 => \N__8008\,
            lcout => \blink_counterZ0Z_12\,
            ltout => OPEN,
            carryin => blink_counter_cry_11,
            carryout => blink_counter_cry_12,
            clk => \N__19595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_13_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8158\,
            in2 => \_gnd_net_\,
            in3 => \N__8152\,
            lcout => \blink_counterZ0Z_13\,
            ltout => OPEN,
            carryin => blink_counter_cry_12,
            carryout => blink_counter_cry_13,
            clk => \N__19595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_14_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8149\,
            in2 => \_gnd_net_\,
            in3 => \N__8143\,
            lcout => \blink_counterZ0Z_14\,
            ltout => OPEN,
            carryin => blink_counter_cry_13,
            carryout => blink_counter_cry_14,
            clk => \N__19595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_15_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8140\,
            in2 => \_gnd_net_\,
            in3 => \N__8134\,
            lcout => \blink_counterZ0Z_15\,
            ltout => OPEN,
            carryin => blink_counter_cry_14,
            carryout => blink_counter_cry_15,
            clk => \N__19595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_16_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8131\,
            in2 => \_gnd_net_\,
            in3 => \N__8125\,
            lcout => \blink_counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_6_23_0_\,
            carryout => blink_counter_cry_16,
            clk => \N__19600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_17_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8122\,
            in2 => \_gnd_net_\,
            in3 => \N__8116\,
            lcout => \blink_counterZ0Z_17\,
            ltout => OPEN,
            carryin => blink_counter_cry_16,
            carryout => blink_counter_cry_17,
            clk => \N__19600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_18_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8113\,
            in2 => \_gnd_net_\,
            in3 => \N__8107\,
            lcout => \blink_counterZ0Z_18\,
            ltout => OPEN,
            carryin => blink_counter_cry_17,
            carryout => blink_counter_cry_18,
            clk => \N__19600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_19_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8104\,
            in2 => \_gnd_net_\,
            in3 => \N__8098\,
            lcout => \blink_counterZ0Z_19\,
            ltout => OPEN,
            carryin => blink_counter_cry_18,
            carryout => blink_counter_cry_19,
            clk => \N__19600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_20_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8095\,
            in2 => \_gnd_net_\,
            in3 => \N__8089\,
            lcout => \blink_counterZ0Z_20\,
            ltout => OPEN,
            carryin => blink_counter_cry_19,
            carryout => blink_counter_cry_20,
            clk => \N__19600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_21_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9294\,
            in2 => \_gnd_net_\,
            in3 => \N__8185\,
            lcout => \blink_counterZ0Z_21\,
            ltout => OPEN,
            carryin => blink_counter_cry_20,
            carryout => blink_counter_cry_21,
            clk => \N__19600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_22_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9273\,
            in2 => \_gnd_net_\,
            in3 => \N__8182\,
            lcout => \blink_counterZ0Z_22\,
            ltout => OPEN,
            carryin => blink_counter_cry_21,
            carryout => blink_counter_cry_22,
            clk => \N__19600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_23_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9201\,
            in2 => \_gnd_net_\,
            in3 => \N__8179\,
            lcout => \blink_counterZ0Z_23\,
            ltout => OPEN,
            carryin => blink_counter_cry_22,
            carryout => blink_counter_cry_23,
            clk => \N__19600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_24_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9249\,
            in2 => \_gnd_net_\,
            in3 => \N__8176\,
            lcout => \blink_counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_6_24_0_\,
            carryout => blink_counter_cry_24,
            clk => \N__19607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_25_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9222\,
            in2 => \_gnd_net_\,
            in3 => \N__8173\,
            lcout => \blink_counterZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_2_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__14104\,
            in1 => \_gnd_net_\,
            in2 => \N__14237\,
            in3 => \N__14176\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_Bytece_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__12210\,
            in1 => \N__9047\,
            in2 => \N__8170\,
            in3 => \N__8232\,
            lcout => \c0.rx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_RNIHTCD_1_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14217\,
            in2 => \_gnd_net_\,
            in3 => \N__14103\,
            lcout => \c0.rx.N_325\,
            ltout => \c0.rx.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_2_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010011000000000"
        )
    port map (
            in0 => \N__14180\,
            in1 => \N__8257\,
            in2 => \N__8161\,
            in3 => \N__8850\,
            lcout => \c0.rx.r_Bit_IndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_5_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14177\,
            in1 => \N__14221\,
            in2 => \_gnd_net_\,
            in3 => \N__14105\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_Bytece_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_5_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__8233\,
            in1 => \N__15717\,
            in2 => \N__8260\,
            in3 => \N__9049\,
            lcout => \c0.rx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNI91B33_0_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__8710\,
            in1 => \N__8649\,
            in2 => \N__8530\,
            in3 => \N__9103\,
            lcout => \c0.rx.N_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_0_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14244\,
            in1 => \N__14110\,
            in2 => \_gnd_net_\,
            in3 => \N__14175\,
            lcout => \c0.rx.r_Rx_Bytece_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_7_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__9052\,
            in1 => \N__14056\,
            in2 => \N__10866\,
            in3 => \N__8231\,
            lcout => \c0.rx_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_6_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14111\,
            in1 => \N__14245\,
            in2 => \_gnd_net_\,
            in3 => \N__14179\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_Bytece_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_6_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__16068\,
            in1 => \N__9051\,
            in2 => \N__8239\,
            in3 => \N__8230\,
            lcout => \c0.rx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNIJ0FM2_2_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8709\,
            in1 => \N__9102\,
            in2 => \_gnd_net_\,
            in3 => \N__8648\,
            lcout => \c0.rx.r_Rx_Byte_1_sqmuxa\,
            ltout => \c0.rx.r_Rx_Byte_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_0_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__10413\,
            in1 => \N__8200\,
            in2 => \N__8194\,
            in3 => \N__9050\,
            lcout => \c0.rx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8272\,
            in2 => \N__8467\,
            in3 => \N__8466\,
            lcout => \c0.rx.r_Clock_Count_RNO_0_0_0\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \c0.rx.un1_r_Clock_Count_5_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_1_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8284\,
            in2 => \_gnd_net_\,
            in3 => \N__8323\,
            lcout => \c0.rx.r_Clock_Count_RNO_0_0_1\,
            ltout => OPEN,
            carryin => \c0.rx.un1_r_Clock_Count_5_cry_0\,
            carryout => \c0.rx.un1_r_Clock_Count_5_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_2_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8434\,
            in2 => \_gnd_net_\,
            in3 => \N__8320\,
            lcout => \c0.rx.r_Clock_Count_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \c0.rx.un1_r_Clock_Count_5_cry_1\,
            carryout => \c0.rx.un1_r_Clock_Count_5_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_3_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8737\,
            in2 => \_gnd_net_\,
            in3 => \N__8317\,
            lcout => \c0.rx.r_Clock_Count_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \c0.rx.un1_r_Clock_Count_5_cry_2\,
            carryout => \c0.rx.un1_r_Clock_Count_5_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_4_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8395\,
            in2 => \_gnd_net_\,
            in3 => \N__8308\,
            lcout => \c0.rx.r_Clock_Count_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \c0.rx.un1_r_Clock_Count_5_cry_3\,
            carryout => \c0.rx.un1_r_Clock_Count_5_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_5_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8377\,
            in2 => \_gnd_net_\,
            in3 => \N__8305\,
            lcout => \c0.rx.r_Clock_Count_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \c0.rx.un1_r_Clock_Count_5_cry_4\,
            carryout => \c0.rx.un1_r_Clock_Count_5_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_6_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8422\,
            in2 => \_gnd_net_\,
            in3 => \N__8296\,
            lcout => \c0.rx.r_Clock_Count_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \c0.rx.un1_r_Clock_Count_5_cry_5\,
            carryout => \c0.rx.un1_r_Clock_Count_5_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_7_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8409\,
            in2 => \_gnd_net_\,
            in3 => \N__8293\,
            lcout => \c0.rx.r_Clock_Count_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNIL4RQ_0_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__8433\,
            in1 => \N__8283\,
            in2 => \_gnd_net_\,
            in3 => \N__8271\,
            lcout => \c0.rx.N_320\,
            ltout => \c0.rx.N_320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNITSB13_3_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110110"
        )
    port map (
            in0 => \N__8734\,
            in1 => \N__8943\,
            in2 => \N__8473\,
            in3 => \N__8351\,
            lcout => \c0.rx.r_Clock_Count_8_f0_0_o2_0_2\,
            ltout => \c0.rx.r_Clock_Count_8_f0_0_o2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNINFV94_0_4_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__8944\,
            in1 => \N__8579\,
            in2 => \N__8470\,
            in3 => \N__8625\,
            lcout => \c0.rx.un1_r_Clock_Count_2_sqmuxa_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNICMJ72_3_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__8735\,
            in1 => \N__8364\,
            in2 => \_gnd_net_\,
            in3 => \N__8352\,
            lcout => \c0.rx.N_386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNINFV94_4_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__8945\,
            in1 => \N__8580\,
            in2 => \N__8452\,
            in3 => \N__8626\,
            lcout => \c0.rx.N_332\,
            ltout => \c0.rx.N_332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_2_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__8443\,
            in1 => \N__8912\,
            in2 => \N__8437\,
            in3 => \N__8833\,
            lcout => \c0.rx.r_Clock_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8421\,
            in1 => \N__8376\,
            in2 => \N__8410\,
            in3 => \N__8394\,
            lcout => \c0.rx.N_317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_5_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8383\,
            in1 => \N__8881\,
            in2 => \N__8786\,
            in3 => \N__8834\,
            lcout => \c0.rx.r_Clock_CountZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNICMJ72_0_3_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8365\,
            in1 => \N__8736\,
            in2 => \_gnd_net_\,
            in3 => \N__8353\,
            lcout => \c0.rx.N_383\,
            ltout => \c0.rx.N_383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_1_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__8644\,
            in1 => \N__8338\,
            in2 => \N__8332\,
            in3 => \N__8524\,
            lcout => \c0.rx.r_SM_Main_dup_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.N_98_ip_RNO_1_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__9140\,
            in1 => \N__8512\,
            in2 => \_gnd_net_\,
            in3 => \N__9093\,
            lcout => \c0.rx.r_SM_Main_illegal_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNO_0_0_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001111"
        )
    port map (
            in0 => \N__8969\,
            in1 => \_gnd_net_\,
            in2 => \N__8526\,
            in3 => \N__9142\,
            lcout => OPEN,
            ltout => \c0.rx.N_138r_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_0_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__9061\,
            in1 => \N__8570\,
            in2 => \N__8533\,
            in3 => \N__8645\,
            lcout => \c0.rx.r_SM_MainZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.N_98_ip_RNO_0_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__9091\,
            in1 => \_gnd_net_\,
            in2 => \N__8525\,
            in3 => \N__9141\,
            lcout => OPEN,
            ltout => \c0.rx.N_91_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.N_98_ip_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111111"
        )
    port map (
            in0 => \N__8673\,
            in1 => \N__8569\,
            in2 => \N__8485\,
            in3 => \N__8482\,
            lcout => \c0.rx.N_98_dup\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNIH6OP_3_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9092\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8672\,
            lcout => \c0.rx.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__9067\,
            in1 => \N__8970\,
            in2 => \N__9154\,
            in3 => \N__8634\,
            lcout => \c0.rx.r_SM_Main_dup_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNO_0_3_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14184\,
            in1 => \N__14125\,
            in2 => \N__14251\,
            in3 => \N__9096\,
            lcout => OPEN,
            ltout => \c0.rx.r_SM_Main_ns_0_i_a2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_3_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__8676\,
            in1 => \N__8707\,
            in2 => \N__8476\,
            in3 => \N__8635\,
            lcout => \c0.rx.r_SM_Main_dup_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNO_1_2_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__9144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9060\,
            lcout => \c0.rx.r_SM_Main_ns_0_i_a2_1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNIHKFL1_1_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8946\,
            in1 => \N__9143\,
            in2 => \N__8650\,
            in3 => \N__8567\,
            lcout => \c0.rx.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_RNO_1_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__8566\,
            in1 => \N__8674\,
            in2 => \_gnd_net_\,
            in3 => \N__9094\,
            lcout => OPEN,
            ltout => \c0.rx.un1_r_Rx_DV7_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_RNO_0_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__8675\,
            in1 => \N__8705\,
            in2 => \N__9118\,
            in3 => \N__8633\,
            lcout => \c0.rx.r_Rx_DV_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNO_0_2_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__8706\,
            in1 => \N__14049\,
            in2 => \_gnd_net_\,
            in3 => \N__9095\,
            lcout => \c0.rx.r_SM_Main_ns_0_i_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNI7GPF_4_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9053\,
            in2 => \_gnd_net_\,
            in3 => \N__8568\,
            lcout => OPEN,
            ltout => \c0.rx.r_Clock_Count_8_f0_0_a2_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.N_98_ip_RNIJK4J3_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8971\,
            in1 => \N__8950\,
            in2 => \N__8923\,
            in3 => \N__8646\,
            lcout => \c0.rx.N_371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_3_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8890\,
            in1 => \N__8854\,
            in2 => \N__8775\,
            in3 => \N__8746\,
            lcout => \c0.rx.r_Clock_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_4_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8708\,
            in1 => \N__8677\,
            in2 => \_gnd_net_\,
            in3 => \N__8647\,
            lcout => \c0.rx.r_SM_Main_dup_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__3_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17075\,
            lcout => \c0.d_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19621\,
            ce => 'H',
            sr => \N__16881\
        );

    \c0.data_out_0__5_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19621\,
            ce => 'H',
            sr => \N__16881\
        );

    \c0.data_out_1__1_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17060\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19631\,
            ce => 'H',
            sr => \N__16880\
        );

    \c0.data_out_7__7_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14875\,
            in1 => \N__14503\,
            in2 => \N__9385\,
            in3 => \N__10090\,
            lcout => \c0.data_out_7_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19590\,
            ce => \N__16838\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNO_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11336\,
            in1 => \N__11048\,
            in2 => \N__13965\,
            in3 => \N__12347\,
            lcout => \c0.i12_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__5_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11170\,
            lcout => \c0.data_in_3_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19591\,
            ce => \N__17716\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__6_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16102\,
            lcout => \c0.data_in_3_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19591\,
            ce => \N__17716\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__6_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11337\,
            lcout => \c0.data_in_2_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19591\,
            ce => \N__17716\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__6_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13613\,
            lcout => \c0.data_in_1_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19591\,
            ce => \N__17716\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_0_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9160\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \c0.i12_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_1_c_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9307\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_0\,
            carryout => \c0.i12_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_2_c_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9676\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_1\,
            carryout => \c0.i12_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_3_c_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9640\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_2\,
            carryout => \c0.i12_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_4_c_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9721\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_3\,
            carryout => \c0.i12_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_5_c_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9688\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_4\,
            carryout => \c0.i12_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_6_c_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9682\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_5\,
            carryout => \c0.i12_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_7_c_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9172\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_6\,
            carryout => \c0.i12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_THRU_LUT4_0_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9163\,
            lcout => \c0.i12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_0_c_RNO_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10254\,
            in1 => \N__12711\,
            in2 => \N__13506\,
            in3 => \N__16113\,
            lcout => \c0.i12_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_1_c_RNO_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15869\,
            in1 => \N__10241\,
            in2 => \N__11127\,
            in3 => \N__10968\,
            lcout => \c0.i12_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_obuf_RNO_1_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001010"
        )
    port map (
            in0 => \N__9301\,
            in1 => \N__9283\,
            in2 => \N__9262\,
            in3 => \N__9231\,
            lcout => \N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_obuf_RNO_0_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__9282\,
            in1 => \N__9258\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \N_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_obuf_RNO_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000101010101"
        )
    port map (
            in0 => \N__9238\,
            in1 => \N__9232\,
            in2 => \N__9211\,
            in3 => \N__9208\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__1_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15870\,
            lcout => \c0.data_in_0_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19609\,
            ce => \N__17723\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__3_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11123\,
            lcout => \c0.data_in_0_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19609\,
            ce => \N__17723\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__4_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_0_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19609\,
            ce => \N__17723\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__6_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13716\,
            lcout => \c0.data_in_0_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19609\,
            ce => \N__17723\,
            sr => \_gnd_net_\
        );

    \c0.tx.N_90_ip_RNO_1_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__10650\,
            in1 => \N__10529\,
            in2 => \_gnd_net_\,
            in3 => \N__9852\,
            lcout => \c0.tx.r_SM_Main_illegal_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.N_90_ip_RNIVJLQ_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__9855\,
            in1 => \N__9940\,
            in2 => \_gnd_net_\,
            in3 => \N__9817\,
            lcout => \c0.tx.N_90_ip_RNIVJLQZ0\,
            ltout => \c0.tx.N_90_ip_RNIVJLQZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.N_90_ip_RNIVJLQ_0_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9370\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx.N_398_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.N_90_ip_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011111111011"
        )
    port map (
            in0 => \N__10316\,
            in1 => \N__9367\,
            in2 => \N__9984\,
            in3 => \N__9358\,
            lcout => \c0.tx.N_90_dup\,
            ltout => \c0.tx.N_90_dup_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNI1GI71_4_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9980\,
            in1 => \N__9854\,
            in2 => \N__9361\,
            in3 => \N__9770\,
            lcout => \c0.tx.r_Clock_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_3_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__10317\,
            in1 => \N__9904\,
            in2 => \N__10618\,
            in3 => \N__9818\,
            lcout => \c0.tx.r_SM_Main_dup_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.N_90_ip_RNO_0_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10651\,
            in1 => \N__10530\,
            in2 => \_gnd_net_\,
            in3 => \N__9853\,
            lcout => \c0.tx.N_83_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_0_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__9979\,
            in1 => \N__9819\,
            in2 => \N__9913\,
            in3 => \N__10652\,
            lcout => \c0.tx.r_SM_MainZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNO_0_0_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9427\,
            in2 => \N__9351\,
            in3 => \N__9352\,
            lcout => \c0.tx.r_Clock_Count_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \c0.tx.un1_r_Clock_Count_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNO_0_1_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9471\,
            in2 => \_gnd_net_\,
            in3 => \N__9310\,
            lcout => \c0.tx.r_Clock_Count_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \c0.tx.un1_r_Clock_Count_cry_0\,
            carryout => \c0.tx.un1_r_Clock_Count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNO_0_2_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9493\,
            in2 => \_gnd_net_\,
            in3 => \N__9508\,
            lcout => \c0.tx.r_Clock_Count_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \c0.tx.un1_r_Clock_Count_cry_1\,
            carryout => \c0.tx.un1_r_Clock_Count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNO_0_3_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9450\,
            in2 => \_gnd_net_\,
            in3 => \N__9505\,
            lcout => \c0.tx.r_Clock_Count_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNI522E_4_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9985\,
            in2 => \_gnd_net_\,
            in3 => \N__9820\,
            lcout => \c0.tx.r_SM_Main_RNI522EZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNI636A_3_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9492\,
            in1 => \N__9472\,
            in2 => \N__9451\,
            in3 => \N__9426\,
            lcout => \c0.tx.N_171_0\,
            ltout => \c0.tx.N_171_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_1_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__9821\,
            in1 => \N__9409\,
            in2 => \N__9397\,
            in3 => \N__9863\,
            lcout => \c0.tx.r_SM_Main_dup_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_0_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__9391\,
            in1 => \N__15529\,
            in2 => \N__10063\,
            in3 => \N__15379\,
            lcout => \c0.tx_data_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_0_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13013\,
            in1 => \N__14470\,
            in2 => \_gnd_net_\,
            in3 => \N__11778\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_0_a2_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__0_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14498\,
            in1 => \N__11517\,
            in2 => \N__9394\,
            in3 => \N__10023\,
            lcout => \c0.data_out_6_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19632\,
            ce => \N__16837\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_7_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__10896\,
            in1 => \N__13329\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__5_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9610\,
            lcout => \c0.d_2_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19638\,
            ce => \N__16836\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__1_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9571\,
            lcout => \c0.d_2_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19638\,
            ce => \N__16836\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__3_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9631\,
            lcout => \c0.d_2_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19638\,
            ce => \N__16836\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__1_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9532\,
            lcout => \c0.d_2_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19646\,
            ce => \N__16834\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__7_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9589\,
            lcout => \c0.d_2_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19646\,
            ce => \N__16834\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__5_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9664\,
            lcout => \c0.d_2_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19646\,
            ce => \N__16834\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__2_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9553\,
            lcout => \c0.d_2_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19646\,
            ce => \N__16834\,
            sr => \_gnd_net_\
        );

    \c0.data_0_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10185\,
            in2 => \_gnd_net_\,
            in3 => \N__9535\,
            lcout => \c0.dataZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \c0.data_cry_0\,
            clk => \N__19652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_1_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9531\,
            in2 => \_gnd_net_\,
            in3 => \N__9520\,
            lcout => \c0.dataZ0Z_1\,
            ltout => OPEN,
            carryin => \c0.data_cry_0\,
            carryout => \c0.data_cry_1\,
            clk => \N__19652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_2_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10149\,
            in2 => \_gnd_net_\,
            in3 => \N__9634\,
            lcout => \c0.dataZ0Z_2\,
            ltout => OPEN,
            carryin => \c0.data_cry_1\,
            carryout => \c0.data_cry_2\,
            clk => \N__19652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_3_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9627\,
            in2 => \_gnd_net_\,
            in3 => \N__9616\,
            lcout => \c0.dataZ0Z_3\,
            ltout => OPEN,
            carryin => \c0.data_cry_2\,
            carryout => \c0.data_cry_3\,
            clk => \N__19652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_4_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10125\,
            in2 => \_gnd_net_\,
            in3 => \N__9613\,
            lcout => \c0.dataZ0Z_4\,
            ltout => OPEN,
            carryin => \c0.data_cry_3\,
            carryout => \c0.data_cry_4\,
            clk => \N__19652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_5_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9606\,
            in2 => \_gnd_net_\,
            in3 => \N__9595\,
            lcout => \c0.dataZ0Z_5\,
            ltout => OPEN,
            carryin => \c0.data_cry_4\,
            carryout => \c0.data_cry_5\,
            clk => \N__19652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_6_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10740\,
            in2 => \_gnd_net_\,
            in3 => \N__9592\,
            lcout => \c0.dataZ0Z_6\,
            ltout => OPEN,
            carryin => \c0.data_cry_5\,
            carryout => \c0.data_cry_6\,
            clk => \N__19652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_7_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9588\,
            in2 => \_gnd_net_\,
            in3 => \N__9577\,
            lcout => \c0.dataZ0Z_7\,
            ltout => OPEN,
            carryin => \c0.data_cry_6\,
            carryout => \c0.data_cry_7\,
            clk => \N__19652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_8_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10113\,
            in2 => \_gnd_net_\,
            in3 => \N__9574\,
            lcout => \c0.dataZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_28_0_\,
            carryout => \c0.data_cry_8\,
            clk => \N__19661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_9_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9567\,
            in2 => \_gnd_net_\,
            in3 => \N__9556\,
            lcout => \c0.dataZ0Z_9\,
            ltout => OPEN,
            carryin => \c0.data_cry_8\,
            carryout => \c0.data_cry_9\,
            clk => \N__19661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_10_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9549\,
            in2 => \_gnd_net_\,
            in3 => \N__9538\,
            lcout => \c0.dataZ0Z_10\,
            ltout => OPEN,
            carryin => \c0.data_cry_9\,
            carryout => \c0.data_cry_10\,
            clk => \N__19661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_11_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10161\,
            in2 => \_gnd_net_\,
            in3 => \N__9670\,
            lcout => \c0.dataZ0Z_11\,
            ltout => OPEN,
            carryin => \c0.data_cry_10\,
            carryout => \c0.data_cry_11\,
            clk => \N__19661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_12_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10038\,
            in2 => \_gnd_net_\,
            in3 => \N__9667\,
            lcout => \c0.dataZ0Z_12\,
            ltout => OPEN,
            carryin => \c0.data_cry_11\,
            carryout => \c0.data_cry_12\,
            clk => \N__19661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_13_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9660\,
            in2 => \_gnd_net_\,
            in3 => \N__9649\,
            lcout => \c0.dataZ0Z_13\,
            ltout => OPEN,
            carryin => \c0.data_cry_12\,
            carryout => \c0.data_cry_13\,
            clk => \N__19661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_14_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10173\,
            in2 => \_gnd_net_\,
            in3 => \N__9646\,
            lcout => \c0.dataZ0Z_14\,
            ltout => OPEN,
            carryin => \c0.data_cry_13\,
            carryout => \c0.data_cry_14\,
            clk => \N__19661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_15_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10137\,
            in2 => \_gnd_net_\,
            in3 => \N__9643\,
            lcout => \c0.dataZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__4_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13663\,
            lcout => \c0.data_in_3_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19586\,
            ce => \N__17715\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__0_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14409\,
            lcout => \c0.data_in_3_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19586\,
            ce => \N__17715\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__7_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11241\,
            lcout => \c0.data_in_3_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19586\,
            ce => \N__17715\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__0_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12270\,
            lcout => \c0.data_in_4_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19586\,
            ce => \N__17715\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11012\,
            in1 => \N__10991\,
            in2 => \N__10956\,
            in3 => \N__12674\,
            lcout => \c0.i12_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__2_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12306\,
            lcout => \c0.data_in_2_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19593\,
            ce => \N__17718\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__5_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11049\,
            lcout => \c0.data_in_2_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19593\,
            ce => \N__17718\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__7_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13964\,
            lcout => \c0.data_in_2_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19593\,
            ce => \N__17718\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__2_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12675\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_1_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19593\,
            ce => \N__17718\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__2_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11181\,
            lcout => \c0.data_in_3_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19593\,
            ce => \N__17718\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11072\,
            in1 => \N__12305\,
            in2 => \N__12388\,
            in3 => \N__15842\,
            lcout => \c0.i12_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_2_c_RNO_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11099\,
            in1 => \N__12323\,
            in2 => \N__12504\,
            in3 => \N__13766\,
            lcout => \c0.i12_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__4_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11196\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_1_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19598\,
            ce => \N__17719\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__5_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11013\,
            lcout => \c0.data_in_1_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19598\,
            ce => \N__17719\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__7_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_1_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19598\,
            ce => \N__17719\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__0_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11079\,
            lcout => \c0.data_in_2_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19598\,
            ce => \N__17719\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__5_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_0_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19598\,
            ce => \N__17719\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__4_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12357\,
            lcout => \c0.data_in_2_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19598\,
            ce => \N__17719\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_5_c_RNO_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11195\,
            in1 => \N__11360\,
            in2 => \N__13617\,
            in3 => \N__13709\,
            lcout => \c0.i12_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__7_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11100\,
            lcout => \c0.data_in_0_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19603\,
            ce => \N__17721\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__0_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12500\,
            lcout => \c0.data_in_1_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19603\,
            ce => \N__17721\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__1_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11361\,
            lcout => \c0.data_in_1_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19603\,
            ce => \N__17721\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__3_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10996\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_1_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19603\,
            ce => \N__17721\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__0_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10242\,
            lcout => \c0.data_in_0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19603\,
            ce => \N__17721\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12693\,
            in1 => \N__14430\,
            in2 => \N__15933\,
            in3 => \N__11142\,
            lcout => \c0.i12_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__2_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15929\,
            lcout => \c0.data_in_0_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19603\,
            ce => \N__17721\,
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_RNO_0_2_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10486\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9734\,
            lcout => OPEN,
            ltout => \c0.tx.r_Bit_Index_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_2_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000010010001000"
        )
    port map (
            in0 => \N__10570\,
            in1 => \N__10398\,
            in2 => \N__9715\,
            in3 => \N__10606\,
            lcout => \c0.tx.r_Bit_IndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_RNO_0_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10319\,
            in1 => \N__9822\,
            in2 => \_gnd_net_\,
            in3 => \N__9778\,
            lcout => OPEN,
            ltout => \c0.tx.r_Tx_Active_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011111111"
        )
    port map (
            in0 => \N__9703\,
            in1 => \_gnd_net_\,
            in2 => \N__9712\,
            in3 => \N__9709\,
            lcout => \c0.tx_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_RNI6GJO_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9936\,
            in2 => \_gnd_net_\,
            in3 => \N__9701\,
            lcout => \c0.byte_transmit_counter15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__9702\,
            in1 => \_gnd_net_\,
            in2 => \N__9947\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_transmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.N_90_ip_RNI1U1E_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9814\,
            in2 => \_gnd_net_\,
            in3 => \N__9856\,
            lcout => \c0.tx.N_90_ip_RNI1U1EZ0\,
            ltout => \c0.tx.N_90_ip_RNI1U1EZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10494\,
            in2 => \N__9691\,
            in3 => \N__9735\,
            lcout => \c0.tx.r_Bit_IndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_4_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10323\,
            in1 => \N__9902\,
            in2 => \_gnd_net_\,
            in3 => \N__9815\,
            lcout => \c0.tx.r_SM_Main_dup_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNO_0_0_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10318\,
            in1 => \N__10648\,
            in2 => \N__9957\,
            in3 => \N__10537\,
            lcout => \c0.tx.r_SM_Main_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_1_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001110000000000"
        )
    port map (
            in0 => \N__9736\,
            in1 => \N__10605\,
            in2 => \N__10503\,
            in3 => \N__10399\,
            lcout => \c0.tx.r_Bit_IndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNO_0_2_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__9901\,
            in1 => \N__10649\,
            in2 => \_gnd_net_\,
            in3 => \N__10538\,
            lcout => OPEN,
            ltout => \c0.tx.r_SM_Main_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_2_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__10468\,
            in1 => \N__9903\,
            in2 => \N__9886\,
            in3 => \N__9816\,
            lcout => \c0.tx.r_SM_Main_dup_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNIVDI71_2_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__9857\,
            in1 => \N__10647\,
            in2 => \N__9823\,
            in3 => \N__9771\,
            lcout => \c0.tx.r_SM_Main_RNIVDI71Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__7_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19624\,
            ce => 'H',
            sr => \N__16879\
        );

    \c0.data_out_2__4_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16960\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19624\,
            ce => 'H',
            sr => \N__16879\
        );

    \c0.data_out_1__7_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16959\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19624\,
            ce => 'H',
            sr => \N__16879\
        );

    \c0.data_out_0__0_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16955\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19624\,
            ce => 'H',
            sr => \N__16879\
        );

    \c0.data_out_0__1_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16956\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19624\,
            ce => 'H',
            sr => \N__16879\
        );

    \c0.data_out_0__4_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16957\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19624\,
            ce => 'H',
            sr => \N__16879\
        );

    \c0.data_out_2__7_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16961\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19624\,
            ce => 'H',
            sr => \N__16879\
        );

    \CONSTANT_ONE_LUT4_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_2_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14466\,
            in1 => \N__12086\,
            in2 => \_gnd_net_\,
            in3 => \N__13328\,
            lcout => \c0.nextCRC16_3_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNINVK01_8_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12637\,
            in1 => \N__13009\,
            in2 => \_gnd_net_\,
            in3 => \N__11862\,
            lcout => \c0.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIIQK01_7_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10895\,
            in1 => \N__11427\,
            in2 => \_gnd_net_\,
            in3 => \N__13327\,
            lcout => \c0.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIQ3DA1_20_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11513\,
            in1 => \N__14465\,
            in2 => \N__12090\,
            in3 => \N__14497\,
            lcout => \c0.nextCRC16_3_0_a2_6_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__1_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10674\,
            in1 => \N__10789\,
            in2 => \N__12850\,
            in3 => \N__10071\,
            lcout => \c0.data_out_7_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19639\,
            ce => \N__16832\,
            sr => \_gnd_net_\
        );

    \c0.d_2_RNI9INJ_33_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11762\,
            in2 => \_gnd_net_\,
            in3 => \N__11790\,
            lcout => \c0.N_24_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNID5VK2_21_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9998\,
            in1 => \N__11992\,
            in2 => \N__14873\,
            in3 => \N__10022\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIKDAK6_20_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10102\,
            in1 => \N__12013\,
            in2 => \N__10096\,
            in3 => \N__10083\,
            lcout => \c0.N_106\,
            ltout => \c0.N_106_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__7_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10822\,
            in2 => \N__10093\,
            in3 => \N__10788\,
            lcout => \c0.data_out_6_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19639\,
            ce => \N__16832\,
            sr => \_gnd_net_\
        );

    \c0.d_2_RNITDBK1_19_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10440\,
            in1 => \N__12803\,
            in2 => \N__13361\,
            in3 => \N__11588\,
            lcout => \c0.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__0_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10675\,
            in1 => \N__10717\,
            in2 => \N__10909\,
            in3 => \N__10072\,
            lcout => \c0.data_out_7_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19639\,
            ce => \N__16832\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__2_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13399\,
            in1 => \N__13485\,
            in2 => \N__10054\,
            in3 => \N__10005\,
            lcout => \c0.data_out_6_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19647\,
            ce => \N__16829\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__4_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10042\,
            lcout => \c0.d_2_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19647\,
            ce => \N__16829\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__1_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14874\,
            in1 => \N__10027\,
            in2 => \N__11998\,
            in3 => \N__10006\,
            lcout => \c0.data_out_6_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19653\,
            ce => \N__16827\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__0_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10186\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19653\,
            ce => \N__16827\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__6_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10174\,
            lcout => \c0.d_2_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19653\,
            ce => \N__16827\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__3_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10162\,
            lcout => \c0.d_2_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19653\,
            ce => \N__16827\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__2_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10150\,
            lcout => \c0.d_2_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19653\,
            ce => \N__16827\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__7_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10138\,
            lcout => \c0.d_2_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19653\,
            ce => \N__16827\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__4_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10126\,
            lcout => \c0.d_2_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19653\,
            ce => \N__16827\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__0_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10114\,
            lcout => \c0.d_2_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19662\,
            ce => \N__16825\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__0_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10931\,
            lcout => \c0.data_in_5_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19592\,
            ce => \N__17717\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__7_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12150\,
            lcout => \c0.data_in_4_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19592\,
            ce => \N__17717\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__3_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11230\,
            lcout => \c0.data_in_4_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19592\,
            ce => \N__17717\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__7_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13584\,
            lcout => \c0.data_in_5_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19592\,
            ce => \N__17717\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__2_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17761\,
            lcout => \c0.data_in_5_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19592\,
            ce => \N__17717\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__0_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17369\,
            lcout => \c0.data_in_6_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19592\,
            ce => \N__17717\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__1_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13640\,
            lcout => \c0.data_in_5_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19599\,
            ce => \N__17720\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__1_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12288\,
            lcout => \c0.data_in_4_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19599\,
            ce => \N__17720\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__1_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17337\,
            lcout => \c0.data_in_6_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19599\,
            ce => \N__17720\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__3_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12386\,
            lcout => \c0.data_in_2_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19599\,
            ce => \N__17720\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__3_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11386\,
            lcout => \c0.data_in_6_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19599\,
            ce => \N__17720\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__2_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12519\,
            lcout => \c0.data_in_4_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19599\,
            ce => \N__17720\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__1_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11031\,
            lcout => \c0.data_in_3_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19599\,
            ce => \N__17720\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__4_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10261\,
            lcout => \c0.d_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19604\,
            ce => \N__17185\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__3_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11381\,
            lcout => \c0.data_in_frame_7_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19604\,
            ce => \N__17185\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__0_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10243\,
            lcout => \c0.d_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19604\,
            ce => \N__17185\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__1_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13641\,
            lcout => \c0.data_in_frame_6_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19604\,
            ce => \N__17185\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__1_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15849\,
            lcout => \c0.data_in_2_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19612\,
            ce => \N__17724\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__3_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12139\,
            lcout => \c0.data_in_3_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19612\,
            ce => \N__17724\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__3_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10225\,
            lcout => \c0.data_in_7_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19612\,
            ce => \N__17724\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__7_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13552\,
            lcout => \c0.data_in_6_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19612\,
            ce => \N__17724\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__1_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10207\,
            lcout => \c0.data_in_7_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19612\,
            ce => \N__17724\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__0_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10420\,
            lcout => \c0.data_in_7_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19612\,
            ce => \N__17724\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__3_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11310\,
            lcout => \c0.data_in_5_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19612\,
            ce => \N__17724\,
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_5_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__13174\,
            in1 => \N__10566\,
            in2 => \N__11398\,
            in3 => \N__10599\,
            lcout => OPEN,
            ltout => \c0.tx.o_Tx_Serial_2_3_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_3_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10600\,
            in1 => \N__14299\,
            in2 => \N__10402\,
            in3 => \N__13156\,
            lcout => \c0.tx.o_Tx_Serial_RNO_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_0_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10397\,
            lcout => \c0.tx.N_390_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_4_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__10567\,
            in1 => \N__13096\,
            in2 => \N__11608\,
            in3 => \N__10601\,
            lcout => OPEN,
            ltout => \c0.tx.o_Tx_Serial_2_6_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_2_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10602\,
            in1 => \N__11404\,
            in2 => \N__10381\,
            in3 => \N__11440\,
            lcout => OPEN,
            ltout => \c0.tx.o_Tx_Serial_RNO_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_1_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__10498\,
            in1 => \N__10378\,
            in2 => \N__10372\,
            in3 => \N__10654\,
            lcout => OPEN,
            ltout => \c0.tx.o_Tx_Serial_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__10272\,
            in1 => \N__10356\,
            in2 => \N__10327\,
            in3 => \N__10324\,
            lcout => \PIN_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19625\,
            ce => 'H',
            sr => \N__10666\
        );

    \c0.tx.r_SM_Main_RNO_0_3_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10568\,
            in1 => \N__10603\,
            in2 => \N__10504\,
            in3 => \N__10653\,
            lcout => \c0.tx.r_SM_Main_recr_i_0_a2_0_2_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNO_1_2_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__10604\,
            in1 => \N__10569\,
            in2 => \N__10546\,
            in3 => \N__10502\,
            lcout => \c0.tx.r_SM_Main_recr_i_i_a2_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__5_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10834\,
            in1 => \N__10765\,
            in2 => \N__10450\,
            in3 => \N__11598\,
            lcout => \c0.data_out_7_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19633\,
            ce => \N__16835\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_5_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__15373\,
            in1 => \N__10459\,
            in2 => \N__15568\,
            in3 => \N__10846\,
            lcout => \c0.tx_data_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_3_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__10780\,
            in1 => \N__15558\,
            in2 => \N__14830\,
            in3 => \N__15371\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_3_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__15197\,
            in1 => \N__15652\,
            in2 => \N__10453\,
            in3 => \N__10426\,
            lcout => \c0.tx_data_1_0_i_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_3_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__10446\,
            in1 => \N__15557\,
            in2 => \N__10711\,
            in3 => \N__15370\,
            lcout => \c0.tx_data_RNO_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_3_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__15372\,
            in1 => \N__11711\,
            in2 => \N__15567\,
            in3 => \N__10900\,
            lcout => \c0.tx_data_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_2_0_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11824\,
            in1 => \N__11710\,
            in2 => \_gnd_net_\,
            in3 => \N__11741\,
            lcout => \c0.nextCRC16_3_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_2_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11831\,
            in1 => \N__12832\,
            in2 => \N__12942\,
            in3 => \N__11649\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_0_a2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__2_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10803\,
            in1 => \N__15030\,
            in2 => \N__10750\,
            in3 => \N__11671\,
            lcout => \c0.data_out_7_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19640\,
            ce => \N__16833\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__6_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10747\,
            lcout => \c0.d_2_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19640\,
            ce => \N__16833\,
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIFMJ01_45_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12984\,
            in1 => \N__14934\,
            in2 => \_gnd_net_\,
            in3 => \N__12864\,
            lcout => \c0.N_99\,
            ltout => \c0.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_3_0_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14993\,
            in1 => \N__13039\,
            in2 => \N__10729\,
            in3 => \N__10802\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_0_a2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_1_0_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10726\,
            in1 => \N__12775\,
            in2 => \N__10720\,
            in3 => \N__14793\,
            lcout => \c0.nextCRC16_3_0_a2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIDLMJ_16_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14959\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12602\,
            lcout => \c0.N_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIM3JT_12_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12035\,
            in1 => \N__14894\,
            in2 => \_gnd_net_\,
            in3 => \N__11947\,
            lcout => \c0.N_81\,
            ltout => \c0.N_81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNII92R1_27_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10710\,
            in1 => \N__13136\,
            in2 => \N__10678\,
            in3 => \N__14819\,
            lcout => \c0.N_105\,
            ltout => \c0.N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__5_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12933\,
            in2 => \N__10849\,
            in3 => \N__13404\,
            lcout => \c0.data_out_6_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19648\,
            ce => \N__16830\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_1_7_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11740\,
            in1 => \N__11835\,
            in2 => \N__12941\,
            in3 => \N__14789\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_0_a2_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_7_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10816\,
            in1 => \N__11666\,
            in2 => \N__10837\,
            in3 => \N__10833\,
            lcout => \c0.nextCRC16_3_0_a2_5_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_2_7_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14895\,
            in1 => \N__13135\,
            in2 => \N__11955\,
            in3 => \N__14818\,
            lcout => \c0.nextCRC16_3_0_a2_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIJ2812_44_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14747\,
            in1 => \N__13293\,
            in2 => \N__13448\,
            in3 => \N__10761\,
            lcout => \c0.N_95\,
            ltout => \c0.N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIJDOU2_14_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15031\,
            in2 => \N__10810\,
            in3 => \N__10807\,
            lcout => \c0.nextCRC16_3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__7_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19654\,
            ce => 'H',
            sr => \N__16877\
        );

    \c0.data_out_0__3_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17019\,
            lcout => \c0.d_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19654\,
            ce => 'H',
            sr => \N__16877\
        );

    \c0.d_2_RNI6EK01_3_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12114\,
            in1 => \N__11638\,
            in2 => \_gnd_net_\,
            in3 => \N__10776\,
            lcout => \c0.N_75\,
            ltout => \c0.N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_0_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13441\,
            in2 => \N__10912\,
            in3 => \N__14748\,
            lcout => \c0.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__2_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17018\,
            lcout => \c0.d_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19654\,
            ce => 'H',
            sr => \N__16877\
        );

    \c0.data_out_6__RNO_0_4_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11940\,
            in2 => \_gnd_net_\,
            in3 => \N__13395\,
            lcout => \c0.nextCRC16_3_3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_6_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12113\,
            in2 => \_gnd_net_\,
            in3 => \N__10894\,
            lcout => \c0.un144_newcrc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__1_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.d_2_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19668\,
            ce => 'H',
            sr => \N__16873\
        );

    \c0.data_out_3__0_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.d_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19668\,
            ce => 'H',
            sr => \N__16873\
        );

    \c0.data_in_7__7_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10870\,
            lcout => \c0.data_in_7_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19605\,
            ce => \N__17722\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__5_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11877\,
            lcout => \c0.data_in_4_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19605\,
            ce => \N__17722\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__5_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11878\,
            lcout => \c0.d_4_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19597\,
            ce => \N__17177\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__6_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16087\,
            lcout => \c0.d_4_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19597\,
            ce => \N__17177\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__0_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10932\,
            lcout => \c0.data_in_frame_6_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19597\,
            ce => \N__17177\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__5_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11020\,
            lcout => \c0.d_4_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19597\,
            ce => \N__17177\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__2_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17757\,
            lcout => \c0.data_in_frame_6_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19597\,
            ce => \N__17177\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__3_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10992\,
            lcout => \c0.d_4_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19597\,
            ce => \N__17177\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__2_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17775\,
            lcout => \c0.data_in_frame_7_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19597\,
            ce => \N__17177\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNINGK21_21_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17582\,
            in1 => \N__18869\,
            in2 => \N__14394\,
            in3 => \N__13688\,
            lcout => \c0.N_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__7_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10975\,
            lcout => \c0.d_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19606\,
            ce => \N__17181\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__7_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10957\,
            lcout => \c0.d_4_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19606\,
            ce => \N__17181\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIT2KP_20_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13689\,
            in1 => \N__12193\,
            in2 => \N__10933\,
            in3 => \N__17960\,
            lcout => \c0.un1_data_in_6__0_0_a2_5_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__4_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11203\,
            lcout => \c0.d_4_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19606\,
            ce => \N__17181\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__2_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19606\,
            ce => \N__17181\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIQ7PC_23_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14390\,
            in1 => \N__16437\,
            in2 => \N__17649\,
            in3 => \N__11303\,
            lcout => \c0.un1_data_in_6__3_0_a2_5_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__5_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11166\,
            lcout => \c0.d_4_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19606\,
            ce => \N__17181\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__0_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11149\,
            lcout => \c0.d_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19613\,
            ce => \N__17182\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__3_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11131\,
            lcout => \c0.d_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19613\,
            ce => \N__17182\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__7_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11104\,
            lcout => \c0.d_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19613\,
            ce => \N__17182\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__0_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11083\,
            lcout => \c0.d_4_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19613\,
            ce => \N__17182\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__5_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11056\,
            lcout => \c0.d_4_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19613\,
            ce => \N__17182\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__1_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11032\,
            lcout => \c0.d_4_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19613\,
            ce => \N__17182\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__7_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11245\,
            lcout => \c0.d_4_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19613\,
            ce => \N__17182\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__3_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11226\,
            lcout => \c0.d_4_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19613\,
            ce => \N__17182\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI5L571_45_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17676\,
            in1 => \N__12738\,
            in2 => \N__11284\,
            in3 => \N__14612\,
            lcout => \c0.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIH9JJ_4_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12198\,
            in1 => \N__18054\,
            in2 => \_gnd_net_\,
            in3 => \N__12472\,
            lcout => \c0.N_108\,
            ltout => \c0.N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNICGS41_17_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__11281\,
            in1 => \_gnd_net_\,
            in2 => \N__11215\,
            in3 => \N__14613\,
            lcout => OPEN,
            ltout => \c0.N_122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIJUS53_16_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16545\,
            in1 => \N__12259\,
            in2 => \N__11212\,
            in3 => \N__12550\,
            lcout => \c0.un1_data_in_7__1_0_a2_24_a2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIVCPC_26_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13927\,
            in1 => \N__17606\,
            in2 => \N__13583\,
            in3 => \N__16046\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__7_0_a2_17_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIIAP41_26_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__16301\,
            in1 => \_gnd_net_\,
            in2 => \N__11209\,
            in3 => \N__13801\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__7_0_a2_17_a2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIP5RG3_15_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16501\,
            in1 => \N__16546\,
            in2 => \N__11206\,
            in3 => \N__16157\,
            lcout => \c0.un1_data_in_6__7_0_a2_17_a2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIN7VG_47_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11282\,
            in1 => \N__18095\,
            in2 => \N__11385\,
            in3 => \N__17514\,
            lcout => \c0.un1_data_in_7__3_0_a2_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__1_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11362\,
            lcout => \c0.d_4_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19626\,
            ce => \N__17187\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__6_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11344\,
            lcout => \c0.d_4_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19626\,
            ce => \N__17187\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_3_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__18361\,
            in1 => \N__11290\,
            in2 => \N__11323\,
            in3 => \N__18571\,
            lcout => \c0.tx2_data_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__3_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11311\,
            lcout => \c0.data_in_frame_6_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19626\,
            ce => \N__17187\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_1_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__11283\,
            in1 => \N__18572\,
            in2 => \N__18374\,
            in3 => \N__15826\,
            lcout => \c0.tx2_data_RNO_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_1_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__16633\,
            in1 => \N__18715\,
            in2 => \N__11263\,
            in3 => \N__18799\,
            lcout => OPEN,
            ltout => \c0.m161_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_1_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__18716\,
            in1 => \N__16597\,
            in2 => \N__11254\,
            in3 => \N__11251\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19634\,
            ce => \N__19978\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_1_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__15985\,
            in1 => \N__18578\,
            in2 => \N__18376\,
            in3 => \N__12479\,
            lcout => \c0.tx2_data_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_2_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__16336\,
            in1 => \N__18370\,
            in2 => \N__18594\,
            in3 => \N__12199\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_2_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__11458\,
            in1 => \N__14335\,
            in2 => \N__11485\,
            in3 => \N__18717\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19634\,
            ce => \N__19978\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_2_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__18577\,
            in1 => \N__11482\,
            in2 => \N__11470\,
            in3 => \N__18369\,
            lcout => \c0.tx2_data_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_7_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__11650\,
            in1 => \N__15565\,
            in2 => \N__11997\,
            in3 => \N__15374\,
            lcout => \c0.tx_data_RNO_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_3_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__11452\,
            in1 => \N__13216\,
            in2 => \N__15212\,
            in3 => \N__11446\,
            lcout => \c0.tx.r_Tx_DataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19641\,
            ce => \N__14279\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_7_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__11431\,
            in1 => \N__15566\,
            in2 => \N__11749\,
            in3 => \N__15375\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_7_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__15198\,
            in1 => \N__15658\,
            in2 => \N__11416\,
            in3 => \N__11413\,
            lcout => OPEN,
            ltout => \c0.tx_data_1_0_i_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_7_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__13339\,
            in1 => \N__15199\,
            in2 => \N__11407\,
            in3 => \N__12559\,
            lcout => \c0.tx.r_Tx_DataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19641\,
            ce => \N__14279\,
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_4_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__13282\,
            in1 => \N__11890\,
            in2 => \N__15213\,
            in3 => \N__11536\,
            lcout => \c0.tx.r_Tx_DataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19641\,
            ce => \N__14279\,
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_5_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__12961\,
            in1 => \N__11614\,
            in2 => \N__15214\,
            in3 => \N__12751\,
            lcout => \c0.tx.r_Tx_DataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19641\,
            ce => \N__14279\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_1_6_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12811\,
            in1 => \N__12879\,
            in2 => \N__11530\,
            in3 => \N__11599\,
            lcout => OPEN,
            ltout => \c0.un144_newcrc_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__6_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11572\,
            in1 => \N__14749\,
            in2 => \N__11563\,
            in3 => \N__12606\,
            lcout => \c0.data_out_7_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19649\,
            ce => \N__16831\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_6_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15346\,
            in1 => \N__11545\,
            in2 => \N__11560\,
            in3 => \N__15531\,
            lcout => \c0.tx_data_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__6_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12886\,
            in1 => \N__11551\,
            in2 => \_gnd_net_\,
            in3 => \N__11712\,
            lcout => \c0.data_out_6_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19649\,
            ce => \N__16831\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_4_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15345\,
            in1 => \N__12878\,
            in2 => \N__14902\,
            in3 => \N__15532\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_4_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__15166\,
            in1 => \N__15657\,
            in2 => \N__11539\,
            in3 => \N__11497\,
            lcout => \c0.tx_data_1_0_i_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_4_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__15344\,
            in1 => \N__12828\,
            in2 => \N__11529\,
            in3 => \N__15530\,
            lcout => \c0.tx_data_RNO_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__4_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11491\,
            in1 => \N__14958\,
            in2 => \N__15001\,
            in3 => \N__11797\,
            lcout => \c0.data_out_7_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19655\,
            ce => \N__16828\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_0_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__11866\,
            in1 => \N__15511\,
            in2 => \N__11842\,
            in3 => \N__15341\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_0_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__15186\,
            in1 => \N__15656\,
            in2 => \N__11806\,
            in3 => \N__11803\,
            lcout => \c0.tx_data_1_0_i_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_0_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__14957\,
            in1 => \N__15510\,
            in2 => \N__12091\,
            in3 => \N__15340\,
            lcout => \c0.tx_data_RNO_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_1_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__15342\,
            in1 => \N__12036\,
            in2 => \N__15540\,
            in3 => \N__11796\,
            lcout => \c0.tx_data_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_2_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__12934\,
            in1 => \N__15515\,
            in2 => \N__11779\,
            in3 => \N__15343\,
            lcout => \c0.tx_data_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_3_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13452\,
            in2 => \_gnd_net_\,
            in3 => \N__11748\,
            lcout => OPEN,
            ltout => \c0.un105_newcrc_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__3_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11620\,
            in1 => \N__11713\,
            in2 => \N__11674\,
            in3 => \N__11667\,
            lcout => \c0.data_out_7_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19663\,
            ce => \N__16826\,
            sr => \_gnd_net_\
        );

    \c0.d_2_RNI9GJ01_29_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14997\,
            in1 => \N__16905\,
            in2 => \_gnd_net_\,
            in3 => \N__13049\,
            lcout => \c0.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_1_3_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13365\,
            in1 => \N__12121\,
            in2 => \N__14938\,
            in3 => \N__11645\,
            lcout => \c0.un105_newcrc_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_0_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__12120\,
            in1 => \N__15516\,
            in2 => \N__11959\,
            in3 => \N__15332\,
            lcout => \c0.tx_data_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_1_4_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14829\,
            in1 => \N__15706\,
            in2 => \N__12082\,
            in3 => \N__12641\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_4_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__4_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14794\,
            in1 => \N__12049\,
            in2 => \N__12043\,
            in3 => \N__12040\,
            lcout => \c0.data_out_6_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19669\,
            ce => \N__16824\,
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIGMI01_10_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13400\,
            in1 => \N__15705\,
            in2 => \_gnd_net_\,
            in3 => \N__13489\,
            lcout => \c0.N_94\,
            ltout => \c0.N_94_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__3_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12642\,
            in1 => \N__11917\,
            in2 => \N__12001\,
            in3 => \N__13020\,
            lcout => \c0.data_out_6_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19669\,
            ce => \N__16824\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_3_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11996\,
            in1 => \N__13140\,
            in2 => \_gnd_net_\,
            in3 => \N__11954\,
            lcout => \c0.nextCRC16_3_0_a2_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_4_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__15471\,
            in1 => \N__11911\,
            in2 => \N__11905\,
            in3 => \N__15334\,
            lcout => \c0.tx_data_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_5__5_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17299\,
            lcout => \c0.data_in_5_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19614\,
            ce => \N__17725\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__4_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12238\,
            lcout => \c0.data_in_7_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19614\,
            ce => \N__17725\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__2_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12217\,
            lcout => \c0.data_in_7_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19614\,
            ce => \N__17725\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__4_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12537\,
            lcout => \c0.data_in_4_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19614\,
            ce => \N__17725\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__4_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16015\,
            lcout => \c0.data_in_5_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19614\,
            ce => \N__17725\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIJLQL_19_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14628\,
            in1 => \N__14700\,
            in2 => \N__13750\,
            in3 => \N__17504\,
            lcout => \c0.N_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI6FQT_21_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17904\,
            in1 => \N__13903\,
            in2 => \N__13541\,
            in3 => \N__17583\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__7_0_a2_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI675O1_33_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12194\,
            in1 => \N__12480\,
            in2 => \N__12169\,
            in3 => \N__12426\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__7_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI8SR93_20_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__12166\,
            in1 => \N__13732\,
            in2 => \N__12157\,
            in3 => \N__16403\,
            lcout => \c0.m163_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__7_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12154\,
            lcout => \c0.d_4_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19602\,
            ce => \N__17174\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__3_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12138\,
            lcout => \c0.d_4_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19602\,
            ce => \N__17174\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIO7RC_40_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16183\,
            in1 => \N__17984\,
            in2 => \N__17221\,
            in3 => \N__18174\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI240O_40_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12251\,
            in2 => \N__12361\,
            in3 => \N__13797\,
            lcout => \c0.un1_data_in_6__6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__4_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19615\,
            ce => \N__17178\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI1VL6_13_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17922\,
            in1 => \N__16039\,
            in2 => \_gnd_net_\,
            in3 => \N__15962\,
            lcout => \c0.N_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__5_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12331\,
            lcout => \c0.d_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19615\,
            ce => \N__17178\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__2_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12310\,
            lcout => \c0.d_4_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19615\,
            ce => \N__17178\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__1_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12292\,
            lcout => \c0.d_4_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19615\,
            ce => \N__17178\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__0_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12277\,
            lcout => \c0.d_4_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19615\,
            ce => \N__17178\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI1LAI2_12_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16302\,
            in1 => \N__12258\,
            in2 => \N__12400\,
            in3 => \N__16161\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__0_0_a2_1_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI20TA7_15_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16505\,
            in1 => \N__16544\,
            in2 => \N__12433\,
            in3 => \N__12409\,
            lcout => \c0.un1_data_in_7__0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIJ66B_11_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18818\,
            in1 => \N__14579\,
            in2 => \N__16438\,
            in3 => \N__13883\,
            lcout => \c0.N_121\,
            ltout => \c0.N_121_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNITCL32_11_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13833\,
            in2 => \N__12430\,
            in3 => \N__12427\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__7_0_a2_17_a2_4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIV4MJ3_10_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15892\,
            in1 => \N__12445\,
            in2 => \N__12412\,
            in3 => \N__16404\,
            lcout => \c0.N_136\,
            ltout => \c0.N_136_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIK2SL3_14_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__16272\,
            in1 => \_gnd_net_\,
            in2 => \N__12403\,
            in3 => \_gnd_net_\,
            lcout => \c0.un1_data_in_7__1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIG6H4_39_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17465\,
            in2 => \_gnd_net_\,
            in3 => \N__18173\,
            lcout => \c0.N_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIH0UG_12_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14667\,
            in1 => \N__16184\,
            in2 => \N__17370\,
            in3 => \N__18036\,
            lcout => \c0.un1_data_in_7__0_0_a2_1_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__3_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12387\,
            lcout => \c0.d_4_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19627\,
            ce => \N__17183\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIQ3V8_12_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14666\,
            in1 => \N__16328\,
            in2 => \N__13934\,
            in3 => \N__18035\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__1_0_a2_24_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIQ7KN_16_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17993\,
            in1 => \N__17333\,
            in2 => \N__12553\,
            in3 => \N__18849\,
            lcout => \c0.un1_data_in_7__1_0_a2_24_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__4_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12544\,
            lcout => \c0.d_4_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19627\,
            ce => \N__17183\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__2_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12526\,
            lcout => \c0.d_4_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19627\,
            ce => \N__17183\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__0_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19627\,
            ce => \N__17183\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIA0HJ_0_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18094\,
            in1 => \N__18894\,
            in2 => \_gnd_net_\,
            in3 => \N__18848\,
            lcout => \c0.N_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI34PL_16_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18096\,
            in1 => \N__18847\,
            in2 => \N__12481\,
            in3 => \N__14611\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI6DG41_18_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12657\,
            in1 => \N__15750\,
            in2 => \N__12448\,
            in3 => \N__13935\,
            lcout => \c0.un1_data_in_7__4_0_a2_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIABPL_18_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17964\,
            in1 => \N__12656\,
            in2 => \N__16371\,
            in3 => \N__17900\,
            lcout => \c0.N_124\,
            ltout => \c0.N_124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_7__RNIBJH41_6_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17251\,
            in1 => \N__18401\,
            in2 => \N__12436\,
            in3 => \N__14709\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__6_0_a2_5_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIDD8G3_18_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001000"
        )
    port map (
            in0 => \N__12745\,
            in1 => \N__13942\,
            in2 => \N__12727\,
            in3 => \N__12724\,
            lcout => \c0.m163_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__3_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12718\,
            lcout => \c0.d_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19635\,
            ce => \N__17186\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__5_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12700\,
            lcout => \c0.d_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19635\,
            ce => \N__17186\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_7_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__13675\,
            in1 => \N__18714\,
            in2 => \N__14374\,
            in3 => \N__18797\,
            lcout => \c0.m60_0_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_2_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__18576\,
            in1 => \N__16050\,
            in2 => \N__12661\,
            in3 => \N__18354\,
            lcout => \c0.tx2_data_RNO_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__2_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12682\,
            lcout => \c0.d_4_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19642\,
            ce => \N__17188\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_6_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__15533\,
            in1 => \N__14983\,
            in2 => \N__14464\,
            in3 => \N__15365\,
            lcout => \c0.tx_data_RNO_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_6_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15368\,
            in1 => \N__12643\,
            in2 => \N__12613\,
            in3 => \N__15537\,
            lcout => \c0.tx_data_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_7_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__15536\,
            in1 => \N__12586\,
            in2 => \N__12574\,
            in3 => \N__15369\,
            lcout => \c0.tx_data_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_5_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__15367\,
            in1 => \N__15535\,
            in2 => \N__13021\,
            in3 => \N__12985\,
            lcout => \c0.tx_data_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_6_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15366\,
            in1 => \N__14502\,
            in2 => \N__15026\,
            in3 => \N__15534\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_6_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__15165\,
            in1 => \N__15651\,
            in2 => \N__12955\,
            in3 => \N__12952\,
            lcout => \c0.tx_data_1_0_i_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIK3C71_13_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14775\,
            in1 => \N__12827\,
            in2 => \N__12946\,
            in3 => \N__12767\,
            lcout => \c0.nextCRC16_3_3_1\,
            ltout => \c0.nextCRC16_3_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_1_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12880\,
            in1 => \N__13054\,
            in2 => \N__12853\,
            in3 => \N__14926\,
            lcout => \c0.nextCRC16_3_0_a2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__5_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17006\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19656\,
            ce => 'H',
            sr => \N__16878\
        );

    \c0.data_out_3__4_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19656\,
            ce => 'H',
            sr => \N__16878\
        );

    \c0.tx_data_RNO_3_5_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__12810\,
            in1 => \N__15556\,
            in2 => \N__12774\,
            in3 => \N__15339\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_5_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__15163\,
            in1 => \N__15640\,
            in2 => \N__12754\,
            in3 => \N__13204\,
            lcout => \c0.tx_data_1_0_i_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_5_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__16909\,
            in1 => \N__15555\,
            in2 => \N__14866\,
            in3 => \N__15338\,
            lcout => \c0.tx_data_RNO_4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_0_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__13198\,
            in1 => \N__13186\,
            in2 => \N__15209\,
            in3 => \N__13180\,
            lcout => \c0.tx.r_Tx_DataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19664\,
            ce => \N__14283\,
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_2_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__13060\,
            in1 => \N__13162\,
            in2 => \N__15210\,
            in3 => \N__13414\,
            lcout => \c0.tx.r_Tx_DataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19664\,
            ce => \N__14283\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_1_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__14933\,
            in1 => \N__15517\,
            in2 => \N__13144\,
            in3 => \N__15364\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_1_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__15650\,
            in1 => \N__15187\,
            in2 => \N__13108\,
            in3 => \N__13459\,
            lcout => OPEN,
            ltout => \c0.tx_data_1_0_i_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_1_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__13105\,
            in1 => \N__15164\,
            in2 => \N__13099\,
            in3 => \N__13246\,
            lcout => \c0.tx.r_Tx_DataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19664\,
            ce => \N__14283\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_2_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__15289\,
            in1 => \N__13084\,
            in2 => \N__15539\,
            in3 => \N__13072\,
            lcout => \c0.tx_data_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_2_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__14776\,
            in1 => \N__15500\,
            in2 => \N__14743\,
            in3 => \N__15284\,
            lcout => \c0.tx_data_RNO_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_1_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__15286\,
            in1 => \N__13050\,
            in2 => \N__15538\,
            in3 => \N__13484\,
            lcout => \c0.tx_data_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_2_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__15704\,
            in1 => \N__15503\,
            in2 => \N__13453\,
            in3 => \N__15285\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_2_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__15167\,
            in1 => \N__15631\,
            in2 => \N__13423\,
            in3 => \N__13420\,
            lcout => \c0.tx_data_1_0_i_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_7_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__13408\,
            in1 => \N__15502\,
            in2 => \N__13366\,
            in3 => \N__15288\,
            lcout => \c0.tx_data_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_4_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__13330\,
            in1 => \N__15501\,
            in2 => \N__13303\,
            in3 => \N__15287\,
            lcout => \c0.tx_data_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_1_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__15473\,
            in1 => \N__13270\,
            in2 => \N__13261\,
            in3 => \N__15333\,
            lcout => \c0.tx_data_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNI7Q6P_6_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15676\,
            in2 => \_gnd_net_\,
            in3 => \N__15682\,
            lcout => OPEN,
            ltout => \c0.m2_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNIQP0V1_3_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13594\,
            in1 => \N__15664\,
            in2 => \N__13237\,
            in3 => \N__15670\,
            lcout => \c0.N_132_mux\,
            ltout => \c0.N_132_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_3_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__13234\,
            in1 => \N__13228\,
            in2 => \N__13219\,
            in3 => \N__15472\,
            lcout => \c0.tx_data_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19676\,
            ce => \N__15075\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15474\,
            in2 => \_gnd_net_\,
            in3 => \N__15335\,
            lcout => \c0.byte_transmit_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19676\,
            ce => \N__15075\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_2_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__15336\,
            in1 => \N__15133\,
            in2 => \N__15528\,
            in3 => \N__15633\,
            lcout => \c0.byte_transmit_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19676\,
            ce => \N__15075\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__4_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15746\,
            lcout => \c0.data_in_frame_7_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19619\,
            ce => \N__17172\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_7_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__13558\,
            in1 => \N__18347\,
            in2 => \N__13522\,
            in3 => \N__18590\,
            lcout => \c0.tx2_data_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__7_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13588\,
            lcout => \c0.data_in_frame_6_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19610\,
            ce => \N__17173\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__7_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13548\,
            lcout => \c0.data_in_frame_7_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19610\,
            ce => \N__17173\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_6_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__18591\,
            in1 => \N__16268\,
            in2 => \N__18372\,
            in3 => \N__13749\,
            lcout => \c0.tx2_data_RNO_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__6_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13513\,
            lcout => \c0.d_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19610\,
            ce => \N__17173\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIUBBH_6_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13748\,
            in2 => \_gnd_net_\,
            in3 => \N__14704\,
            lcout => \c0.N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__6_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13723\,
            lcout => \c0.d_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19610\,
            ce => \N__17173\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_7_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__18589\,
            in1 => \N__16516\,
            in2 => \N__18371\,
            in3 => \N__13696\,
            lcout => \c0.tx2_data_RNO_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__4_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13659\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19620\,
            ce => \N__17175\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIJ8G4_36_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13901\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17648\,
            lcout => OPEN,
            ltout => \c0.N_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_6__RNIKD2F_1_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13642\,
            in1 => \N__16435\,
            in2 => \N__13621\,
            in3 => \N__14705\,
            lcout => \c0.un1_data_in_6__1_0_a2_4_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI76N6_22_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13900\,
            in1 => \N__17647\,
            in2 => \_gnd_net_\,
            in3 => \N__18117\,
            lcout => \c0.N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__6_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13618\,
            lcout => \c0.d_4_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19620\,
            ce => \N__17175\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__6_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16098\,
            lcout => \c0.d_4_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19620\,
            ce => \N__17175\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_4_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__18588\,
            in1 => \N__13936\,
            in2 => \N__18375\,
            in3 => \N__13902\,
            lcout => \c0.tx2_data_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_6_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__16436\,
            in1 => \N__18587\,
            in2 => \N__16372\,
            in3 => \N__18365\,
            lcout => \c0.tx2_data_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI23VN_11_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13793\,
            in1 => \N__14586\,
            in2 => \N__13810\,
            in3 => \N__13884\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNITNPS1_11_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000001001"
        )
    port map (
            in0 => \N__13885\,
            in1 => \N__13870\,
            in2 => \N__13858\,
            in3 => \N__15891\,
            lcout => OPEN,
            ltout => \c0.m163_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_6__RNIAQG64_1_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__13855\,
            in1 => \N__13849\,
            in2 => \N__13843\,
            in3 => \N__13840\,
            lcout => OPEN,
            ltout => \c0.m163_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIFGESA_24_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16282\,
            in1 => \N__16381\,
            in2 => \N__13822\,
            in3 => \N__13819\,
            lcout => \c0.m163_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIN4PC_25_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17291\,
            in1 => \N__14665\,
            in2 => \N__15980\,
            in3 => \N__15818\,
            lcout => \c0.un1_data_in_6__5_0_a2_5_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI9TE4_12_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16327\,
            in2 => \_gnd_net_\,
            in3 => \N__18034\,
            lcout => \c0.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__4_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13777\,
            lcout => \c0.d_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19628\,
            ce => \N__17179\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIC7M21_1_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18402\,
            in1 => \N__16245\,
            in2 => \N__16675\,
            in3 => \N__14365\,
            lcout => \c0.N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNIGB9N4_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000000000"
        )
    port map (
            in0 => \N__14032\,
            in1 => \N__14026\,
            in2 => \N__15946\,
            in3 => \N__19287\,
            lcout => OPEN,
            ltout => \c0.m163_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIGIT3F_14_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111101111"
        )
    port map (
            in0 => \N__14020\,
            in1 => \N__14011\,
            in2 => \N__14002\,
            in3 => \N__13999\,
            lcout => OPEN,
            ltout => \c0.m163_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI7JOT41_15_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__13993\,
            in1 => \N__16132\,
            in2 => \N__13987\,
            in3 => \N__13984\,
            lcout => \c0.N_164_0\,
            ltout => \c0.N_164_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_RNIG45P61_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__19339\,
            in1 => \N__20013\,
            in2 => \N__13978\,
            in3 => \N__17809\,
            lcout => \c0.N_173_0\,
            ltout => \c0.N_173_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_active_RNIABU671_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19721\,
            in2 => \N__13975\,
            in3 => \_gnd_net_\,
            lcout => \c0.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIM5UG_19_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18400\,
            in1 => \N__16243\,
            in2 => \N__17275\,
            in3 => \N__14640\,
            lcout => \c0.un1_data_in_7__5_0_a2_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__7_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13972\,
            lcout => \c0.d_4_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19643\,
            ce => \N__17184\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIB3JJ_2_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18399\,
            in1 => \N__16242\,
            in2 => \_gnd_net_\,
            in3 => \N__14360\,
            lcout => \c0.d_4_RNIB3JJZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__2_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14437\,
            lcout => \c0.d_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19643\,
            ce => \N__17184\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__0_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14419\,
            lcout => \c0.d_4_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19643\,
            ce => \N__17184\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_7_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__16244\,
            in1 => \N__18305\,
            in2 => \N__18570\,
            in3 => \N__14398\,
            lcout => \c0.tx2_data_RNO_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_2_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__15910\,
            in1 => \N__18514\,
            in2 => \N__18353\,
            in3 => \N__14361\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_2_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__18657\,
            in1 => \N__14347\,
            in2 => \N__14338\,
            in3 => \N__18784\,
            lcout => \c0.m131_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_6_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__14323\,
            in1 => \N__14311\,
            in2 => \N__15211\,
            in3 => \N__14305\,
            lcout => \c0.tx.r_Tx_DataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19650\,
            ce => \N__14287\,
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNIC9J951_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19342\,
            in2 => \_gnd_net_\,
            in3 => \N__18142\,
            lcout => \c0.tx2_transmit_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_RNIRD3K_1_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__14247\,
            in1 => \N__14185\,
            in2 => \_gnd_net_\,
            in3 => \N__14124\,
            lcout => \c0.rx.N_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_3_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__16198\,
            in1 => \N__18357\,
            in2 => \N__18595\,
            in3 => \N__14713\,
            lcout => \c0.tx2_data_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_3_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__18355\,
            in1 => \N__14674\,
            in2 => \N__14647\,
            in3 => \N__18582\,
            lcout => \c0.tx2_data_RNO_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_3_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__18586\,
            in1 => \N__14617\,
            in2 => \N__14593\,
            in3 => \N__18356\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_3_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__18798\,
            in1 => \N__14566\,
            in2 => \N__14560\,
            in3 => \N__18719\,
            lcout => OPEN,
            ltout => \c0.m105_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_3_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__14557\,
            in1 => \N__18721\,
            in2 => \N__14551\,
            in3 => \N__14548\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19657\,
            ce => \N__19973\,
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_3_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__14509\,
            in1 => \N__14536\,
            in2 => \_gnd_net_\,
            in3 => \N__19822\,
            lcout => \c0.tx2.o_Tx_Serial_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_7_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__18720\,
            in1 => \N__17452\,
            in2 => \N__14530\,
            in3 => \N__14515\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19657\,
            ce => \N__19973\,
            sr => \_gnd_net_\
        );

    \c0.data_out_0__6_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17008\,
            lcout => \c0.d_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19665\,
            ce => 'H',
            sr => \N__16875\
        );

    \c0.data_out_2__6_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17010\,
            lcout => \c0.d_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19665\,
            ce => 'H',
            sr => \N__16875\
        );

    \c0.data_out_1__6_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17009\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19665\,
            ce => 'H',
            sr => \N__16875\
        );

    \c0.data_out_3__6_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17011\,
            lcout => \c0.d_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19665\,
            ce => 'H',
            sr => \N__16875\
        );

    \c0.data_out_2__0_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17087\,
            lcout => \c0.d_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19670\,
            ce => 'H',
            sr => \N__16874\
        );

    \c0.data_out_2__1_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19670\,
            ce => 'H',
            sr => \N__16874\
        );

    \c0.data_out_1__4_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17086\,
            lcout => \c0.d_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19670\,
            ce => 'H',
            sr => \N__16874\
        );

    \c0.data_out_2__5_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17090\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19670\,
            ce => 'H',
            sr => \N__16874\
        );

    \c0.data_out_1__3_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17085\,
            lcout => \c0.d_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19670\,
            ce => 'H',
            sr => \N__16874\
        );

    \c0.data_out_3__2_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.d_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19670\,
            ce => 'H',
            sr => \N__16874\
        );

    \c0.data_out_2__2_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17089\,
            lcout => \c0.d_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19670\,
            ce => 'H',
            sr => \N__16874\
        );

    \c0.data_out_1__2_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17091\,
            lcout => \c0.d_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19673\,
            ce => 'H',
            sr => \N__16872\
        );

    \c0.byte_transmit_counter_1_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__15632\,
            in1 => \N__15478\,
            in2 => \_gnd_net_\,
            in3 => \N__15337\,
            lcout => \c0.byte_transmit_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19677\,
            ce => \N__15079\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_6_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19677\,
            ce => \N__15079\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_7_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19677\,
            ce => \N__15079\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_3_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19677\,
            ce => \N__15079\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19677\,
            ce => \N__15079\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNIL77O2_1_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__15610\,
            in1 => \N__15429\,
            in2 => \_gnd_net_\,
            in3 => \N__15282\,
            lcout => OPEN,
            ltout => \c0.N_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNI4QES5_2_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100000000"
        )
    port map (
            in0 => \N__15283\,
            in1 => \N__15110\,
            in2 => \N__15082\,
            in3 => \N__15063\,
            lcout => \c0.data_out_0__1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__4_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16011\,
            lcout => \c0.data_in_frame_6_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19629\,
            ce => \N__17170\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_4_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__15802\,
            in1 => \N__18348\,
            in2 => \N__18593\,
            in3 => \N__15796\,
            lcout => \c0.tx2_data_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_4_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__18709\,
            in1 => \N__17941\,
            in2 => \N__18016\,
            in3 => \N__18795\,
            lcout => OPEN,
            ltout => \c0.m120_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_4_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__15790\,
            in1 => \N__15784\,
            in2 => \N__15778\,
            in3 => \N__18711\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19617\,
            ce => \N__19977\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_6_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__18796\,
            in1 => \N__15775\,
            in2 => \N__18073\,
            in3 => \N__18710\,
            lcout => OPEN,
            ltout => \c0.m90_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_6_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__15769\,
            in1 => \N__18718\,
            in2 => \N__15763\,
            in3 => \N__15760\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19617\,
            ce => \N__19977\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_6_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__18592\,
            in1 => \N__17227\,
            in2 => \N__18373\,
            in3 => \N__17197\,
            lcout => \c0.tx2_data_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_6__4_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15754\,
            lcout => \c0.data_in_6_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19630\,
            ce => \N__17726\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__5_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17270\,
            lcout => \c0.data_in_6_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19630\,
            ce => \N__17726\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__5_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15727\,
            lcout => \c0.data_in_7_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19630\,
            ce => \N__17726\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__6_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16080\,
            lcout => \c0.data_in_4_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19630\,
            ce => \N__17726\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__6_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17216\,
            lcout => \c0.data_in_5_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19630\,
            ce => \N__17726\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__6_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17246\,
            lcout => \c0.data_in_6_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19630\,
            ce => \N__17726\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__6_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16069\,
            lcout => \c0.data_in_7_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19630\,
            ce => \N__17726\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIFRNC_10_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15906\,
            in1 => \N__16051\,
            in2 => \N__16010\,
            in3 => \N__15981\,
            lcout => \c0.un1_data_in_6__4_0_a2_5_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__2_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15937\,
            lcout => \c0.d_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19636\,
            ce => \N__17176\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIH6GJ_10_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15905\,
            in1 => \N__16646\,
            in2 => \_gnd_net_\,
            in3 => \N__15819\,
            lcout => \c0.N_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__1_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15877\,
            lcout => \c0.d_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19636\,
            ce => \N__17176\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__1_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15853\,
            lcout => \c0.d_4_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19636\,
            ce => \N__17176\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNISRG61_39_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16647\,
            in1 => \N__18876\,
            in2 => \N__17484\,
            in3 => \N__17745\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__2_0_a2_6_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIK7NH1_24_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16434\,
            in1 => \N__16405\,
            in2 => \N__16384\,
            in3 => \N__18819\,
            lcout => \c0.un1_data_in_6__2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI5G09_46_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17619\,
            in1 => \N__16367\,
            in2 => \N__18004\,
            in3 => \N__16335\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__2_0_a2_0_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI9IAQ1_14_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__16306\,
            in1 => \_gnd_net_\,
            in2 => \N__16285\,
            in3 => \N__16222\,
            lcout => \c0.un1_data_in_7__2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIQ1PT_14_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16273\,
            in1 => \N__16670\,
            in2 => \N__17791\,
            in3 => \N__16246\,
            lcout => \c0.un1_data_in_7__2_0_a2_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI9FFL_29_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16213\,
            in1 => \N__16197\,
            in2 => \_gnd_net_\,
            in3 => \N__17620\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__3_0_a2_0_a2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI6GFI3_15_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000010100"
        )
    port map (
            in0 => \N__16162\,
            in1 => \N__16480\,
            in2 => \N__16141\,
            in3 => \N__16138\,
            lcout => \c0.m163_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__1_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16123\,
            lcout => \c0.d_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19644\,
            ce => \N__17180\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI26S41_15_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16532\,
            in2 => \_gnd_net_\,
            in3 => \N__16515\,
            lcout => \c0.N_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18531\,
            in2 => \N__16474\,
            in3 => \N__16473\,
            lcout => \c0.byte_transmit_counter2Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \c0.un1_byte_transmit_counter2_1_cry_0\,
            clk => \N__19651\,
            ce => 'H',
            sr => \N__19365\
        );

    \c0.byte_transmit_counter2_1_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18764\,
            in2 => \_gnd_net_\,
            in3 => \N__16459\,
            lcout => \c0.byte_transmit_counter2Z0Z_1\,
            ltout => OPEN,
            carryin => \c0.un1_byte_transmit_counter2_1_cry_0\,
            carryout => \c0.un1_byte_transmit_counter2_1_cry_1\,
            clk => \N__19651\,
            ce => 'H',
            sr => \N__19365\
        );

    \c0.byte_transmit_counter2_2_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18708\,
            in2 => \_gnd_net_\,
            in3 => \N__16456\,
            lcout => \c0.byte_transmit_counter2Z0Z_2\,
            ltout => OPEN,
            carryin => \c0.un1_byte_transmit_counter2_1_cry_1\,
            carryout => \c0.un1_byte_transmit_counter2_1_cry_2\,
            clk => \N__19651\,
            ce => 'H',
            sr => \N__19365\
        );

    \c0.byte_transmit_counter2_3_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17863\,
            in2 => \_gnd_net_\,
            in3 => \N__16453\,
            lcout => \c0.byte_transmit_counter2Z0Z_3\,
            ltout => OPEN,
            carryin => \c0.un1_byte_transmit_counter2_1_cry_2\,
            carryout => \c0.un1_byte_transmit_counter2_1_cry_3\,
            clk => \N__19651\,
            ce => 'H',
            sr => \N__19365\
        );

    \c0.byte_transmit_counter2_4_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17824\,
            in2 => \_gnd_net_\,
            in3 => \N__16450\,
            lcout => \c0.byte_transmit_counter2Z0Z_4\,
            ltout => OPEN,
            carryin => \c0.un1_byte_transmit_counter2_1_cry_3\,
            carryout => \c0.un1_byte_transmit_counter2_1_cry_4\,
            clk => \N__19651\,
            ce => 'H',
            sr => \N__19365\
        );

    \c0.byte_transmit_counter2_5_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17839\,
            in2 => \_gnd_net_\,
            in3 => \N__16447\,
            lcout => \c0.byte_transmit_counter2Z0Z_5\,
            ltout => OPEN,
            carryin => \c0.un1_byte_transmit_counter2_1_cry_4\,
            carryout => \c0.un1_byte_transmit_counter2_1_cry_5\,
            clk => \N__19651\,
            ce => 'H',
            sr => \N__19365\
        );

    \c0.byte_transmit_counter2_6_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17851\,
            in2 => \_gnd_net_\,
            in3 => \N__16444\,
            lcout => \c0.byte_transmit_counter2Z0Z_6\,
            ltout => OPEN,
            carryin => \c0.un1_byte_transmit_counter2_1_cry_5\,
            carryout => \c0.un1_byte_transmit_counter2_1_cry_6\,
            clk => \N__19651\,
            ce => 'H',
            sr => \N__19365\
        );

    \c0.byte_transmit_counter2_7_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17875\,
            in2 => \_gnd_net_\,
            in3 => \N__16441\,
            lcout => \c0.byte_transmit_counter2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19651\,
            ce => 'H',
            sr => \N__19365\
        );

    \c0.tx2_data_RNO_3_1_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__16674\,
            in1 => \N__18526\,
            in2 => \N__18333\,
            in3 => \N__16651\,
            lcout => \c0.tx2_data_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_2_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__19818\,
            in1 => \N__17554\,
            in2 => \_gnd_net_\,
            in3 => \N__16624\,
            lcout => \c0.tx2.o_Tx_Serial_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_1_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__18282\,
            in1 => \N__18527\,
            in2 => \N__16615\,
            in3 => \N__17311\,
            lcout => \c0.tx2_data_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__16570\,
            in1 => \N__17103\,
            in2 => \_gnd_net_\,
            in3 => \N__18968\,
            lcout => \c0.tx2.r_Clock_Count_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_5_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__16588\,
            in1 => \N__18601\,
            in2 => \_gnd_net_\,
            in3 => \N__19817\,
            lcout => \c0.tx2.o_Tx_Serial_RNOZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19722\,
            in1 => \N__19353\,
            in2 => \_gnd_net_\,
            in3 => \N__16579\,
            lcout => \c0.tx2_transmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_0_c_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16569\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \c0.tx2.r_Clock_Count12_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16558\,
            in2 => \N__17112\,
            in3 => \N__19001\,
            lcout => \c0.tx2.r_Clock_Count_i_1\,
            ltout => OPEN,
            carryin => \c0.tx2.r_Clock_Count12_cry_0\,
            carryout => \c0.tx2.r_Clock_Count12_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19019\,
            in1 => \N__16552\,
            in2 => \N__17114\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx2.r_Clock_Count_i_2\,
            ltout => OPEN,
            carryin => \c0.tx2.r_Clock_Count12_cry_1\,
            carryout => \c0.tx2.r_Clock_Count12_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17125\,
            in2 => \N__17113\,
            in3 => \N__18983\,
            lcout => \c0.tx2.r_Clock_Count_i_3\,
            ltout => OPEN,
            carryin => \c0.tx2.r_Clock_Count12_cry_2\,
            carryout => \c0.tx2.r_Clock_Count12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17119\,
            lcout => \c0.tx2.r_Clock_Count12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__5_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17093\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19666\,
            ce => 'H',
            sr => \N__16876\
        );

    \c0.tx2.o_Tx_Serial_RNO_6_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__16732\,
            in1 => \N__16720\,
            in2 => \_gnd_net_\,
            in3 => \N__19811\,
            lcout => OPEN,
            ltout => \c0.tx2.o_Tx_Serial_RNOZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_4_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__19741\,
            in1 => \N__19191\,
            in2 => \N__16708\,
            in3 => \N__16705\,
            lcout => OPEN,
            ltout => \c0.tx2.m195_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_1_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__16696\,
            in1 => \N__19193\,
            in2 => \N__16690\,
            in3 => \N__16687\,
            lcout => OPEN,
            ltout => \c0.tx2.N_196_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_0_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19048\,
            in2 => \N__16678\,
            in3 => \N__19138\,
            lcout => \c0.tx2.N_205_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNI7NQN_2_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__19870\,
            in1 => \_gnd_net_\,
            in2 => \N__19141\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx2.N_493\,
            ltout => \c0.tx2.N_493_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011100"
        )
    port map (
            in0 => \N__19249\,
            in1 => \N__19192\,
            in2 => \N__17413\,
            in3 => \N__19764\,
            lcout => \c0.tx2.r_Bit_IndexZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011011100"
        )
    port map (
            in0 => \N__19078\,
            in1 => \N__19946\,
            in2 => \N__19720\,
            in3 => \N__19248\,
            lcout => \c0.tx2_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011110001"
        )
    port map (
            in0 => \N__19222\,
            in1 => \N__19875\,
            in2 => \N__17391\,
            in3 => \N__17410\,
            lcout => \PIN_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19674\,
            ce => 'H',
            sr => \N__19771\
        );

    \c0.data_in_frame_7__0_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17374\,
            lcout => \c0.data_in_frame_7_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19623\,
            ce => \N__17171\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__1_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17341\,
            lcout => \c0.data_in_frame_7_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19623\,
            ce => \N__17171\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__5_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17292\,
            lcout => \c0.data_in_frame_6_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19623\,
            ce => \N__17171\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__5_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17271\,
            lcout => \c0.data_in_frame_7_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19623\,
            ce => \N__17171\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__6_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17247\,
            lcout => \c0.data_in_frame_7_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19623\,
            ce => \N__17171\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__6_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17217\,
            lcout => \c0.data_in_frame_6_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19623\,
            ce => \N__17171\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__2_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17790\,
            lcout => \c0.data_in_6_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19637\,
            ce => \N__17727\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_5_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__18567\,
            in1 => \N__17677\,
            in2 => \N__17656\,
            in3 => \N__18301\,
            lcout => \c0.tx2_data_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_5_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__18569\,
            in1 => \N__17618\,
            in2 => \N__18352\,
            in3 => \N__17590\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_4Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_5_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__18712\,
            in1 => \N__17881\,
            in2 => \N__17566\,
            in3 => \N__18791\,
            lcout => OPEN,
            ltout => \c0.m75_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_5_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__18713\,
            in1 => \N__17563\,
            in2 => \N__17557\,
            in3 => \N__17521\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19645\,
            ce => \N__19969\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_5_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__18304\,
            in1 => \N__17542\,
            in2 => \N__17533\,
            in3 => \N__18568\,
            lcout => \c0.tx2_data_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_7_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__18565\,
            in1 => \N__17515\,
            in2 => \N__17485\,
            in3 => \N__18302\,
            lcout => \c0.tx2_data_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_0_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__18303\,
            in1 => \N__17440\,
            in2 => \N__17425\,
            in3 => \N__18566\,
            lcout => \c0.tx2_data_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_0_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011101111"
        )
    port map (
            in0 => \N__17805\,
            in1 => \N__20012\,
            in2 => \N__19340\,
            in3 => \N__18141\,
            lcout => \c0.N_170_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_6_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__18519\,
            in1 => \N__18124\,
            in2 => \N__18106\,
            in3 => \N__18278\,
            lcout => \c0.tx2_data_RNO_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_4_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__18513\,
            in1 => \N__18061\,
            in2 => \N__18331\,
            in3 => \N__18043\,
            lcout => \c0.tx2_data_RNO_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_4_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__18003\,
            in1 => \N__18518\,
            in2 => \N__18332\,
            in3 => \N__17968\,
            lcout => \c0.tx2_data_RNO_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_5_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__18520\,
            in1 => \N__17929\,
            in2 => \N__17911\,
            in3 => \N__18274\,
            lcout => \c0.tx2_data_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNI8GE8_7_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17874\,
            in2 => \_gnd_net_\,
            in3 => \N__17862\,
            lcout => OPEN,
            ltout => \c0.m45_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNIK84L_4_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__17850\,
            in1 => \N__17838\,
            in2 => \N__17827\,
            in3 => \N__17823\,
            lcout => \c0.N_204_mux\,
            ltout => \c0.N_204_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNIKKP11_1_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__18654\,
            in1 => \N__18762\,
            in2 => \N__17812\,
            in3 => \N__18482\,
            lcout => \c0.N_215_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_0_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__18483\,
            in1 => \N__18901\,
            in2 => \N__18329\,
            in3 => \N__18883\,
            lcout => \c0.tx2_data_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_0_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__18532\,
            in1 => \N__18856\,
            in2 => \N__18829\,
            in3 => \N__18267\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_0_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__18763\,
            in1 => \N__18730\,
            in2 => \N__18724\,
            in3 => \N__18655\,
            lcout => OPEN,
            ltout => \c0.m146_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_0_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__18656\,
            in1 => \N__18613\,
            in2 => \N__18604\,
            in3 => \N__18157\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19659\,
            ce => \N__19968\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_0_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__18484\,
            in1 => \N__18406\,
            in2 => \N__18330\,
            in3 => \N__18181\,
            lcout => \c0.tx2_data_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_0_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18947\,
            in1 => \N__18970\,
            in2 => \N__18933\,
            in3 => \N__18934\,
            lcout => \c0.tx2.r_Clock_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \c0.tx2.un1_r_Clock_Count_cry_0\,
            clk => \N__19667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_1_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__18954\,
            in1 => \_gnd_net_\,
            in2 => \N__19006\,
            in3 => \N__18151\,
            lcout => \c0.tx2.r_Clock_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \c0.tx2.un1_r_Clock_Count_cry_0\,
            carryout => \c0.tx2.un1_r_Clock_Count_cry_1\,
            clk => \N__19667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_2_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__18948\,
            in1 => \_gnd_net_\,
            in2 => \N__19024\,
            in3 => \N__18148\,
            lcout => \c0.tx2.r_Clock_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \c0.tx2.un1_r_Clock_Count_cry_1\,
            carryout => \c0.tx2.un1_r_Clock_Count_cry_2\,
            clk => \N__19667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_3_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18955\,
            in1 => \N__18987\,
            in2 => \_gnd_net_\,
            in3 => \N__18145\,
            lcout => \c0.tx2.r_Clock_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_RNIE5AU_3_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19020\,
            in1 => \N__19002\,
            in2 => \N__18988\,
            in3 => \N__18969\,
            lcout => \c0.tx2.N_171_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNI9USD1_4_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__19246\,
            in1 => \N__19221\,
            in2 => \N__19912\,
            in3 => \N__19857\,
            lcout => \c0.tx2.N_16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNI9USD1_0_4_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19856\,
            in1 => \N__19219\,
            in2 => \N__19915\,
            in3 => \N__19245\,
            lcout => \c0.tx2.r_Clock_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_0_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110010"
        )
    port map (
            in0 => \N__19220\,
            in1 => \N__19134\,
            in2 => \N__19258\,
            in3 => \N__19858\,
            lcout => \c0.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.N_90_ip_RNO_0_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19133\,
            in1 => \N__19164\,
            in2 => \_gnd_net_\,
            in3 => \N__19899\,
            lcout => OPEN,
            ltout => \c0.tx2.N_83_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.N_90_ip_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111111"
        )
    port map (
            in0 => \N__19218\,
            in1 => \N__19045\,
            in2 => \N__18916\,
            in3 => \N__18907\,
            lcout => \c0.N_90_dup\,
            ltout => \c0.N_90_dup_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNO_0_1_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19105\,
            in2 => \N__18913\,
            in3 => \N__19903\,
            lcout => OPEN,
            ltout => \c0.tx2.i97_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_1_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__19166\,
            in1 => \N__19952\,
            in2 => \N__18910\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx2.r_SM_Main_dup_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.N_90_ip_RNO_1_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__19132\,
            in1 => \N__19165\,
            in2 => \_gnd_net_\,
            in3 => \N__19898\,
            lcout => \c0.tx2.r_SM_Main_illegal_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNO_0_0_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19047\,
            in1 => \N__20011\,
            in2 => \_gnd_net_\,
            in3 => \N__19167\,
            lcout => \c0.tx2.N_214_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_RNIPHKF1_0_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__19861\,
            in1 => \N__19139\,
            in2 => \N__19198\,
            in3 => \N__19247\,
            lcout => \c0.tx2.N_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNI8OQN_3_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19046\,
            in2 => \_gnd_net_\,
            in3 => \N__19859\,
            lcout => \c0.tx2.N_17_0\,
            ltout => \c0.tx2.N_17_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_4_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19225\,
            in3 => \N__19106\,
            lcout => \c0.tx2.r_SM_Main_dup_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_RNIN3O01_1_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19747\,
            in1 => \N__19194\,
            in2 => \_gnd_net_\,
            in3 => \N__19815\,
            lcout => \c0.tx2.N_212_0\,
            ltout => \c0.tx2.N_212_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNO_0_2_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000100"
        )
    port map (
            in0 => \N__19860\,
            in1 => \N__19140\,
            in2 => \N__19171\,
            in3 => \N__19168\,
            lcout => OPEN,
            ltout => \c0.tx2.N_496_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_2_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__19056\,
            in1 => \_gnd_net_\,
            in2 => \N__19144\,
            in3 => \N__19107\,
            lcout => \c0.tx2.r_SM_Main_dup_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_3_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19108\,
            in1 => \N__19077\,
            in2 => \N__19066\,
            in3 => \N__19057\,
            lcout => \c0.tx2.r_SM_Main_dup_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_RNILRI51_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19913\,
            in2 => \N__19876\,
            in3 => \N__20014\,
            lcout => \c0.N_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNI5LQN_0_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__19914\,
            in1 => \N__19871\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx2.N_9_1\,
            ltout => \c0.tx2.N_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_2_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__19746\,
            in1 => \N__19780\,
            in2 => \N__19825\,
            in3 => \N__19816\,
            lcout => \c0.tx2.r_Bit_IndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_1_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__19745\,
            in1 => \N__19779\,
            in2 => \_gnd_net_\,
            in3 => \N__19763\,
            lcout => \c0.tx2.r_Bit_IndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__19723\,
            in1 => \N__19326\,
            in2 => \_gnd_net_\,
            in3 => \N__19684\,
            lcout => \c0.wait_for_transmissionZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19660\,
            ce => 'H',
            sr => \N__19369\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19341\,
            in2 => \_gnd_net_\,
            in3 => \N__19291\,
            lcout => \c0.data_in_frame_0__0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
