-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 12 2019 19:18:20

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : inout std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : inout std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : inout std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__52613\ : std_logic;
signal \N__52612\ : std_logic;
signal \N__52611\ : std_logic;
signal \N__52604\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52595\ : std_logic;
signal \N__52594\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52585\ : std_logic;
signal \N__52584\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52576\ : std_logic;
signal \N__52575\ : std_logic;
signal \N__52568\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52566\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52548\ : std_logic;
signal \N__52545\ : std_logic;
signal \N__52544\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52527\ : std_logic;
signal \N__52524\ : std_logic;
signal \N__52521\ : std_logic;
signal \N__52518\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52511\ : std_logic;
signal \N__52508\ : std_logic;
signal \N__52505\ : std_logic;
signal \N__52502\ : std_logic;
signal \N__52499\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52494\ : std_logic;
signal \N__52491\ : std_logic;
signal \N__52488\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52480\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52464\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52461\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52458\ : std_logic;
signal \N__52457\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52455\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52453\ : std_logic;
signal \N__52452\ : std_logic;
signal \N__52451\ : std_logic;
signal \N__52448\ : std_logic;
signal \N__52445\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52415\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52409\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52406\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52396\ : std_logic;
signal \N__52393\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52374\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52361\ : std_logic;
signal \N__52358\ : std_logic;
signal \N__52355\ : std_logic;
signal \N__52352\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52335\ : std_logic;
signal \N__52322\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52306\ : std_logic;
signal \N__52303\ : std_logic;
signal \N__52302\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52300\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52296\ : std_logic;
signal \N__52295\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52290\ : std_logic;
signal \N__52289\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52261\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52251\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52231\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52227\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52202\ : std_logic;
signal \N__52197\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52187\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52175\ : std_logic;
signal \N__52172\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52141\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52137\ : std_logic;
signal \N__52136\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52131\ : std_logic;
signal \N__52128\ : std_logic;
signal \N__52125\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52116\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52098\ : std_logic;
signal \N__52097\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52089\ : std_logic;
signal \N__52088\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52085\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52082\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52080\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52076\ : std_logic;
signal \N__52073\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52071\ : std_logic;
signal \N__52070\ : std_logic;
signal \N__52067\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52065\ : std_logic;
signal \N__52064\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52062\ : std_logic;
signal \N__52061\ : std_logic;
signal \N__52060\ : std_logic;
signal \N__52057\ : std_logic;
signal \N__52056\ : std_logic;
signal \N__52055\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52045\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52043\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52040\ : std_logic;
signal \N__52039\ : std_logic;
signal \N__52038\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52025\ : std_logic;
signal \N__52022\ : std_logic;
signal \N__52019\ : std_logic;
signal \N__52016\ : std_logic;
signal \N__52013\ : std_logic;
signal \N__52010\ : std_logic;
signal \N__52005\ : std_logic;
signal \N__51998\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51995\ : std_logic;
signal \N__51994\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51990\ : std_logic;
signal \N__51987\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51976\ : std_logic;
signal \N__51973\ : std_logic;
signal \N__51972\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51970\ : std_logic;
signal \N__51967\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51957\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51938\ : std_logic;
signal \N__51935\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51913\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51898\ : std_logic;
signal \N__51893\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51864\ : std_logic;
signal \N__51857\ : std_logic;
signal \N__51854\ : std_logic;
signal \N__51851\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51829\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51812\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51774\ : std_logic;
signal \N__51771\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51767\ : std_logic;
signal \N__51764\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51761\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51752\ : std_logic;
signal \N__51749\ : std_logic;
signal \N__51746\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51739\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51733\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51718\ : std_logic;
signal \N__51715\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51702\ : std_logic;
signal \N__51701\ : std_logic;
signal \N__51698\ : std_logic;
signal \N__51695\ : std_logic;
signal \N__51692\ : std_logic;
signal \N__51689\ : std_logic;
signal \N__51686\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51667\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51655\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51651\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51647\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51644\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51634\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51632\ : std_logic;
signal \N__51631\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51621\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51618\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51616\ : std_logic;
signal \N__51615\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51613\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51609\ : std_logic;
signal \N__51608\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51586\ : std_logic;
signal \N__51583\ : std_logic;
signal \N__51580\ : std_logic;
signal \N__51577\ : std_logic;
signal \N__51576\ : std_logic;
signal \N__51571\ : std_logic;
signal \N__51564\ : std_logic;
signal \N__51561\ : std_logic;
signal \N__51558\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51545\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51532\ : std_logic;
signal \N__51525\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51512\ : std_logic;
signal \N__51509\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51463\ : std_logic;
signal \N__51462\ : std_logic;
signal \N__51459\ : std_logic;
signal \N__51456\ : std_logic;
signal \N__51453\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51447\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51423\ : std_logic;
signal \N__51420\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51411\ : std_logic;
signal \N__51408\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51404\ : std_logic;
signal \N__51401\ : std_logic;
signal \N__51398\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51384\ : std_logic;
signal \N__51381\ : std_logic;
signal \N__51378\ : std_logic;
signal \N__51373\ : std_logic;
signal \N__51370\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51340\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51338\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51327\ : std_logic;
signal \N__51322\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51313\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51305\ : std_logic;
signal \N__51304\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51295\ : std_logic;
signal \N__51292\ : std_logic;
signal \N__51289\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51279\ : std_logic;
signal \N__51278\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51275\ : std_logic;
signal \N__51274\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51271\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51250\ : std_logic;
signal \N__51249\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51246\ : std_logic;
signal \N__51245\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51243\ : std_logic;
signal \N__51240\ : std_logic;
signal \N__51237\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51225\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51222\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51219\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51215\ : std_logic;
signal \N__51214\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51209\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51206\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51202\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51199\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51196\ : std_logic;
signal \N__51195\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51193\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51187\ : std_logic;
signal \N__51186\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51184\ : std_logic;
signal \N__51183\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51180\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51177\ : std_logic;
signal \N__51174\ : std_logic;
signal \N__51171\ : std_logic;
signal \N__51170\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51162\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51154\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51147\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51138\ : std_logic;
signal \N__51137\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51135\ : std_logic;
signal \N__51132\ : std_logic;
signal \N__51131\ : std_logic;
signal \N__51130\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51117\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51109\ : std_logic;
signal \N__51106\ : std_logic;
signal \N__51105\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51103\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51089\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51073\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51061\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51018\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51005\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__51001\ : std_logic;
signal \N__50996\ : std_logic;
signal \N__50995\ : std_logic;
signal \N__50992\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50974\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50965\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50951\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50948\ : std_logic;
signal \N__50947\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50942\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50939\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50936\ : std_logic;
signal \N__50935\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50929\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50926\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50923\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50863\ : std_logic;
signal \N__50854\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50812\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50737\ : std_logic;
signal \N__50728\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50644\ : std_logic;
signal \N__50641\ : std_logic;
signal \N__50638\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50636\ : std_logic;
signal \N__50635\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50628\ : std_logic;
signal \N__50623\ : std_logic;
signal \N__50620\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50614\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50591\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50579\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50576\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50569\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50566\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50564\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50531\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50519\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50503\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50475\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50451\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49673\ : std_logic;
signal \N__49670\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49595\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49300\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__49290\ : std_logic;
signal \N__49287\ : std_logic;
signal \N__49284\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49029\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48906\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48630\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47023\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43036\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41392\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36436\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n17299_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal tx2_enable : std_logic;
signal n17298 : std_logic;
signal \bfn_1_28_0_\ : std_logic;
signal \c0.tx2.n15675\ : std_logic;
signal \c0.tx2.n15676\ : std_logic;
signal n17457 : std_logic;
signal \c0.tx2.n15677\ : std_logic;
signal \c0.tx2.n15678\ : std_logic;
signal \c0.tx2.n15679\ : std_logic;
signal \c0.tx2.n15680\ : std_logic;
signal \c0.tx2.n15681\ : std_logic;
signal \c0.tx2.n15682\ : std_logic;
signal \bfn_1_29_0_\ : std_logic;
signal n17640 : std_logic;
signal n16824 : std_logic;
signal n10_adj_2412 : std_logic;
signal n17458 : std_logic;
signal \bfn_1_30_0_\ : std_logic;
signal \c0.tx.n15660\ : std_logic;
signal \c0.tx.n15661\ : std_logic;
signal \c0.tx.n15662\ : std_logic;
signal \c0.tx.n15663\ : std_logic;
signal \c0.tx.n15664\ : std_logic;
signal \c0.tx.n15665\ : std_logic;
signal \c0.tx.n15666\ : std_logic;
signal \c0.tx.n15667\ : std_logic;
signal \bfn_1_31_0_\ : std_logic;
signal \n17537_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2090_2_cascade_\ : std_logic;
signal n17631 : std_logic;
signal \n16810_cascade_\ : std_logic;
signal \c0.rx.n13452_cascade_\ : std_logic;
signal n16867 : std_logic;
signal n17222 : std_logic;
signal \c0.rx.n16850\ : std_logic;
signal \c0.FRAME_MATCHER_state_7\ : std_logic;
signal \c0.n16443\ : std_logic;
signal \c0.FRAME_MATCHER_state_13\ : std_logic;
signal \c0.n16447\ : std_logic;
signal \c0.FRAME_MATCHER_state_11\ : std_logic;
signal \c0.n16451\ : std_logic;
signal \c0.n16445\ : std_logic;
signal n26 : std_logic;
signal \bfn_2_25_0_\ : std_logic;
signal n25 : std_logic;
signal n15590 : std_logic;
signal n24 : std_logic;
signal n15591 : std_logic;
signal n23 : std_logic;
signal n15592 : std_logic;
signal n22 : std_logic;
signal n15593 : std_logic;
signal n21 : std_logic;
signal n15594 : std_logic;
signal n20 : std_logic;
signal n15595 : std_logic;
signal n19 : std_logic;
signal n15596 : std_logic;
signal n15597 : std_logic;
signal n18 : std_logic;
signal \bfn_2_26_0_\ : std_logic;
signal n17_adj_2422 : std_logic;
signal n15598 : std_logic;
signal n16 : std_logic;
signal n15599 : std_logic;
signal n15 : std_logic;
signal n15600 : std_logic;
signal n14_adj_2424 : std_logic;
signal n15601 : std_logic;
signal n13 : std_logic;
signal n15602 : std_logic;
signal n12_adj_2419 : std_logic;
signal n15603 : std_logic;
signal n11 : std_logic;
signal n15604 : std_logic;
signal n15605 : std_logic;
signal n10_adj_2420 : std_logic;
signal \bfn_2_27_0_\ : std_logic;
signal n9 : std_logic;
signal n15606 : std_logic;
signal n8 : std_logic;
signal n15607 : std_logic;
signal n7 : std_logic;
signal n15608 : std_logic;
signal n6_adj_2421 : std_logic;
signal n15609 : std_logic;
signal blink_counter_21 : std_logic;
signal n15610 : std_logic;
signal blink_counter_22 : std_logic;
signal n15611 : std_logic;
signal blink_counter_23 : std_logic;
signal n15612 : std_logic;
signal n15613 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_2_28_0_\ : std_logic;
signal n15614 : std_logic;
signal blink_counter_25 : std_logic;
signal n17570 : std_logic;
signal n17629 : std_logic;
signal n17504 : std_logic;
signal \r_Clock_Count_2_adj_2452\ : std_logic;
signal \r_Clock_Count_3_adj_2451\ : std_logic;
signal n9403 : std_logic;
signal \n17140_cascade_\ : std_logic;
signal n16817 : std_logic;
signal n12_adj_2410 : std_logic;
signal \r_Clock_Count_5_adj_2449\ : std_logic;
signal \r_Clock_Count_1_adj_2453\ : std_logic;
signal \c0.tx2.n10\ : std_logic;
signal n15837 : std_logic;
signal \n15837_cascade_\ : std_logic;
signal \r_SM_Main_2_N_2033_1_cascade_\ : std_logic;
signal \r_Clock_Count_7_adj_2447\ : std_logic;
signal \r_Clock_Count_8_adj_2446\ : std_logic;
signal n9929 : std_logic;
signal n17494 : std_logic;
signal n17542 : std_logic;
signal n17484 : std_logic;
signal \n17_adj_2416_cascade_\ : std_logic;
signal \r_Clock_Count_2\ : std_logic;
signal \r_Clock_Count_3\ : std_logic;
signal \r_Clock_Count_0\ : std_logic;
signal \r_Clock_Count_5\ : std_logic;
signal \c0.tx.n10_cascade_\ : std_logic;
signal n16863 : std_logic;
signal \n16863_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2096_0_cascade_\ : std_logic;
signal n6_adj_2461 : std_logic;
signal n17641 : std_logic;
signal \n17144_cascade_\ : std_logic;
signal n16828 : std_logic;
signal \bfn_2_32_0_\ : std_logic;
signal \c0.rx.n15668\ : std_logic;
signal \r_Clock_Count_2_adj_2435\ : std_logic;
signal n16860 : std_logic;
signal \c0.rx.n15669\ : std_logic;
signal \c0.rx.n15670\ : std_logic;
signal n16854 : std_logic;
signal \c0.rx.n15671\ : std_logic;
signal \c0.rx.n15672\ : std_logic;
signal \c0.rx.n15673\ : std_logic;
signal \r_Clock_Count_7_adj_2430\ : std_logic;
signal n16852 : std_logic;
signal \c0.rx.n15674\ : std_logic;
signal n16855 : std_logic;
signal \c0.FRAME_MATCHER_state_15\ : std_logic;
signal \c0.n16349\ : std_logic;
signal \n1651_cascade_\ : std_logic;
signal n1651 : std_logic;
signal \n6_cascade_\ : std_logic;
signal n4 : std_logic;
signal \n8_adj_2459_cascade_\ : std_logic;
signal \FRAME_MATCHER_state_31_N_1440_1\ : std_logic;
signal n3_adj_2408 : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_5_cascade_\ : std_logic;
signal \c0.n3_adj_2256\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_4_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_3_cascade_\ : std_logic;
signal \c0.n3_adj_2258\ : std_logic;
signal \c0.n16379\ : std_logic;
signal \c0.n3_adj_2242\ : std_logic;
signal \c0.n3_adj_2243\ : std_logic;
signal \c0.n3_adj_2244\ : std_logic;
signal \c0.n17172_cascade_\ : std_logic;
signal data_in_0_7 : std_logic;
signal data_in_1_5 : std_logic;
signal data_in_0_4 : std_logic;
signal \n9472_cascade_\ : std_logic;
signal \c0.rx.n10086_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2090_2\ : std_logic;
signal \n14060_cascade_\ : std_logic;
signal \n7866_cascade_\ : std_logic;
signal \n10425_cascade_\ : std_logic;
signal n12 : std_logic;
signal n13276 : std_logic;
signal \n10_adj_2415_cascade_\ : std_logic;
signal n15701 : std_logic;
signal n16844 : std_logic;
signal n17461 : std_logic;
signal \r_Clock_Count_1\ : std_logic;
signal n17601 : std_logic;
signal n17602 : std_logic;
signal \r_Clock_Count_4_adj_2433\ : std_logic;
signal \c0.rx.n6\ : std_logic;
signal n16853 : std_logic;
signal \r_Clock_Count_1_adj_2436\ : std_logic;
signal n4_adj_2411 : std_logic;
signal n17260 : std_logic;
signal n10425 : std_logic;
signal n16857 : std_logic;
signal \r_Clock_Count_5_adj_2432\ : std_logic;
signal n16858 : std_logic;
signal \r_Clock_Count_3_adj_2434\ : std_logic;
signal n9406 : std_logic;
signal \c0.n3_adj_2217\ : std_logic;
signal \c0.n3_adj_2215\ : std_logic;
signal \c0.n3_adj_2210\ : std_logic;
signal \c0.n3_adj_2249\ : std_logic;
signal \c0.n9393\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_2_cascade_\ : std_logic;
signal \c0.n3_adj_2259\ : std_logic;
signal \c0.n10_adj_2329\ : std_logic;
signal \c0.n16895\ : std_logic;
signal \c0.n16895_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_1_cascade_\ : std_logic;
signal \c0.n3_adj_2260\ : std_logic;
signal \bfn_4_22_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_1\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_1\ : std_logic;
signal \c0.n15622\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_2\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_2\ : std_logic;
signal \c0.n15623\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_3\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_3\ : std_logic;
signal \c0.n15624\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_4\ : std_logic;
signal \c0.n15625\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_5\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_5\ : std_logic;
signal \c0.n15626\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_6\ : std_logic;
signal \c0.n15627\ : std_logic;
signal \c0.n15628\ : std_logic;
signal \c0.n15629\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_8\ : std_logic;
signal \bfn_4_23_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_9\ : std_logic;
signal \c0.n15630\ : std_logic;
signal \c0.n15631\ : std_logic;
signal \c0.n15632\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_12\ : std_logic;
signal \c0.n15633\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_13\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_13\ : std_logic;
signal \c0.n15634\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_14\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_14\ : std_logic;
signal \c0.n15635\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_15\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_15\ : std_logic;
signal \c0.n15636\ : std_logic;
signal \c0.n15637\ : std_logic;
signal \bfn_4_24_0_\ : std_logic;
signal \c0.n15638\ : std_logic;
signal \c0.n15639\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_19\ : std_logic;
signal \c0.n15640\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_20\ : std_logic;
signal \c0.n15641\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_21\ : std_logic;
signal \c0.n15642\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_22\ : std_logic;
signal \c0.n15643\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_23\ : std_logic;
signal \c0.n15644\ : std_logic;
signal \c0.n15645\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_24\ : std_logic;
signal \bfn_4_25_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_25\ : std_logic;
signal \c0.n15646\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_26\ : std_logic;
signal \c0.n15647\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_27\ : std_logic;
signal \c0.n15648\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_28\ : std_logic;
signal \c0.n15649\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_29\ : std_logic;
signal \c0.n15650\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_30\ : std_logic;
signal \c0.n15651\ : std_logic;
signal \c0.n15652\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_31\ : std_logic;
signal data_in_0_6 : std_logic;
signal \c0.n17274_cascade_\ : std_logic;
signal \c0.n17889\ : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_2_1 : std_logic;
signal data_in_2_4 : std_logic;
signal data_in_1_4 : std_logic;
signal n17567 : std_logic;
signal \r_Clock_Count_4_adj_2450\ : std_logic;
signal data_in_2_3 : std_logic;
signal n16856 : std_logic;
signal \r_Clock_Count_6_adj_2431\ : std_logic;
signal \n16893_cascade_\ : std_logic;
signal n5 : std_logic;
signal n17636 : std_logic;
signal \r_SM_Main_2_N_2033_1\ : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \r_Bit_Index_1_adj_2438\ : std_logic;
signal \r_Clock_Count_7\ : std_logic;
signal \r_Clock_Count_6\ : std_logic;
signal \r_Clock_Count_8\ : std_logic;
signal n9937 : std_logic;
signal \c0.tx.n15683_cascade_\ : std_logic;
signal \c0.tx.n14082\ : std_logic;
signal n17573 : std_logic;
signal \r_Clock_Count_4\ : std_logic;
signal \c0.n12993_cascade_\ : std_logic;
signal \c0.n12993\ : std_logic;
signal \c0.n13298\ : std_logic;
signal \c0.n20_adj_2267\ : std_logic;
signal \c0.n21_adj_2271_cascade_\ : std_logic;
signal \n29_cascade_\ : std_logic;
signal tx_enable : std_logic;
signal \c0.n12991\ : std_logic;
signal \c0.n12991_cascade_\ : std_logic;
signal \c0.n19_adj_2270\ : std_logic;
signal n16859 : std_logic;
signal n17_adj_2416 : std_logic;
signal \r_Clock_Count_0_adj_2437\ : std_logic;
signal tx_o : std_logic;
signal data_in_1_0 : std_logic;
signal \n3977_cascade_\ : std_logic;
signal \c0.n3_adj_2233\ : std_logic;
signal \c0.n3_adj_2219\ : std_logic;
signal \c0.n16441\ : std_logic;
signal \c0.n3_adj_2229\ : std_logic;
signal \c0.n3_adj_2231\ : std_logic;
signal \c0.n3_adj_2227\ : std_logic;
signal \c0.n3_adj_2223\ : std_logic;
signal \c0.n3_adj_2225\ : std_logic;
signal \c0.n1439_cascade_\ : std_logic;
signal \c0.n3_adj_2221\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_7\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_7\ : std_logic;
signal \c0.n3_adj_2250\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_6\ : std_logic;
signal \c0.n3_adj_2253\ : std_logic;
signal \c0.n3_adj_2237\ : std_logic;
signal \c0.n3_adj_2235\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_11\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_11\ : std_logic;
signal \c0.n3_adj_2246\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_10\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_9\ : std_logic;
signal \c0.n3_adj_2248\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_8\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_19\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_20\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_21\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_23\ : std_logic;
signal \c0.n18_adj_2198_cascade_\ : std_logic;
signal \c0.n127_adj_2136_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_27\ : std_logic;
signal n9472 : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_30\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_25\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_28\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_24\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_26\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_22\ : std_logic;
signal \c0.n12_adj_2200\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_31\ : std_logic;
signal n4_adj_2460 : std_logic;
signal n4_adj_2417 : std_logic;
signal data_in_0_2 : std_logic;
signal data_in_1_3 : std_logic;
signal n13082 : std_logic;
signal \c0.n16891_cascade_\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \c0.rx.n9323\ : std_logic;
signal n9477 : std_logic;
signal n4_adj_2409 : std_logic;
signal \n9477_cascade_\ : std_logic;
signal n16893 : std_logic;
signal \c0.tx.n17462\ : std_logic;
signal \c0.tx.r_Bit_Index_0\ : std_logic;
signal n17397 : std_logic;
signal \c0.tx.r_Bit_Index_2\ : std_logic;
signal \c0.tx.n17975_cascade_\ : std_logic;
signal \c0.tx.o_Tx_Serial_N_2064_cascade_\ : std_logic;
signal n3_adj_2406 : std_logic;
signal \c0.n1419_cascade_\ : std_logic;
signal \c0.n1419\ : std_logic;
signal n53 : std_logic;
signal \c0.delay_counter_0\ : std_logic;
signal \c0.n17637\ : std_logic;
signal \bfn_5_31_0_\ : std_logic;
signal \c0.delay_counter_1\ : std_logic;
signal \c0.n6531\ : std_logic;
signal \c0.n15514\ : std_logic;
signal \c0.n6530\ : std_logic;
signal \c0.n15515\ : std_logic;
signal \c0.delay_counter_3\ : std_logic;
signal \c0.n6529\ : std_logic;
signal \c0.n15516\ : std_logic;
signal \c0.n6528\ : std_logic;
signal \c0.n15517\ : std_logic;
signal \c0.delay_counter_5\ : std_logic;
signal \c0.n17574\ : std_logic;
signal \c0.n15518\ : std_logic;
signal \c0.delay_counter_6\ : std_logic;
signal \c0.n6526\ : std_logic;
signal \c0.n15519\ : std_logic;
signal \c0.delay_counter_7\ : std_logic;
signal \c0.n17638\ : std_logic;
signal \c0.n15520\ : std_logic;
signal \c0.n15521\ : std_logic;
signal \c0.n6524\ : std_logic;
signal \bfn_5_32_0_\ : std_logic;
signal \c0.delay_counter_9\ : std_logic;
signal \c0.n6523\ : std_logic;
signal \c0.n15522\ : std_logic;
signal \c0.delay_counter_10\ : std_logic;
signal \c0.n6522\ : std_logic;
signal \c0.n15523\ : std_logic;
signal \c0.delay_counter_11\ : std_logic;
signal \c0.n6521\ : std_logic;
signal \c0.n15524\ : std_logic;
signal \c0.delay_counter_12\ : std_logic;
signal \c0.n17575\ : std_logic;
signal \c0.n15525\ : std_logic;
signal \c0.n17639\ : std_logic;
signal \c0.n15526\ : std_logic;
signal \c0.delay_counter_14\ : std_logic;
signal \c0.n15527\ : std_logic;
signal \c0.n17635\ : std_logic;
signal \c0.n16331\ : std_logic;
signal \c0.n16381\ : std_logic;
signal \c0.FRAME_MATCHER_i_19\ : std_logic;
signal \c0.FRAME_MATCHER_i_24\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_16\ : std_logic;
signal \n1716_cascade_\ : std_logic;
signal n14 : std_logic;
signal n16775 : std_logic;
signal n3977 : std_logic;
signal \n16775_cascade_\ : std_logic;
signal n9453 : std_logic;
signal \c0.FRAME_MATCHER_i_1\ : std_logic;
signal n2275 : std_logic;
signal \n2275_cascade_\ : std_logic;
signal \c0.n7212_cascade_\ : std_logic;
signal \c0.n17452_cascade_\ : std_logic;
signal \c0.n17454\ : std_logic;
signal \c0.n7_cascade_\ : std_logic;
signal \c0.n16335\ : std_logic;
signal \c0.FRAME_MATCHER_state_5\ : std_logic;
signal \c0.FRAME_MATCHER_state_6\ : std_logic;
signal \c0.FRAME_MATCHER_state_29\ : std_logic;
signal \c0.n59_cascade_\ : std_logic;
signal \c0.n5_adj_2262_cascade_\ : std_logic;
signal \c0.n16876_cascade_\ : std_logic;
signal \c0.n60_cascade_\ : std_logic;
signal \c0.n16363\ : std_logic;
signal \c0.FRAME_MATCHER_state_30\ : std_logic;
signal \c0.FRAME_MATCHER_state_23\ : std_logic;
signal \c0.n9451_cascade_\ : std_logic;
signal \n12933_cascade_\ : std_logic;
signal \c0.n9451\ : std_logic;
signal \c0.n9\ : std_logic;
signal \c0.n17258\ : std_logic;
signal \c0.n28_cascade_\ : std_logic;
signal \c0.n60\ : std_logic;
signal \c0.n16879\ : std_logic;
signal \c0.n33\ : std_logic;
signal \c0.n16879_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_6\ : std_logic;
signal \c0.FRAME_MATCHER_i_7\ : std_logic;
signal \c0.FRAME_MATCHER_i_9\ : std_logic;
signal n9445 : std_logic;
signal \c0.n9488\ : std_logic;
signal \c0.n12_adj_2158\ : std_logic;
signal \c0.n9488_cascade_\ : std_logic;
signal \c0.n17262\ : std_logic;
signal \c0.n17256\ : std_logic;
signal data_in_0_0 : std_logic;
signal \c0.n9485\ : std_logic;
signal \c0.n10_adj_2149_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_29\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_29\ : std_logic;
signal data_in_3_0 : std_logic;
signal data_in_0_5 : std_logic;
signal data_in_3_4 : std_logic;
signal \c0.n17264\ : std_logic;
signal \c0.n9493\ : std_logic;
signal \c0.n12_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31\ : std_logic;
signal \n127_adj_2418_cascade_\ : std_logic;
signal \c0.n17240\ : std_logic;
signal data_in_1_1 : std_logic;
signal \c0.n9482\ : std_logic;
signal \c0.n9490\ : std_logic;
signal n16795 : std_logic;
signal \n127_cascade_\ : std_logic;
signal \c0.n2\ : std_logic;
signal \c0.n2_cascade_\ : std_logic;
signal n9435 : std_logic;
signal n7198 : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_18\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_18\ : std_logic;
signal \c0.FRAME_MATCHER_i_18\ : std_logic;
signal \c0.n3_adj_2239\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_17\ : std_logic;
signal \c0.n127_adj_2136\ : std_logic;
signal n127 : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_16\ : std_logic;
signal n127_adj_2418 : std_logic;
signal \c0.FRAME_MATCHER_i_16\ : std_logic;
signal \c0.n7212\ : std_logic;
signal \c0.n3_adj_2241\ : std_logic;
signal \c0.data_in_frame_9_2\ : std_logic;
signal \c0.n15939\ : std_logic;
signal \c0.data_in_frame_10_0\ : std_logic;
signal \c0.n17013_cascade_\ : std_logic;
signal \c0.n17013\ : std_logic;
signal \c0.data_in_frame_9_7\ : std_logic;
signal data_in_3_6 : std_logic;
signal data_in_2_0 : std_logic;
signal \c0.n17268\ : std_logic;
signal data_in_1_7 : std_logic;
signal data_in_0_3 : std_logic;
signal \c0.n19_adj_2199\ : std_logic;
signal \c0.data_in_frame_10_1\ : std_logic;
signal \c0.n9743\ : std_logic;
signal \c0.n16954_cascade_\ : std_logic;
signal \c0.data_in_frame_10_6\ : std_logic;
signal \c0.n18_adj_2174_cascade_\ : std_logic;
signal \c0.n17015\ : std_logic;
signal \c0.data_in_frame_9_4\ : std_logic;
signal \c0.n6_adj_2152\ : std_logic;
signal \c0.n13272\ : std_logic;
signal \c0.n16882_cascade_\ : std_logic;
signal \c0.data_in_frame_10_4\ : std_logic;
signal \c0.data_in_frame_9_6\ : std_logic;
signal \c0.data_in_frame_2_7\ : std_logic;
signal \c0.n25_adj_2324\ : std_logic;
signal \n4_adj_2458_cascade_\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal n14060 : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal n17395 : std_logic;
signal \c0.tx_active_prev\ : std_logic;
signal \c0.n65\ : std_logic;
signal \bfn_6_30_0_\ : std_logic;
signal \c0.n15653\ : std_logic;
signal \c0.n15654\ : std_logic;
signal \c0.n15655\ : std_logic;
signal \c0.n15656\ : std_logic;
signal \c0.n15657\ : std_logic;
signal \c0.n15658\ : std_logic;
signal \c0.n15659\ : std_logic;
signal \c0.n8938_cascade_\ : std_logic;
signal \c0.n22_adj_2164\ : std_logic;
signal \c0.n22_adj_2164_cascade_\ : std_logic;
signal \c0.tx_transmit_N_1949_1\ : std_logic;
signal \c0.n15868_cascade_\ : std_logic;
signal \c0.n8631\ : std_logic;
signal \n10141_cascade_\ : std_logic;
signal \c0.n446\ : std_logic;
signal \c0.n446_cascade_\ : std_logic;
signal \c0.n456\ : std_logic;
signal \c0.n16371\ : std_logic;
signal \c0.n16453\ : std_logic;
signal \c0.n59\ : std_logic;
signal \c0.n61_cascade_\ : std_logic;
signal \c0.n10_adj_2336\ : std_logic;
signal \c0.n16133_cascade_\ : std_logic;
signal \c0.n16898\ : std_logic;
signal \c0.FRAME_MATCHER_state_19\ : std_logic;
signal \c0.n52\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_4\ : std_logic;
signal \c0.n3_adj_2257\ : std_logic;
signal \c0.FRAME_MATCHER_i_20\ : std_logic;
signal \c0.FRAME_MATCHER_i_4\ : std_logic;
signal \c0.FRAME_MATCHER_i_5\ : std_logic;
signal \c0.FRAME_MATCHER_i_21\ : std_logic;
signal \c0.n30_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_13\ : std_logic;
signal \c0.n56\ : std_logic;
signal \c0.FRAME_MATCHER_state_10\ : std_logic;
signal \c0.n6_adj_2213\ : std_logic;
signal \c0.n16869\ : std_logic;
signal \c0.n16869_cascade_\ : std_logic;
signal \c0.n16871_cascade_\ : std_logic;
signal \c0.n16876\ : std_logic;
signal \c0.n50\ : std_logic;
signal \c0.n46\ : std_logic;
signal \c0.n56_adj_2146_cascade_\ : std_logic;
signal \c0.n51\ : std_logic;
signal \c0.n9346\ : std_logic;
signal \c0.FRAME_MATCHER_i_3\ : std_logic;
signal \c0.FRAME_MATCHER_i_2\ : std_logic;
signal \c0.FRAME_MATCHER_i_28\ : std_logic;
signal \c0.n45\ : std_logic;
signal \c0.FRAME_MATCHER_i_27\ : std_logic;
signal \c0.FRAME_MATCHER_i_30\ : std_logic;
signal \c0.FRAME_MATCHER_i_8\ : std_logic;
signal \c0.FRAME_MATCHER_i_26\ : std_logic;
signal \c0.n47_adj_2144\ : std_logic;
signal \c0.FRAME_MATCHER_i_22\ : std_logic;
signal \c0.FRAME_MATCHER_i_23\ : std_logic;
signal \c0.FRAME_MATCHER_i_25\ : std_logic;
signal \c0.n49\ : std_logic;
signal \c0.FRAME_MATCHER_state_22\ : std_logic;
signal \c0.n16365\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_12\ : std_logic;
signal \c0.FRAME_MATCHER_i_12\ : std_logic;
signal \c0.n3_adj_2245\ : std_logic;
signal \c0.n16351\ : std_logic;
signal \c0.FRAME_MATCHER_state_21\ : std_logic;
signal \c0.n16367\ : std_logic;
signal \c0.FRAME_MATCHER_state_26\ : std_logic;
signal \c0.n16357\ : std_logic;
signal \c0.FRAME_MATCHER_state_27\ : std_logic;
signal \c0.n16355\ : std_logic;
signal data_in_0_1 : std_logic;
signal \c0.n17266\ : std_logic;
signal data_in_3_5 : std_logic;
signal data_in_2_5 : std_logic;
signal data_in_2_7 : std_logic;
signal \c0.n8_adj_2157\ : std_logic;
signal data_in_3_7 : std_logic;
signal data_in_3_3 : std_logic;
signal data_in_frame_7_0 : std_logic;
signal data_in_frame_7_6 : std_logic;
signal n16896 : std_logic;
signal rx_data_6 : std_logic;
signal rx_data_0 : std_logic;
signal \c0.n2351_cascade_\ : std_logic;
signal data_in_frame_6_7 : std_logic;
signal data_in_frame_6_1 : std_logic;
signal \c0.n2352_cascade_\ : std_logic;
signal data_in_frame_6_3 : std_logic;
signal data_in_frame_6_4 : std_logic;
signal \c0.n23_adj_2145\ : std_logic;
signal \c0.n9541_cascade_\ : std_logic;
signal \c0.n16943\ : std_logic;
signal data_in_frame_0_2 : std_logic;
signal \c0.data_in_frame_2_5\ : std_logic;
signal \c0.data_in_frame_2_3\ : std_logic;
signal \c0.n2336_cascade_\ : std_logic;
signal \c0.data_in_frame_1_5\ : std_logic;
signal \c0.n20_adj_2340_cascade_\ : std_logic;
signal data_in_3_2 : std_logic;
signal data_in_2_2 : std_logic;
signal data_in_1_2 : std_logic;
signal \c0.data_in_frame_10_3\ : std_logic;
signal data_in_frame_6_6 : std_logic;
signal data_in_frame_7_7 : std_logic;
signal data_in_frame_7_2 : std_logic;
signal data_in_frame_6_2 : std_logic;
signal \c0.n22_cascade_\ : std_logic;
signal \c0.n27\ : std_logic;
signal rx_data_7 : std_logic;
signal \c0.data_in_frame_1_0\ : std_logic;
signal n17634 : std_logic;
signal \r_Clock_Count_6_adj_2448\ : std_logic;
signal \c0.n9585\ : std_logic;
signal \c0.data_in_frame_2_2\ : std_logic;
signal \c0.n22_adj_2301\ : std_logic;
signal \c0.n9585_cascade_\ : std_logic;
signal data_in_frame_7_1 : std_logic;
signal data_in_frame_7_4 : std_logic;
signal rx_data_2 : std_logic;
signal data_in_frame_0_0 : std_logic;
signal \c0.data_in_frame_1_6\ : std_logic;
signal \c0.data_in_frame_10_2\ : std_logic;
signal data_in_frame_0_1 : std_logic;
signal \c0.n17460\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \c0.delay_counter_13\ : std_logic;
signal \c0.delay_counter_8\ : std_logic;
signal \c0.delay_counter_4\ : std_logic;
signal \c0.delay_counter_2\ : std_logic;
signal \c0.n17236\ : std_logic;
signal \c0.n42_adj_2165\ : std_logic;
signal \c0.byte_transmit_counter_5\ : std_logic;
signal \c0.n17254\ : std_logic;
signal \c0.n17254_cascade_\ : std_logic;
signal \c0.n17290\ : std_logic;
signal \c0.tx_transmit_N_1949_5\ : std_logic;
signal \c0.n5_adj_2319\ : std_logic;
signal \c0.tx_transmit_N_1949_6\ : std_logic;
signal \c0.byte_transmit_counter_6\ : std_logic;
signal \c0.n23_adj_2309\ : std_logic;
signal \c0.n17278\ : std_logic;
signal \c0.n17276\ : std_logic;
signal \c0.tx_transmit_N_1949_0\ : std_logic;
signal \c0.n16839_cascade_\ : std_logic;
signal \c0.tx_transmit_N_1949_4\ : std_logic;
signal \c0.n8938\ : std_logic;
signal \c0.tx_transmit_N_1949_3\ : std_logic;
signal \c0.n16839\ : std_logic;
signal \c0.tx_transmit_N_1949_7\ : std_logic;
signal \c0.byte_transmit_counter_7\ : std_logic;
signal \n17834_cascade_\ : std_logic;
signal n17162 : std_logic;
signal \n9358_cascade_\ : std_logic;
signal \n41_cascade_\ : std_logic;
signal n35 : std_logic;
signal n29 : std_logic;
signal n445 : std_logic;
signal n10031 : std_logic;
signal \n17479_cascade_\ : std_logic;
signal n16886 : std_logic;
signal n38 : std_logic;
signal \c0.n44_adj_2163\ : std_logic;
signal n9357 : std_logic;
signal \c0.tx_transmit_N_1949_2\ : std_logic;
signal \c0.n4_adj_2311\ : std_logic;
signal \c0.n17475\ : std_logic;
signal \c0.tx2_transmit_N_1997_cascade_\ : std_logic;
signal \c0.tx2.n113\ : std_logic;
signal \c0.tx2.n113_cascade_\ : std_logic;
signal \c0.r_SM_Main_2_N_2036_0_adj_2261\ : std_logic;
signal n491 : std_logic;
signal \n491_cascade_\ : std_logic;
signal n17 : std_logic;
signal \c0.n16369\ : std_logic;
signal \c0.n12_adj_2189\ : std_logic;
signal \c0.FRAME_MATCHER_state_20\ : std_logic;
signal n9460 : std_logic;
signal \n9460_cascade_\ : std_logic;
signal n9462 : std_logic;
signal \c0.FRAME_MATCHER_state_18\ : std_logic;
signal \c0.n16343\ : std_logic;
signal data_in_2_6 : std_logic;
signal rx_data_ready : std_logic;
signal data_in_1_6 : std_logic;
signal \c0.n8603\ : std_logic;
signal \c0.FRAME_MATCHER_i_11\ : std_logic;
signal \c0.FRAME_MATCHER_i_14\ : std_logic;
signal \c0.FRAME_MATCHER_i_15\ : std_logic;
signal \c0.n48\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_10\ : std_logic;
signal \c0.FRAME_MATCHER_i_10\ : std_logic;
signal \c0.n3_adj_2247\ : std_logic;
signal \c0.n9819_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_25\ : std_logic;
signal \c0.n16359\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_17\ : std_logic;
signal \c0.FRAME_MATCHER_i_17\ : std_logic;
signal \c0.n3_adj_2240\ : std_logic;
signal data_in_frame_0_7 : std_logic;
signal \c0.data_in_frame_1_7\ : std_logic;
signal \c0.data_in_frame_1_4\ : std_logic;
signal \c0.n27_adj_2342\ : std_logic;
signal \c0.n23_adj_2341_cascade_\ : std_logic;
signal \c0.data_in_frame_1_3\ : std_logic;
signal \c0.n21_adj_2171\ : std_logic;
signal \c0.n15930\ : std_logic;
signal \c0.data_in_frame_10_7\ : std_logic;
signal \c0.n17352_cascade_\ : std_logic;
signal \c0.n27_adj_2196\ : std_logic;
signal \c0.n25\ : std_logic;
signal \c0.n15846_cascade_\ : std_logic;
signal \c0.n15929\ : std_logic;
signal \c0.n26_adj_2184\ : std_logic;
signal \c0.n15938\ : std_logic;
signal \c0.data_in_frame_1_2\ : std_logic;
signal \c0.data_in_frame_9_3\ : std_logic;
signal \c0.data_in_frame_1_1\ : std_logic;
signal \c0.n17014\ : std_logic;
signal \c0.n23_adj_2156_cascade_\ : std_logic;
signal \c0.n17001\ : std_logic;
signal \c0.n28_adj_2183\ : std_logic;
signal data_in_frame_0_6 : std_logic;
signal \c0.n2340\ : std_logic;
signal \c0.data_in_frame_9_0\ : std_logic;
signal \c0.n17004\ : std_logic;
signal \c0.n19\ : std_logic;
signal data_in_frame_7_3 : std_logic;
signal \c0.n2336\ : std_logic;
signal data_in_frame_7_5 : std_logic;
signal \c0.n9541\ : std_logic;
signal data_in_frame_6_0 : std_logic;
signal data_in_frame_6_5 : std_logic;
signal \c0.n20_cascade_\ : std_logic;
signal \c0.n2342\ : std_logic;
signal \c0.data_in_frame_9_1\ : std_logic;
signal \c0.n8_adj_2310\ : std_logic;
signal \c0.data_in_frame_9_5\ : std_logic;
signal tx2_o : std_logic;
signal \c0.tx2.n18113_cascade_\ : std_logic;
signal n10398 : std_logic;
signal n17194 : std_logic;
signal \n10398_cascade_\ : std_logic;
signal \c0.tx2.n17906\ : std_logic;
signal \c0.tx2.n18116\ : std_logic;
signal \c0.tx2.o_Tx_Serial_N_2064_cascade_\ : std_logic;
signal \r_SM_Main_0_adj_2445\ : std_logic;
signal n3 : std_logic;
signal n5029 : std_logic;
signal \r_Bit_Index_2_adj_2455\ : std_logic;
signal \c0.tx2.n13281\ : std_logic;
signal \c0.n2_adj_2266_cascade_\ : std_logic;
signal \c0.n18098_cascade_\ : std_logic;
signal \c0.n10_adj_2139_cascade_\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal n17394 : std_logic;
signal \c0.n8_adj_2160\ : std_logic;
signal \c0.n15_cascade_\ : std_logic;
signal \c0.n12_adj_2150_cascade_\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal n10_adj_2426 : std_logic;
signal \n10_adj_2407_cascade_\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \c0.n17590_cascade_\ : std_logic;
signal n18026 : std_logic;
signal \c0.n16347\ : std_logic;
signal \c0.n16761\ : std_logic;
signal \c0.FRAME_MATCHER_state_28\ : std_logic;
signal \c0.n16353\ : std_logic;
signal \c0.FRAME_MATCHER_state_24\ : std_logic;
signal \c0.n16361\ : std_logic;
signal \c0.FRAME_MATCHER_state_17\ : std_logic;
signal \c0.n16345\ : std_logic;
signal \c0.FRAME_MATCHER_state_4\ : std_logic;
signal \c0.n4\ : std_logic;
signal \c0.n16339\ : std_logic;
signal \c0.FRAME_MATCHER_state_14\ : std_logic;
signal \c0.n16871\ : std_logic;
signal \c0.n16772\ : std_logic;
signal \c0.n17349_cascade_\ : std_logic;
signal \c0.n1439\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1312_0\ : std_logic;
signal \c0.n5_adj_2322\ : std_logic;
signal \c0.n5_cascade_\ : std_logic;
signal \c0.n17328_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_8\ : std_logic;
signal \c0.n16905\ : std_logic;
signal \c0.n17337_cascade_\ : std_logic;
signal data_in_frame_0_4 : std_logic;
signal data_in_frame_0_5 : std_logic;
signal \c0.n2338\ : std_logic;
signal \c0.data_in_frame_2_6\ : std_logic;
signal \c0.data_in_frame_2_0\ : std_logic;
signal \c0.n2338_cascade_\ : std_logic;
signal \c0.n2352\ : std_logic;
signal \c0.n26_adj_2344\ : std_logic;
signal \c0.n17_adj_2346_cascade_\ : std_logic;
signal \c0.n30_adj_2345\ : std_logic;
signal \n31_cascade_\ : std_logic;
signal \c0.tx2.tx2_active\ : std_logic;
signal \c0.n17334_cascade_\ : std_logic;
signal \c0.n2334\ : std_logic;
signal \c0.n2351\ : std_logic;
signal \c0.n18_adj_2343\ : std_logic;
signal rx_data_3 : std_logic;
signal n16897 : std_logic;
signal data_in_frame_0_3 : std_logic;
signal \c0.n17918_cascade_\ : std_logic;
signal \c0.n17343\ : std_logic;
signal \c0.n17769\ : std_logic;
signal \c0.n18\ : std_logic;
signal \c0.n17\ : std_logic;
signal \c0.n26_adj_2147\ : std_logic;
signal \c0.n30_adj_2148\ : std_logic;
signal rx_data_5 : std_logic;
signal \c0.n16882\ : std_logic;
signal \c0.data_in_frame_10_5\ : std_logic;
signal \r_SM_Main_1_adj_2444\ : std_logic;
signal \c0.tx2.n6480\ : std_logic;
signal \c0.tx2.n1\ : std_logic;
signal \c0.tx2.n10101\ : std_logic;
signal data_out_frame2_18_5 : std_logic;
signal \r_SM_Main_2_adj_2439\ : std_logic;
signal n13440 : std_logic;
signal \r_SM_Main_1_adj_2440\ : std_logic;
signal rx_data_1 : std_logic;
signal \c0.data_in_frame_2_1\ : std_logic;
signal \c0.n16891\ : std_logic;
signal \c0.n8\ : std_logic;
signal rx_data_4 : std_logic;
signal \c0.data_in_frame_2_4\ : std_logic;
signal \c0.r_SM_Main_2_N_2036_0\ : std_logic;
signal tx_active : std_logic;
signal n17230 : std_logic;
signal data_out_1_7 : std_logic;
signal \c0.n10\ : std_logic;
signal \r_SM_Main_2_adj_2443\ : std_logic;
signal n17544 : std_logic;
signal \r_Clock_Count_0_adj_2454\ : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal n17398 : std_logic;
signal \c0.n29_cascade_\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \c0.data_out_0_6\ : std_logic;
signal \c0.n9_adj_2143_cascade_\ : std_logic;
signal \c0.n23\ : std_logic;
signal \c0.n17547\ : std_logic;
signal \c0.n5_adj_2326_cascade_\ : std_logic;
signal \c0.n18023\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \c0.n18014\ : std_logic;
signal \c0.n17585\ : std_logic;
signal n10_adj_2423 : std_logic;
signal \n18044_cascade_\ : std_logic;
signal n10_adj_2414 : std_logic;
signal data_out_0_1 : std_logic;
signal \c0.n18080\ : std_logic;
signal data_out_3_7 : std_logic;
signal \c0.n2_adj_2137\ : std_logic;
signal \c0.data_out_1_4\ : std_logic;
signal n16776 : std_logic;
signal n17208 : std_logic;
signal n8828 : std_logic;
signal \c0.FRAME_MATCHER_state_16\ : std_logic;
signal \c0.n47\ : std_logic;
signal \c0.n6_adj_2140\ : std_logic;
signal \FRAME_MATCHER_state_1\ : std_logic;
signal \c0.n5_adj_2339\ : std_logic;
signal \c0.n16814_cascade_\ : std_logic;
signal \c0.tx2.n89\ : std_logic;
signal \c0.FRAME_MATCHER_state_31\ : std_logic;
signal \c0.n16377\ : std_logic;
signal n9452 : std_logic;
signal n12933 : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1280_0\ : std_logic;
signal \c0.FRAME_MATCHER_i_0\ : std_logic;
signal \c0.n3\ : std_logic;
signal \c0.FRAME_MATCHER_state_12\ : std_logic;
signal \c0.n4_adj_2360\ : std_logic;
signal \c0.n16449\ : std_logic;
signal data_out_frame2_18_2 : std_logic;
signal \c0.n18119_cascade_\ : std_logic;
signal \c0.n18122_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_2\ : std_logic;
signal \c0.n17340\ : std_logic;
signal \c0.n13496\ : std_logic;
signal data_out_frame2_7_3 : std_logic;
signal \FRAME_MATCHER_state_2\ : std_logic;
signal \c0.FRAME_MATCHER_state_3\ : std_logic;
signal \c0.n62\ : std_logic;
signal \c0.n13464\ : std_logic;
signal \c0.n2_adj_2330_cascade_\ : std_logic;
signal \c0.n9758\ : std_logic;
signal \c0.n17915\ : std_logic;
signal data_out_frame2_18_1 : std_logic;
signal \c0.n17909_cascade_\ : std_logic;
signal \c0.n6\ : std_logic;
signal \c0.n18107\ : std_logic;
signal \c0.n17579\ : std_logic;
signal \c0.n17912\ : std_logic;
signal \c0.n18110\ : std_logic;
signal \c0.n22_adj_2359_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_1\ : std_logic;
signal \c0.n17548\ : std_logic;
signal \c0.n17589\ : std_logic;
signal \c0.n2_adj_2298\ : std_logic;
signal \c0.n18029_cascade_\ : std_logic;
signal \c0.n8_adj_2138\ : std_logic;
signal \c0.n5_adj_2299\ : std_logic;
signal \r_SM_Main_0_adj_2441\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2096_0\ : std_logic;
signal \r_Rx_Data\ : std_logic;
signal n1 : std_logic;
signal data_out_3_5 : std_logic;
signal data_out_2_5 : std_logic;
signal \c0.n9530\ : std_logic;
signal data_out_1_6 : std_logic;
signal data_out_2_0 : std_logic;
signal \c0.n9509\ : std_logic;
signal \c0.data_out_7_5\ : std_logic;
signal \c0.n26\ : std_logic;
signal n18032 : std_logic;
signal n10 : std_logic;
signal \c0.n5_adj_2142\ : std_logic;
signal data_out_3_0 : std_logic;
signal \c0.data_out_3_6\ : std_logic;
signal \c0.n10054_cascade_\ : std_logic;
signal \c0.data_out_7_7\ : std_logic;
signal \c0.n5_adj_2188_cascade_\ : std_logic;
signal \c0.n18041\ : std_logic;
signal \c0.n5_adj_2208\ : std_logic;
signal \c0.n17543_cascade_\ : std_logic;
signal \c0.n18011\ : std_logic;
signal \c0.n17445\ : std_logic;
signal \c0.n17456_cascade_\ : std_logic;
signal \c0.n10054\ : std_logic;
signal n9361 : std_logic;
signal n17154 : std_logic;
signal \FRAME_MATCHER_state_0\ : std_logic;
signal \c0.tx2_transmit_N_1997\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \c0.n15615\ : std_logic;
signal \c0.n15616\ : std_logic;
signal \c0.n15617\ : std_logic;
signal \c0.n15618\ : std_logic;
signal \c0.byte_transmit_counter2_5\ : std_logic;
signal \c0.n15619\ : std_logic;
signal \c0.byte_transmit_counter2_6\ : std_logic;
signal \c0.n15620\ : std_logic;
signal \c0.n15621\ : std_logic;
signal \c0.byte_transmit_counter2_7\ : std_logic;
signal \c0.n10052\ : std_logic;
signal \c0.n10297\ : std_logic;
signal \c0.n7\ : std_logic;
signal \c0.FRAME_MATCHER_state_9\ : std_logic;
signal \c0.n16455\ : std_logic;
signal \c0.n17927\ : std_logic;
signal data_out_frame2_17_2 : std_logic;
signal \c0.n17930_cascade_\ : std_logic;
signal \c0.n22_adj_2358\ : std_logic;
signal \c0.n17936\ : std_logic;
signal \c0.n6_adj_2201\ : std_logic;
signal \c0.n17942\ : std_logic;
signal \c0.n17560\ : std_logic;
signal \c0.n17301_cascade_\ : std_logic;
signal \c0.n17303_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_0\ : std_logic;
signal data_out_frame2_18_0 : std_logic;
signal data_out_frame2_17_0 : std_logic;
signal \c0.n18101_cascade_\ : std_logic;
signal \c0.n18104_cascade_\ : std_logic;
signal \c0.n22_adj_2337\ : std_logic;
signal \c0.n17939\ : std_logic;
signal data_out_frame2_6_3 : std_logic;
signal \c0.n16_adj_2197\ : std_logic;
signal \c0.n22_adj_2194\ : std_logic;
signal \c0.n9754\ : std_logic;
signal \c0.n9901_cascade_\ : std_logic;
signal data_out_frame2_5_3 : std_logic;
signal \c0.n16148\ : std_logic;
signal \c0.n17331_cascade_\ : std_logic;
signal \c0.n15846\ : std_logic;
signal \c0.n17891\ : std_logic;
signal data_out_frame2_10_2 : std_logic;
signal \c0.n12_adj_2305\ : std_logic;
signal \c0.n17990\ : std_logic;
signal \c0.n17993_cascade_\ : std_logic;
signal \c0.n17894\ : std_logic;
signal \c0.n17393_cascade_\ : std_logic;
signal \c0.n17571\ : std_logic;
signal \c0.n17963_cascade_\ : std_logic;
signal \c0.n17966_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_5\ : std_logic;
signal data_out_0_5 : std_logic;
signal data_out_0_3 : std_logic;
signal data_out_2_2 : std_logic;
signal \c0.n2_adj_2291\ : std_logic;
signal data_out_3_2 : std_logic;
signal data_out_frame2_9_4 : std_logic;
signal \c0.n9_adj_2347\ : std_logic;
signal \c0.n17897\ : std_logic;
signal \c0.n8_adj_2348_cascade_\ : std_logic;
signal \c0.n17900\ : std_logic;
signal \r_Bit_Index_1_adj_2456\ : std_logic;
signal \r_Bit_Index_0_adj_2457\ : std_logic;
signal \c0.tx2.n17903\ : std_logic;
signal \c0.n16975\ : std_logic;
signal \c0.n16978_cascade_\ : std_logic;
signal \c0.n16912\ : std_logic;
signal \c0.n21\ : std_logic;
signal \c0.n17588\ : std_logic;
signal \c0.n1\ : std_logic;
signal \n18038_cascade_\ : std_logic;
signal n8730 : std_logic;
signal \n10_adj_2413_cascade_\ : std_logic;
signal byte_transmit_counter_4 : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \c0.data_out_1_1\ : std_logic;
signal \c0.n10181\ : std_logic;
signal \c0.data_out_6_6\ : std_logic;
signal \c0.n5_adj_2300\ : std_logic;
signal \c0.n17555_cascade_\ : std_logic;
signal \c0.n18035\ : std_logic;
signal \c0.n17569\ : std_logic;
signal \c0.data_out_frame2_0_2\ : std_logic;
signal \c0.n17578\ : std_logic;
signal \c0.data_out_frame2_0_4\ : std_logic;
signal \c0.n6_adj_2335\ : std_logic;
signal \c0.n5_adj_2317\ : std_logic;
signal \c0.n16957\ : std_logic;
signal \c0.n17106\ : std_logic;
signal \c0.n16957_cascade_\ : std_logic;
signal \c0.n15_adj_2269\ : std_logic;
signal \c0.data_out_frame2_20_1\ : std_logic;
signal \c0.n17061\ : std_logic;
signal \c0.data_out_frame2_20_0\ : std_logic;
signal \c0.n9810\ : std_logic;
signal \c0.n17_adj_2193\ : std_logic;
signal \c0.n16_cascade_\ : std_logic;
signal \c0.n17112_cascade_\ : std_logic;
signal \c0.n14_adj_2308_cascade_\ : std_logic;
signal \c0.data_out_frame2_19_5\ : std_logic;
signal \c0.n17933\ : std_logic;
signal data_out_frame2_15_3 : std_logic;
signal data_out_frame2_13_4 : std_logic;
signal \c0.n11\ : std_logic;
signal \c0.n17981\ : std_logic;
signal \c0.n17984_cascade_\ : std_logic;
signal \c0.n22_adj_2354\ : std_logic;
signal data_out_frame2_17_5 : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal n15528 : std_logic;
signal n15529 : std_logic;
signal n15530 : std_logic;
signal n15531 : std_logic;
signal n15532 : std_logic;
signal n15533 : std_logic;
signal n15534 : std_logic;
signal n15535 : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal n15536 : std_logic;
signal n15537 : std_logic;
signal n15538 : std_logic;
signal n15539 : std_logic;
signal n15540 : std_logic;
signal n15541 : std_logic;
signal n15542 : std_logic;
signal n15543 : std_logic;
signal \bfn_13_27_0_\ : std_logic;
signal n15544 : std_logic;
signal n15545 : std_logic;
signal n15546 : std_logic;
signal n15547 : std_logic;
signal n15548 : std_logic;
signal n15549 : std_logic;
signal n15550 : std_logic;
signal n15551 : std_logic;
signal \bfn_13_28_0_\ : std_logic;
signal n15552 : std_logic;
signal n15553 : std_logic;
signal n15554 : std_logic;
signal n15555 : std_logic;
signal n15556 : std_logic;
signal n15557 : std_logic;
signal n15558 : std_logic;
signal rand_setpoint_0 : std_logic;
signal \bfn_13_29_0_\ : std_logic;
signal rand_data_1 : std_logic;
signal n15559 : std_logic;
signal rand_data_2 : std_logic;
signal n15560 : std_logic;
signal rand_setpoint_3 : std_logic;
signal n15561 : std_logic;
signal rand_setpoint_4 : std_logic;
signal n15562 : std_logic;
signal n15563 : std_logic;
signal n15564 : std_logic;
signal n15565 : std_logic;
signal n15566 : std_logic;
signal rand_setpoint_8 : std_logic;
signal \bfn_13_30_0_\ : std_logic;
signal rand_setpoint_9 : std_logic;
signal n15567 : std_logic;
signal rand_data_10 : std_logic;
signal n15568 : std_logic;
signal rand_setpoint_11 : std_logic;
signal n15569 : std_logic;
signal rand_setpoint_12 : std_logic;
signal n15570 : std_logic;
signal rand_setpoint_13 : std_logic;
signal n15571 : std_logic;
signal rand_setpoint_14 : std_logic;
signal n15572 : std_logic;
signal rand_setpoint_15 : std_logic;
signal n15573 : std_logic;
signal n15574 : std_logic;
signal \bfn_13_31_0_\ : std_logic;
signal n15575 : std_logic;
signal n15576 : std_logic;
signal rand_data_19 : std_logic;
signal n15577 : std_logic;
signal n15578 : std_logic;
signal n15579 : std_logic;
signal rand_setpoint_22 : std_logic;
signal n15580 : std_logic;
signal n15581 : std_logic;
signal n15582 : std_logic;
signal \bfn_13_32_0_\ : std_logic;
signal rand_setpoint_25 : std_logic;
signal n15583 : std_logic;
signal n15584 : std_logic;
signal n15585 : std_logic;
signal n15586 : std_logic;
signal n15587 : std_logic;
signal rand_setpoint_30 : std_logic;
signal n15588 : std_logic;
signal n15589 : std_logic;
signal rand_setpoint_31 : std_logic;
signal \c0.data_out_7_4\ : std_logic;
signal \c0.n22_adj_2357_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_3\ : std_logic;
signal \c0.n6_adj_2187\ : std_logic;
signal \c0.n18128\ : std_logic;
signal \c0.n16936\ : std_logic;
signal \c0.n18_adj_2331\ : std_logic;
signal \c0.n17100_cascade_\ : std_logic;
signal \c0.n16_adj_2332_cascade_\ : std_logic;
signal \c0.n20_adj_2333\ : std_logic;
signal \c0.data_out_frame2_19_0\ : std_logic;
signal \c0.n9886\ : std_logic;
signal \c0.n12_adj_2263_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_2\ : std_logic;
signal \c0.n17112\ : std_logic;
signal \c0.n16_adj_2312_cascade_\ : std_logic;
signal \c0.n17097\ : std_logic;
signal data_out_frame2_6_0 : std_logic;
signal \c0.n5_adj_2334\ : std_logic;
signal \c0.data_out_frame2_0_1\ : std_logic;
signal \c0.n17124\ : std_logic;
signal \c0.n14_adj_2264\ : std_logic;
signal data_out_frame2_16_2 : std_logic;
signal \c0.n17031\ : std_logic;
signal \c0.n17091\ : std_logic;
signal \c0.n17031_cascade_\ : std_logic;
signal \c0.n9692\ : std_logic;
signal \c0.n17085\ : std_logic;
signal data_out_frame2_9_3 : std_logic;
signal \c0.n17085_cascade_\ : std_logic;
signal \c0.n17073\ : std_logic;
signal data_out_frame2_18_4 : std_logic;
signal \c0.data_out_frame2_19_4\ : std_logic;
signal \c0.n9707\ : std_logic;
signal \c0.n16963\ : std_logic;
signal \c0.n9579\ : std_logic;
signal \c0.n9579_cascade_\ : std_logic;
signal \c0.n10_adj_2307\ : std_logic;
signal \c0.n17957\ : std_logic;
signal \c0.n16908\ : std_logic;
signal \c0.n16908_cascade_\ : std_logic;
signal \c0.n6_adj_2286\ : std_logic;
signal data_out_frame2_14_4 : std_logic;
signal \c0.n5543\ : std_logic;
signal \c0.n5545\ : std_logic;
signal n31 : std_logic;
signal rand_data_4 : std_logic;
signal \n10197_cascade_\ : std_logic;
signal data_out_frame2_15_4 : std_logic;
signal data_out_frame2_12_5 : std_logic;
signal \c0.n17049\ : std_logic;
signal data_out_frame2_5_2 : std_logic;
signal \c0.n9865\ : std_logic;
signal \c0.n6_adj_2306_cascade_\ : std_logic;
signal rand_data_27 : std_logic;
signal rand_data_9 : std_logic;
signal data_out_frame2_17_1 : std_logic;
signal data_out_frame2_10_4 : std_logic;
signal \c0.n10_adj_2191\ : std_logic;
signal \c0.n14\ : std_logic;
signal \c0.n17528\ : std_logic;
signal data_out_9_2 : std_logic;
signal \c0.n17064\ : std_logic;
signal \c0.n12_adj_2289_cascade_\ : std_logic;
signal \c0.data_out_7_6\ : std_logic;
signal \c0.n9716_cascade_\ : std_logic;
signal \c0.n9728\ : std_logic;
signal \c0.n10_adj_2162_cascade_\ : std_logic;
signal \data_out_9__2__N_367\ : std_logic;
signal \data_out_9__2__N_367_cascade_\ : std_logic;
signal rand_setpoint_7 : std_logic;
signal \c0.n8_adj_2169_cascade_\ : std_logic;
signal n10_adj_2427 : std_logic;
signal \c0.n9496\ : std_logic;
signal \c0.n9716\ : std_logic;
signal rand_setpoint_2 : std_logic;
signal \c0.n17594\ : std_logic;
signal \c0.n8_adj_2176\ : std_logic;
signal \c0.data_out_1_2\ : std_logic;
signal data_out_2_7 : std_logic;
signal rand_setpoint_20 : std_logic;
signal \c0.n17518\ : std_logic;
signal rand_setpoint_19 : std_logic;
signal \c0.n17514\ : std_logic;
signal rand_setpoint_18 : std_logic;
signal \c0.n17507\ : std_logic;
signal rand_setpoint_17 : std_logic;
signal \c0.n17506_cascade_\ : std_logic;
signal rand_setpoint_26 : std_logic;
signal rand_setpoint_29 : std_logic;
signal rand_setpoint_24 : std_logic;
signal rand_setpoint_27 : std_logic;
signal rand_setpoint_28 : std_logic;
signal data_out_frame2_7_1 : std_logic;
signal data_out_frame2_10_5 : std_logic;
signal \c0.n9763\ : std_logic;
signal data_out_frame2_8_2 : std_logic;
signal \c0.n9916\ : std_logic;
signal data_out_frame2_12_4 : std_logic;
signal \c0.n17037\ : std_logic;
signal \c0.n16933_cascade_\ : std_logic;
signal \c0.n17_adj_2313\ : std_logic;
signal \c0.n17960\ : std_logic;
signal \c0.n18125\ : std_logic;
signal \c0.n15_adj_2320_cascade_\ : std_logic;
signal \c0.n17088\ : std_logic;
signal \c0.data_out_frame2_19_2\ : std_logic;
signal \c0.n14_adj_2323\ : std_logic;
signal \c0.n17052\ : std_logic;
signal \c0.n17121\ : std_logic;
signal \c0.n19_adj_2254\ : std_logic;
signal \c0.n21_adj_2255_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_3\ : std_logic;
signal data_out_frame2_14_5 : std_logic;
signal \c0.n17022\ : std_logic;
signal \c0.n26_adj_2273\ : std_logic;
signal \c0.data_out_frame2_0_5\ : std_logic;
signal \c0.n17103\ : std_logic;
signal \c0.n17067\ : std_logic;
signal \c0.n17100\ : std_logic;
signal \c0.n9749\ : std_logic;
signal data_out_frame2_5_1 : std_logic;
signal \c0.n9776\ : std_logic;
signal \c0.n9555\ : std_logic;
signal \c0.n16946\ : std_logic;
signal \c0.n22_adj_2207_cascade_\ : std_logic;
signal \c0.n18_adj_2251\ : std_logic;
signal \c0.n9892_cascade_\ : std_logic;
signal \c0.n17079\ : std_logic;
signal \c0.n20_adj_2202\ : std_logic;
signal \c0.n17079_cascade_\ : std_logic;
signal \c0.n24\ : std_logic;
signal \c0.data_out_frame2_20_5\ : std_logic;
signal data_out_frame2_10_7 : std_logic;
signal rand_data_28 : std_logic;
signal data_out_frame2_15_2 : std_logic;
signal data_out_frame2_16_1 : std_logic;
signal rand_data_20 : std_logic;
signal \c0.n9814\ : std_logic;
signal \c0.n16987\ : std_logic;
signal \c0.n25_adj_2275\ : std_logic;
signal rand_data_17 : std_logic;
signal data_out_frame2_6_4 : std_logic;
signal \c0.n5_adj_2141_cascade_\ : std_logic;
signal \c0.n17987\ : std_logic;
signal \c0.n17951\ : std_logic;
signal data_out_frame2_13_3 : std_logic;
signal \c0.n17954\ : std_logic;
signal \c0.n18056\ : std_logic;
signal data_out_frame2_7_0 : std_logic;
signal \c0.n17346\ : std_logic;
signal rand_data_26 : std_logic;
signal data_out_frame2_14_2 : std_logic;
signal rand_data_0 : std_logic;
signal data_out_frame2_9_0 : std_logic;
signal \c0.n32_adj_2297\ : std_logic;
signal \c0.data_out_6_4\ : std_logic;
signal \c0.data_out_10_0\ : std_logic;
signal \c0.n16966\ : std_logic;
signal \c0.n16966_cascade_\ : std_logic;
signal \c0.n16918\ : std_logic;
signal \c0.n10_adj_2288_cascade_\ : std_logic;
signal \c0.n17109\ : std_logic;
signal \c0.n16990\ : std_logic;
signal \c0.data_out_6_1\ : std_logic;
signal rand_setpoint_5 : std_logic;
signal data_out_8_5 : std_logic;
signal \c0.n28_adj_2287\ : std_logic;
signal rand_setpoint_6 : std_logic;
signal data_out_8_6 : std_logic;
signal \c0.data_out_10_7\ : std_logic;
signal \c0.n8_adj_2166\ : std_logic;
signal n10_adj_2425 : std_logic;
signal \c0.n17055\ : std_logic;
signal \c0.data_out_9_5\ : std_logic;
signal \c0.data_out_10_1\ : std_logic;
signal \c0.data_out_8_2\ : std_logic;
signal \c0.data_out_10_5\ : std_logic;
signal rand_setpoint_1 : std_logic;
signal \c0.data_out_7_1\ : std_logic;
signal \c0.data_out_9_0\ : std_logic;
signal \c0.data_out_5_2\ : std_logic;
signal \c0.n9522\ : std_logic;
signal data_out_8_1 : std_logic;
signal \c0.n18077\ : std_logic;
signal \c0.data_out_7__2__N_447\ : std_logic;
signal rand_setpoint_23 : std_logic;
signal \c0.n17532_cascade_\ : std_logic;
signal \c0.data_out_6_7\ : std_logic;
signal \c0.data_out_5_5\ : std_logic;
signal \c0.n17025\ : std_logic;
signal \c0.n17534\ : std_logic;
signal \c0.data_out_frame2_0_3\ : std_logic;
signal \c0.n17576\ : std_logic;
signal data_out_frame2_8_3 : std_logic;
signal \c0.n9839\ : std_logic;
signal data_out_frame2_18_6 : std_logic;
signal \c0.n16994\ : std_logic;
signal rand_data_21 : std_logic;
signal \c0.n28_adj_2294\ : std_logic;
signal \c0.n32_cascade_\ : std_logic;
signal \c0.n31\ : std_logic;
signal \c0.n29_adj_2296\ : std_logic;
signal \c0.n16933\ : std_logic;
signal \c0.n16915_cascade_\ : std_logic;
signal data_out_frame2_7_2 : std_logic;
signal \c0.n19_adj_2303\ : std_logic;
signal \c0.n20_adj_2302_cascade_\ : std_logic;
signal \c0.n21_adj_2304\ : std_logic;
signal \c0.data_out_frame2_19_6\ : std_logic;
signal \c0.data_out_frame2_0_0\ : std_logic;
signal \c0.n16972_cascade_\ : std_logic;
signal data_out_frame2_11_2 : std_logic;
signal \c0.n10_adj_2281\ : std_logic;
signal \c0.n17969\ : std_logic;
signal data_out_frame2_16_4 : std_logic;
signal \c0.data_out_frame2_20_4\ : std_logic;
signal \c0.n17972_cascade_\ : std_logic;
signal \c0.n17040\ : std_logic;
signal \c0.n16972\ : std_logic;
signal \c0.n30_adj_2295\ : std_logic;
signal data_out_frame2_7_7 : std_logic;
signal \c0.n5_adj_2351\ : std_logic;
signal data_out_frame2_11_3 : std_logic;
signal \c0.n9695\ : std_logic;
signal \c0.n9695_cascade_\ : std_logic;
signal rand_data_22 : std_logic;
signal data_out_frame2_11_7 : std_logic;
signal data_out_frame2_11_5 : std_logic;
signal \c0.n9919\ : std_logic;
signal \c0.n9901\ : std_logic;
signal \c0.n10_adj_2292\ : std_logic;
signal data_out_frame2_7_4 : std_logic;
signal \c0.n9913\ : std_logic;
signal \c0.n17034\ : std_logic;
signal \c0.n17034_cascade_\ : std_logic;
signal \c0.n9688\ : std_logic;
signal data_out_frame2_12_1 : std_logic;
signal \c0.n9688_cascade_\ : std_logic;
signal \c0.n6_adj_2325\ : std_logic;
signal data_out_frame2_11_1 : std_logic;
signal data_out_frame2_6_1 : std_logic;
signal \c0.n17115\ : std_logic;
signal rand_data_5 : std_logic;
signal data_out_frame2_16_5 : std_logic;
signal data_out_frame2_8_5 : std_logic;
signal data_out_frame2_10_3 : std_logic;
signal \c0.n20_adj_2252\ : std_logic;
signal \c0.n17322\ : std_logic;
signal \c0.n17323_cascade_\ : std_logic;
signal \c0.n18053\ : std_logic;
signal rand_data_16 : std_logic;
signal data_out_frame2_9_1 : std_logic;
signal \c0.n17921\ : std_logic;
signal \c0.n17924\ : std_logic;
signal data_out_frame2_18_7 : std_logic;
signal \c0.data_out_frame2_19_7\ : std_logic;
signal \c0.n18059_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_7\ : std_logic;
signal \c0.n18062_cascade_\ : std_logic;
signal data_out_frame2_11_4 : std_logic;
signal data_out_frame2_17_7 : std_logic;
signal data_out_frame2_14_0 : std_logic;
signal \c0.n9853\ : std_logic;
signal \c0.n9589\ : std_logic;
signal \c0.n9853_cascade_\ : std_logic;
signal data_out_frame2_13_0 : std_logic;
signal \c0.n17046\ : std_logic;
signal \c0.n17581\ : std_logic;
signal \c0.n10259\ : std_logic;
signal \c0.data_out_7_3\ : std_logic;
signal \c0.n8_adj_2153\ : std_logic;
signal \c0.n17070\ : std_logic;
signal \c0.n9737\ : std_logic;
signal \c0.n12_adj_2285\ : std_logic;
signal \c0.data_out_6_3\ : std_logic;
signal \c0.data_out_2_3\ : std_logic;
signal n2652 : std_logic;
signal \c0.n5_adj_2350\ : std_logic;
signal \c0.n17546_cascade_\ : std_logic;
signal \c0.n17592\ : std_logic;
signal \c0.n18017_cascade_\ : std_logic;
signal \c0.n17593\ : std_logic;
signal \c0.n10_adj_2154\ : std_logic;
signal \c0.n18020_cascade_\ : std_logic;
signal byte_transmit_counter_3 : std_logic;
signal \c0.n10_adj_2155\ : std_logic;
signal \c0.n10_adj_2268\ : std_logic;
signal \c0.data_out_8_3\ : std_logic;
signal data_out_8_4 : std_logic;
signal \c0.data_out_9_1\ : std_logic;
signal data_out_3_4 : std_logic;
signal \c0.n17591\ : std_logic;
signal rand_setpoint_16 : std_logic;
signal n2547 : std_logic;
signal \UART_TRANSMITTER_state_2\ : std_logic;
signal \c0.data_out_5_3\ : std_logic;
signal \c0.data_out_5_4\ : std_logic;
signal \c0.n9783\ : std_logic;
signal data_out_frame2_10_6 : std_logic;
signal data_out_frame2_5_4 : std_logic;
signal \c0.n17495\ : std_logic;
signal data_out_frame2_9_6 : std_logic;
signal \c0.n18047\ : std_logic;
signal \c0.n9859\ : std_logic;
signal data_out_frame2_13_2 : std_logic;
signal \c0.n17133\ : std_logic;
signal \c0.n27_adj_2277\ : std_logic;
signal data_out_frame2_8_6 : std_logic;
signal data_out_frame2_6_6 : std_logic;
signal \c0.n18050\ : std_logic;
signal \c0.n9671\ : std_logic;
signal \c0.n17016\ : std_logic;
signal \c0.n6_adj_2293\ : std_logic;
signal \c0.n16960\ : std_logic;
signal \c0.n24_adj_2272\ : std_logic;
signal data_out_frame2_9_2 : std_logic;
signal data_out_frame2_16_0 : std_logic;
signal \c0.n9892\ : std_logic;
signal \c0.n20_adj_2205\ : std_logic;
signal \c0.n18071\ : std_logic;
signal \c0.n18074_cascade_\ : std_logic;
signal data_out_frame2_12_7 : std_logic;
signal data_out_frame2_13_7 : std_logic;
signal \c0.n18065_cascade_\ : std_logic;
signal \c0.n18068\ : std_logic;
signal data_out_frame2_14_6 : std_logic;
signal data_out_frame2_12_6 : std_logic;
signal \c0.n18005_cascade_\ : std_logic;
signal \c0.n18008\ : std_logic;
signal data_out_frame2_10_0 : std_logic;
signal \c0.n17347\ : std_logic;
signal rand_data_18 : std_logic;
signal data_out_frame2_6_2 : std_logic;
signal data_out_frame2_15_6 : std_logic;
signal data_out_frame2_7_6 : std_logic;
signal \c0.n17127\ : std_logic;
signal data_out_frame2_8_7 : std_logic;
signal data_out_frame2_11_6 : std_logic;
signal data_out_frame2_14_7 : std_logic;
signal rand_data_12 : std_logic;
signal data_out_frame2_17_4 : std_logic;
signal rand_data_23 : std_logic;
signal data_out_frame2_6_7 : std_logic;
signal rand_data_31 : std_logic;
signal data_out_frame2_5_7 : std_logic;
signal rand_data_15 : std_logic;
signal data_out_frame2_9_7 : std_logic;
signal data_out_frame2_9_5 : std_logic;
signal \c0.n16926\ : std_logic;
signal rand_data_24 : std_logic;
signal data_out_frame2_5_0 : std_logic;
signal rand_data_25 : std_logic;
signal data_out_frame2_6_5 : std_logic;
signal data_out_frame2_5_5 : std_logic;
signal \c0.n5_adj_2349_cascade_\ : std_logic;
signal \c0.n6_adj_2280\ : std_logic;
signal rand_data_13 : std_logic;
signal \c0.n6_adj_2278\ : std_logic;
signal \c0.n18089\ : std_logic;
signal \c0.n17561\ : std_logic;
signal data_out_frame2_7_5 : std_logic;
signal \c0.n9678\ : std_logic;
signal \c0.n18092\ : std_logic;
signal \c0.n22_adj_2352\ : std_logic;
signal \c0.tx2.r_Tx_Data_7\ : std_logic;
signal n4445 : std_logic;
signal data_out_0_0 : std_logic;
signal data_out_frame2_12_3 : std_logic;
signal rand_data_29 : std_logic;
signal data_out_frame2_13_5 : std_logic;
signal \c0.data_out_5_1\ : std_logic;
signal \c0.n17043\ : std_logic;
signal \c0.n16949\ : std_logic;
signal data_out_8_7 : std_logic;
signal \c0.data_out_7__3__N_441\ : std_logic;
signal \c0.n10_adj_2276\ : std_logic;
signal \c0.data_out_9_3\ : std_logic;
signal \c0.n16981\ : std_logic;
signal \c0.n16969\ : std_logic;
signal \c0.n6_adj_2274\ : std_logic;
signal \c0.data_out_9_4\ : std_logic;
signal \c0.data_out_10_4\ : std_logic;
signal \c0.data_out_7_2\ : std_logic;
signal \c0.n17058\ : std_logic;
signal \c0.n17028\ : std_logic;
signal \c0.n17058_cascade_\ : std_logic;
signal \c0.n17094\ : std_logic;
signal \c0.n19_adj_2283\ : std_logic;
signal \c0.n21_adj_2284_cascade_\ : std_logic;
signal \c0.n20_adj_2282\ : std_logic;
signal \c0.data_out_9_7\ : std_logic;
signal \c0.n17007\ : std_logic;
signal \c0.n9505\ : std_logic;
signal \c0.n17076\ : std_logic;
signal data_out_8_0 : std_logic;
signal \c0.data_out_10_3\ : std_logic;
signal \c0.data_out_9_6\ : std_logic;
signal \c0.data_out_10_2\ : std_logic;
signal \c0.n16998\ : std_logic;
signal \c0.data_out_6_2\ : std_logic;
signal \c0.data_out_10_6\ : std_logic;
signal \data_out_10__7__N_110\ : std_logic;
signal rand_setpoint_21 : std_logic;
signal \c0.n17522\ : std_logic;
signal \UART_TRANSMITTER_state_1\ : std_logic;
signal \c0.data_out_6_5\ : std_logic;
signal n10055 : std_logic;
signal rand_setpoint_10 : std_logic;
signal \UART_TRANSMITTER_state_0\ : std_logic;
signal \c0.n17450\ : std_logic;
signal \c0.n17999\ : std_logic;
signal \c0.n8621\ : std_logic;
signal \c0.n18002\ : std_logic;
signal \c0.data_out_frame2_20_6\ : std_logic;
signal \c0.byte_transmit_counter2_2\ : std_logic;
signal \c0.n22_adj_2353\ : std_logic;
signal \c0.tx2.r_Tx_Data_6\ : std_logic;
signal \c0.n16915\ : std_logic;
signal \c0.n17082\ : std_logic;
signal \c0.n17118\ : std_logic;
signal \c0.n17019\ : std_logic;
signal \c0.n5_adj_2321\ : std_logic;
signal \c0.n18083\ : std_logic;
signal \c0.n6_adj_2290_cascade_\ : std_logic;
signal \c0.n18086\ : std_logic;
signal data_out_frame2_10_1 : std_logic;
signal data_out_frame2_12_0 : std_logic;
signal data_out_frame2_8_1 : std_logic;
signal data_out_frame2_14_3 : std_logic;
signal \c0.n9895_cascade_\ : std_logic;
signal data_out_frame2_15_1 : std_logic;
signal \c0.n26_adj_2314\ : std_logic;
signal \c0.n25_adj_2316\ : std_logic;
signal \c0.n23_adj_2318_cascade_\ : std_logic;
signal \c0.n24_adj_2315\ : std_logic;
signal rand_data_14 : std_logic;
signal data_out_frame2_17_6 : std_logic;
signal \c0.data_out_frame2_19_3\ : std_logic;
signal \c0.n17945_cascade_\ : std_logic;
signal data_out_frame2_16_3 : std_logic;
signal \c0.n17948\ : std_logic;
signal rand_data_30 : std_logic;
signal data_out_frame2_5_6 : std_logic;
signal rand_data_11 : std_logic;
signal data_out_frame2_17_3 : std_logic;
signal rand_data_8 : std_logic;
signal \c0.data_out_frame2_0_6\ : std_logic;
signal \c0.byte_transmit_counter2_1\ : std_logic;
signal \c0.byte_transmit_counter2_0\ : std_logic;
signal \c0.n17563\ : std_logic;
signal rand_data_6 : std_logic;
signal data_out_frame2_16_6 : std_logic;
signal rand_data_3 : std_logic;
signal data_out_frame2_18_3 : std_logic;
signal data_out_frame2_15_5 : std_logic;
signal data_out_frame2_11_0 : std_logic;
signal data_out_frame2_13_6 : std_logic;
signal \c0.n16923\ : std_logic;
signal data_out_frame2_13_1 : std_logic;
signal \c0.n9910\ : std_logic;
signal \c0.n9826\ : std_logic;
signal \c0.data_out_frame2_0_7\ : std_logic;
signal \c0.n9910_cascade_\ : std_logic;
signal \c0.n9843\ : std_logic;
signal data_out_frame2_14_1 : std_logic;
signal data_out_frame2_8_0 : std_logic;
signal data_out_frame2_15_0 : std_logic;
signal data_out_frame2_8_4 : std_logic;
signal \c0.n16_adj_2327\ : std_logic;
signal data_out_frame2_12_2 : std_logic;
signal \c0.n17_adj_2328_cascade_\ : std_logic;
signal \c0.n17010\ : std_logic;
signal \c0.data_out_frame2_19_1\ : std_logic;
signal data_out_frame2_15_7 : std_logic;
signal \c0.n16940\ : std_logic;
signal \c0.data_out_7_0\ : std_logic;
signal data_out_6_0 : std_logic;
signal byte_transmit_counter_2 : std_logic;
signal \c0.n5_adj_2265_cascade_\ : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal \c0.n18095\ : std_logic;
signal \c0.data_out_6__1__N_537\ : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal \c0.n17632\ : std_logic;
signal \c0.byte_transmit_counter2_4\ : std_logic;
signal \c0.n15_adj_2356\ : std_logic;
signal \c0.byte_transmit_counter2_3\ : std_logic;
signal \c0.n22_adj_2355\ : std_logic;
signal \c0.tx2.r_Tx_Data_4\ : std_logic;
signal \c0.tx2.n8737\ : std_logic;
signal rand_data_7 : std_logic;
signal n10197 : std_logic;
signal data_out_frame2_16_7 : std_logic;
signal \CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52613\,
            DIN => \N__52612\,
            DOUT => \N__52611\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__52613\,
            PADOUT => \N__52612\,
            PADIN => \N__52611\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__17170\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52604\,
            DIN => \N__52603\,
            DOUT => \N__52602\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__52604\,
            PADOUT => \N__52603\,
            PADIN => \N__52602\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__52595\,
            DIN => \N__52594\,
            DOUT => \N__52593\,
            PACKAGEPIN => PIN_2
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__52595\,
            PADOUT => \N__52594\,
            PADIN => \N__52593\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \c0.rx.r_Rx_Data_R\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__50505\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx2_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__52586\,
            DIN => \N__52585\,
            DOUT => \N__52584\,
            PACKAGEPIN => PIN_3
        );

    \tx2_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__52586\,
            PADOUT => \N__52585\,
            PADIN => \N__52584\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__28696\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__17155\
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__52577\,
            DIN => \N__52576\,
            DOUT => \N__52575\,
            PACKAGEPIN => PIN_1
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__52577\,
            PADOUT => \N__52576\,
            PADIN => \N__52575\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__20074\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20191\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52568\,
            DIN => \N__52567\,
            DOUT => \N__52566\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__52568\,
            PADOUT => \N__52567\,
            PADIN => \N__52566\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__13232\ : InMux
    port map (
            O => \N__52549\,
            I => \N__52545\
        );

    \I__13231\ : InMux
    port map (
            O => \N__52548\,
            I => \N__52541\
        );

    \I__13230\ : LocalMux
    port map (
            O => \N__52545\,
            I => \N__52538\
        );

    \I__13229\ : InMux
    port map (
            O => \N__52544\,
            I => \N__52535\
        );

    \I__13228\ : LocalMux
    port map (
            O => \N__52541\,
            I => \N__52532\
        );

    \I__13227\ : Span4Mux_h
    port map (
            O => \N__52538\,
            I => \N__52527\
        );

    \I__13226\ : LocalMux
    port map (
            O => \N__52535\,
            I => \N__52527\
        );

    \I__13225\ : Span4Mux_h
    port map (
            O => \N__52532\,
            I => \N__52524\
        );

    \I__13224\ : Span4Mux_h
    port map (
            O => \N__52527\,
            I => \N__52521\
        );

    \I__13223\ : Span4Mux_h
    port map (
            O => \N__52524\,
            I => \N__52518\
        );

    \I__13222\ : Odrv4
    port map (
            O => \N__52521\,
            I => \c0.data_out_7_0\
        );

    \I__13221\ : Odrv4
    port map (
            O => \N__52518\,
            I => \c0.data_out_7_0\
        );

    \I__13220\ : InMux
    port map (
            O => \N__52513\,
            I => \N__52508\
        );

    \I__13219\ : InMux
    port map (
            O => \N__52512\,
            I => \N__52505\
        );

    \I__13218\ : InMux
    port map (
            O => \N__52511\,
            I => \N__52502\
        );

    \I__13217\ : LocalMux
    port map (
            O => \N__52508\,
            I => \N__52499\
        );

    \I__13216\ : LocalMux
    port map (
            O => \N__52505\,
            I => \N__52494\
        );

    \I__13215\ : LocalMux
    port map (
            O => \N__52502\,
            I => \N__52491\
        );

    \I__13214\ : Span4Mux_h
    port map (
            O => \N__52499\,
            I => \N__52488\
        );

    \I__13213\ : InMux
    port map (
            O => \N__52498\,
            I => \N__52483\
        );

    \I__13212\ : InMux
    port map (
            O => \N__52497\,
            I => \N__52483\
        );

    \I__13211\ : Span4Mux_v
    port map (
            O => \N__52494\,
            I => \N__52480\
        );

    \I__13210\ : Span4Mux_h
    port map (
            O => \N__52491\,
            I => \N__52477\
        );

    \I__13209\ : Sp12to4
    port map (
            O => \N__52488\,
            I => \N__52474\
        );

    \I__13208\ : LocalMux
    port map (
            O => \N__52483\,
            I => data_out_6_0
        );

    \I__13207\ : Odrv4
    port map (
            O => \N__52480\,
            I => data_out_6_0
        );

    \I__13206\ : Odrv4
    port map (
            O => \N__52477\,
            I => data_out_6_0
        );

    \I__13205\ : Odrv12
    port map (
            O => \N__52474\,
            I => data_out_6_0
        );

    \I__13204\ : InMux
    port map (
            O => \N__52465\,
            I => \N__52448\
        );

    \I__13203\ : InMux
    port map (
            O => \N__52464\,
            I => \N__52445\
        );

    \I__13202\ : InMux
    port map (
            O => \N__52463\,
            I => \N__52438\
        );

    \I__13201\ : InMux
    port map (
            O => \N__52462\,
            I => \N__52438\
        );

    \I__13200\ : InMux
    port map (
            O => \N__52461\,
            I => \N__52438\
        );

    \I__13199\ : InMux
    port map (
            O => \N__52460\,
            I => \N__52434\
        );

    \I__13198\ : InMux
    port map (
            O => \N__52459\,
            I => \N__52429\
        );

    \I__13197\ : InMux
    port map (
            O => \N__52458\,
            I => \N__52429\
        );

    \I__13196\ : InMux
    port map (
            O => \N__52457\,
            I => \N__52426\
        );

    \I__13195\ : InMux
    port map (
            O => \N__52456\,
            I => \N__52419\
        );

    \I__13194\ : InMux
    port map (
            O => \N__52455\,
            I => \N__52419\
        );

    \I__13193\ : InMux
    port map (
            O => \N__52454\,
            I => \N__52419\
        );

    \I__13192\ : InMux
    port map (
            O => \N__52453\,
            I => \N__52416\
        );

    \I__13191\ : InMux
    port map (
            O => \N__52452\,
            I => \N__52410\
        );

    \I__13190\ : InMux
    port map (
            O => \N__52451\,
            I => \N__52410\
        );

    \I__13189\ : LocalMux
    port map (
            O => \N__52448\,
            I => \N__52399\
        );

    \I__13188\ : LocalMux
    port map (
            O => \N__52445\,
            I => \N__52399\
        );

    \I__13187\ : LocalMux
    port map (
            O => \N__52438\,
            I => \N__52396\
        );

    \I__13186\ : CascadeMux
    port map (
            O => \N__52437\,
            I => \N__52393\
        );

    \I__13185\ : LocalMux
    port map (
            O => \N__52434\,
            I => \N__52388\
        );

    \I__13184\ : LocalMux
    port map (
            O => \N__52429\,
            I => \N__52388\
        );

    \I__13183\ : LocalMux
    port map (
            O => \N__52426\,
            I => \N__52385\
        );

    \I__13182\ : LocalMux
    port map (
            O => \N__52419\,
            I => \N__52380\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__52416\,
            I => \N__52380\
        );

    \I__13180\ : InMux
    port map (
            O => \N__52415\,
            I => \N__52377\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__52410\,
            I => \N__52374\
        );

    \I__13178\ : InMux
    port map (
            O => \N__52409\,
            I => \N__52369\
        );

    \I__13177\ : InMux
    port map (
            O => \N__52408\,
            I => \N__52369\
        );

    \I__13176\ : InMux
    port map (
            O => \N__52407\,
            I => \N__52364\
        );

    \I__13175\ : InMux
    port map (
            O => \N__52406\,
            I => \N__52364\
        );

    \I__13174\ : InMux
    port map (
            O => \N__52405\,
            I => \N__52361\
        );

    \I__13173\ : InMux
    port map (
            O => \N__52404\,
            I => \N__52358\
        );

    \I__13172\ : Span4Mux_s2_v
    port map (
            O => \N__52399\,
            I => \N__52355\
        );

    \I__13171\ : Span4Mux_v
    port map (
            O => \N__52396\,
            I => \N__52352\
        );

    \I__13170\ : InMux
    port map (
            O => \N__52393\,
            I => \N__52348\
        );

    \I__13169\ : Span4Mux_s2_v
    port map (
            O => \N__52388\,
            I => \N__52345\
        );

    \I__13168\ : Span4Mux_v
    port map (
            O => \N__52385\,
            I => \N__52338\
        );

    \I__13167\ : Span4Mux_s2_v
    port map (
            O => \N__52380\,
            I => \N__52338\
        );

    \I__13166\ : LocalMux
    port map (
            O => \N__52377\,
            I => \N__52338\
        );

    \I__13165\ : Span4Mux_h
    port map (
            O => \N__52374\,
            I => \N__52335\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__52369\,
            I => \N__52322\
        );

    \I__13163\ : LocalMux
    port map (
            O => \N__52364\,
            I => \N__52322\
        );

    \I__13162\ : LocalMux
    port map (
            O => \N__52361\,
            I => \N__52322\
        );

    \I__13161\ : LocalMux
    port map (
            O => \N__52358\,
            I => \N__52322\
        );

    \I__13160\ : Sp12to4
    port map (
            O => \N__52355\,
            I => \N__52322\
        );

    \I__13159\ : Sp12to4
    port map (
            O => \N__52352\,
            I => \N__52322\
        );

    \I__13158\ : InMux
    port map (
            O => \N__52351\,
            I => \N__52319\
        );

    \I__13157\ : LocalMux
    port map (
            O => \N__52348\,
            I => byte_transmit_counter_2
        );

    \I__13156\ : Odrv4
    port map (
            O => \N__52345\,
            I => byte_transmit_counter_2
        );

    \I__13155\ : Odrv4
    port map (
            O => \N__52338\,
            I => byte_transmit_counter_2
        );

    \I__13154\ : Odrv4
    port map (
            O => \N__52335\,
            I => byte_transmit_counter_2
        );

    \I__13153\ : Odrv12
    port map (
            O => \N__52322\,
            I => byte_transmit_counter_2
        );

    \I__13152\ : LocalMux
    port map (
            O => \N__52319\,
            I => byte_transmit_counter_2
        );

    \I__13151\ : CascadeMux
    port map (
            O => \N__52306\,
            I => \c0.n5_adj_2265_cascade_\
        );

    \I__13150\ : InMux
    port map (
            O => \N__52303\,
            I => \N__52297\
        );

    \I__13149\ : InMux
    port map (
            O => \N__52302\,
            I => \N__52291\
        );

    \I__13148\ : InMux
    port map (
            O => \N__52301\,
            I => \N__52285\
        );

    \I__13147\ : CascadeMux
    port map (
            O => \N__52300\,
            I => \N__52282\
        );

    \I__13146\ : LocalMux
    port map (
            O => \N__52297\,
            I => \N__52279\
        );

    \I__13145\ : InMux
    port map (
            O => \N__52296\,
            I => \N__52272\
        );

    \I__13144\ : InMux
    port map (
            O => \N__52295\,
            I => \N__52272\
        );

    \I__13143\ : InMux
    port map (
            O => \N__52294\,
            I => \N__52272\
        );

    \I__13142\ : LocalMux
    port map (
            O => \N__52291\,
            I => \N__52269\
        );

    \I__13141\ : InMux
    port map (
            O => \N__52290\,
            I => \N__52266\
        );

    \I__13140\ : InMux
    port map (
            O => \N__52289\,
            I => \N__52261\
        );

    \I__13139\ : InMux
    port map (
            O => \N__52288\,
            I => \N__52258\
        );

    \I__13138\ : LocalMux
    port map (
            O => \N__52285\,
            I => \N__52254\
        );

    \I__13137\ : InMux
    port map (
            O => \N__52282\,
            I => \N__52251\
        );

    \I__13136\ : Span4Mux_h
    port map (
            O => \N__52279\,
            I => \N__52246\
        );

    \I__13135\ : LocalMux
    port map (
            O => \N__52272\,
            I => \N__52246\
        );

    \I__13134\ : Span4Mux_v
    port map (
            O => \N__52269\,
            I => \N__52243\
        );

    \I__13133\ : LocalMux
    port map (
            O => \N__52266\,
            I => \N__52240\
        );

    \I__13132\ : InMux
    port map (
            O => \N__52265\,
            I => \N__52237\
        );

    \I__13131\ : CascadeMux
    port map (
            O => \N__52264\,
            I => \N__52233\
        );

    \I__13130\ : LocalMux
    port map (
            O => \N__52261\,
            I => \N__52227\
        );

    \I__13129\ : LocalMux
    port map (
            O => \N__52258\,
            I => \N__52224\
        );

    \I__13128\ : InMux
    port map (
            O => \N__52257\,
            I => \N__52221\
        );

    \I__13127\ : Span4Mux_v
    port map (
            O => \N__52254\,
            I => \N__52216\
        );

    \I__13126\ : LocalMux
    port map (
            O => \N__52251\,
            I => \N__52216\
        );

    \I__13125\ : Span4Mux_v
    port map (
            O => \N__52246\,
            I => \N__52213\
        );

    \I__13124\ : Span4Mux_h
    port map (
            O => \N__52243\,
            I => \N__52208\
        );

    \I__13123\ : Span4Mux_v
    port map (
            O => \N__52240\,
            I => \N__52208\
        );

    \I__13122\ : LocalMux
    port map (
            O => \N__52237\,
            I => \N__52205\
        );

    \I__13121\ : CascadeMux
    port map (
            O => \N__52236\,
            I => \N__52202\
        );

    \I__13120\ : InMux
    port map (
            O => \N__52233\,
            I => \N__52197\
        );

    \I__13119\ : InMux
    port map (
            O => \N__52232\,
            I => \N__52197\
        );

    \I__13118\ : InMux
    port map (
            O => \N__52231\,
            I => \N__52192\
        );

    \I__13117\ : InMux
    port map (
            O => \N__52230\,
            I => \N__52192\
        );

    \I__13116\ : Span4Mux_v
    port map (
            O => \N__52227\,
            I => \N__52187\
        );

    \I__13115\ : Span4Mux_v
    port map (
            O => \N__52224\,
            I => \N__52187\
        );

    \I__13114\ : LocalMux
    port map (
            O => \N__52221\,
            I => \N__52176\
        );

    \I__13113\ : Sp12to4
    port map (
            O => \N__52216\,
            I => \N__52176\
        );

    \I__13112\ : Sp12to4
    port map (
            O => \N__52213\,
            I => \N__52176\
        );

    \I__13111\ : Sp12to4
    port map (
            O => \N__52208\,
            I => \N__52176\
        );

    \I__13110\ : Span12Mux_s4_v
    port map (
            O => \N__52205\,
            I => \N__52176\
        );

    \I__13109\ : InMux
    port map (
            O => \N__52202\,
            I => \N__52172\
        );

    \I__13108\ : LocalMux
    port map (
            O => \N__52197\,
            I => \N__52165\
        );

    \I__13107\ : LocalMux
    port map (
            O => \N__52192\,
            I => \N__52165\
        );

    \I__13106\ : Sp12to4
    port map (
            O => \N__52187\,
            I => \N__52165\
        );

    \I__13105\ : Span12Mux_h
    port map (
            O => \N__52176\,
            I => \N__52162\
        );

    \I__13104\ : InMux
    port map (
            O => \N__52175\,
            I => \N__52159\
        );

    \I__13103\ : LocalMux
    port map (
            O => \N__52172\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__13102\ : Odrv12
    port map (
            O => \N__52165\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__13101\ : Odrv12
    port map (
            O => \N__52162\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__13100\ : LocalMux
    port map (
            O => \N__52159\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__13099\ : InMux
    port map (
            O => \N__52150\,
            I => \N__52147\
        );

    \I__13098\ : LocalMux
    port map (
            O => \N__52147\,
            I => \N__52144\
        );

    \I__13097\ : Odrv12
    port map (
            O => \N__52144\,
            I => \c0.n18095\
        );

    \I__13096\ : InMux
    port map (
            O => \N__52141\,
            I => \N__52137\
        );

    \I__13095\ : InMux
    port map (
            O => \N__52140\,
            I => \N__52132\
        );

    \I__13094\ : LocalMux
    port map (
            O => \N__52137\,
            I => \N__52128\
        );

    \I__13093\ : InMux
    port map (
            O => \N__52136\,
            I => \N__52125\
        );

    \I__13092\ : InMux
    port map (
            O => \N__52135\,
            I => \N__52122\
        );

    \I__13091\ : LocalMux
    port map (
            O => \N__52132\,
            I => \N__52119\
        );

    \I__13090\ : InMux
    port map (
            O => \N__52131\,
            I => \N__52116\
        );

    \I__13089\ : Span4Mux_h
    port map (
            O => \N__52128\,
            I => \N__52113\
        );

    \I__13088\ : LocalMux
    port map (
            O => \N__52125\,
            I => \N__52110\
        );

    \I__13087\ : LocalMux
    port map (
            O => \N__52122\,
            I => \c0.data_out_6__1__N_537\
        );

    \I__13086\ : Odrv12
    port map (
            O => \N__52119\,
            I => \c0.data_out_6__1__N_537\
        );

    \I__13085\ : LocalMux
    port map (
            O => \N__52116\,
            I => \c0.data_out_6__1__N_537\
        );

    \I__13084\ : Odrv4
    port map (
            O => \N__52113\,
            I => \c0.data_out_6__1__N_537\
        );

    \I__13083\ : Odrv4
    port map (
            O => \N__52110\,
            I => \c0.data_out_6__1__N_537\
        );

    \I__13082\ : InMux
    port map (
            O => \N__52099\,
            I => \N__52093\
        );

    \I__13081\ : CascadeMux
    port map (
            O => \N__52098\,
            I => \N__52077\
        );

    \I__13080\ : CascadeMux
    port map (
            O => \N__52097\,
            I => \N__52073\
        );

    \I__13079\ : InMux
    port map (
            O => \N__52096\,
            I => \N__52067\
        );

    \I__13078\ : LocalMux
    port map (
            O => \N__52093\,
            I => \N__52057\
        );

    \I__13077\ : InMux
    port map (
            O => \N__52092\,
            I => \N__52045\
        );

    \I__13076\ : InMux
    port map (
            O => \N__52091\,
            I => \N__52045\
        );

    \I__13075\ : InMux
    port map (
            O => \N__52090\,
            I => \N__52045\
        );

    \I__13074\ : InMux
    port map (
            O => \N__52089\,
            I => \N__52045\
        );

    \I__13073\ : InMux
    port map (
            O => \N__52088\,
            I => \N__52035\
        );

    \I__13072\ : InMux
    port map (
            O => \N__52087\,
            I => \N__52030\
        );

    \I__13071\ : InMux
    port map (
            O => \N__52086\,
            I => \N__52030\
        );

    \I__13070\ : InMux
    port map (
            O => \N__52085\,
            I => \N__52025\
        );

    \I__13069\ : InMux
    port map (
            O => \N__52084\,
            I => \N__52025\
        );

    \I__13068\ : InMux
    port map (
            O => \N__52083\,
            I => \N__52022\
        );

    \I__13067\ : InMux
    port map (
            O => \N__52082\,
            I => \N__52019\
        );

    \I__13066\ : CascadeMux
    port map (
            O => \N__52081\,
            I => \N__52016\
        );

    \I__13065\ : InMux
    port map (
            O => \N__52080\,
            I => \N__52013\
        );

    \I__13064\ : InMux
    port map (
            O => \N__52077\,
            I => \N__52010\
        );

    \I__13063\ : InMux
    port map (
            O => \N__52076\,
            I => \N__52005\
        );

    \I__13062\ : InMux
    port map (
            O => \N__52073\,
            I => \N__52005\
        );

    \I__13061\ : InMux
    port map (
            O => \N__52072\,
            I => \N__51998\
        );

    \I__13060\ : InMux
    port map (
            O => \N__52071\,
            I => \N__51998\
        );

    \I__13059\ : InMux
    port map (
            O => \N__52070\,
            I => \N__51998\
        );

    \I__13058\ : LocalMux
    port map (
            O => \N__52067\,
            I => \N__51990\
        );

    \I__13057\ : InMux
    port map (
            O => \N__52066\,
            I => \N__51987\
        );

    \I__13056\ : InMux
    port map (
            O => \N__52065\,
            I => \N__51984\
        );

    \I__13055\ : InMux
    port map (
            O => \N__52064\,
            I => \N__51979\
        );

    \I__13054\ : InMux
    port map (
            O => \N__52063\,
            I => \N__51979\
        );

    \I__13053\ : InMux
    port map (
            O => \N__52062\,
            I => \N__51976\
        );

    \I__13052\ : InMux
    port map (
            O => \N__52061\,
            I => \N__51973\
        );

    \I__13051\ : InMux
    port map (
            O => \N__52060\,
            I => \N__51967\
        );

    \I__13050\ : Span4Mux_v
    port map (
            O => \N__52057\,
            I => \N__51964\
        );

    \I__13049\ : InMux
    port map (
            O => \N__52056\,
            I => \N__51957\
        );

    \I__13048\ : InMux
    port map (
            O => \N__52055\,
            I => \N__51957\
        );

    \I__13047\ : InMux
    port map (
            O => \N__52054\,
            I => \N__51957\
        );

    \I__13046\ : LocalMux
    port map (
            O => \N__52045\,
            I => \N__51954\
        );

    \I__13045\ : InMux
    port map (
            O => \N__52044\,
            I => \N__51951\
        );

    \I__13044\ : InMux
    port map (
            O => \N__52043\,
            I => \N__51948\
        );

    \I__13043\ : InMux
    port map (
            O => \N__52042\,
            I => \N__51939\
        );

    \I__13042\ : InMux
    port map (
            O => \N__52041\,
            I => \N__51939\
        );

    \I__13041\ : InMux
    port map (
            O => \N__52040\,
            I => \N__51939\
        );

    \I__13040\ : InMux
    port map (
            O => \N__52039\,
            I => \N__51939\
        );

    \I__13039\ : InMux
    port map (
            O => \N__52038\,
            I => \N__51935\
        );

    \I__13038\ : LocalMux
    port map (
            O => \N__52035\,
            I => \N__51924\
        );

    \I__13037\ : LocalMux
    port map (
            O => \N__52030\,
            I => \N__51924\
        );

    \I__13036\ : LocalMux
    port map (
            O => \N__52025\,
            I => \N__51924\
        );

    \I__13035\ : LocalMux
    port map (
            O => \N__52022\,
            I => \N__51924\
        );

    \I__13034\ : LocalMux
    port map (
            O => \N__52019\,
            I => \N__51924\
        );

    \I__13033\ : InMux
    port map (
            O => \N__52016\,
            I => \N__51921\
        );

    \I__13032\ : LocalMux
    port map (
            O => \N__52013\,
            I => \N__51918\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__52010\,
            I => \N__51913\
        );

    \I__13030\ : LocalMux
    port map (
            O => \N__52005\,
            I => \N__51913\
        );

    \I__13029\ : LocalMux
    port map (
            O => \N__51998\,
            I => \N__51910\
        );

    \I__13028\ : InMux
    port map (
            O => \N__51997\,
            I => \N__51905\
        );

    \I__13027\ : InMux
    port map (
            O => \N__51996\,
            I => \N__51905\
        );

    \I__13026\ : InMux
    port map (
            O => \N__51995\,
            I => \N__51898\
        );

    \I__13025\ : InMux
    port map (
            O => \N__51994\,
            I => \N__51898\
        );

    \I__13024\ : InMux
    port map (
            O => \N__51993\,
            I => \N__51898\
        );

    \I__13023\ : Span4Mux_v
    port map (
            O => \N__51990\,
            I => \N__51893\
        );

    \I__13022\ : LocalMux
    port map (
            O => \N__51987\,
            I => \N__51893\
        );

    \I__13021\ : LocalMux
    port map (
            O => \N__51984\,
            I => \N__51888\
        );

    \I__13020\ : LocalMux
    port map (
            O => \N__51979\,
            I => \N__51888\
        );

    \I__13019\ : LocalMux
    port map (
            O => \N__51976\,
            I => \N__51882\
        );

    \I__13018\ : LocalMux
    port map (
            O => \N__51973\,
            I => \N__51882\
        );

    \I__13017\ : InMux
    port map (
            O => \N__51972\,
            I => \N__51879\
        );

    \I__13016\ : InMux
    port map (
            O => \N__51971\,
            I => \N__51874\
        );

    \I__13015\ : InMux
    port map (
            O => \N__51970\,
            I => \N__51874\
        );

    \I__13014\ : LocalMux
    port map (
            O => \N__51967\,
            I => \N__51871\
        );

    \I__13013\ : Span4Mux_h
    port map (
            O => \N__51964\,
            I => \N__51864\
        );

    \I__13012\ : LocalMux
    port map (
            O => \N__51957\,
            I => \N__51864\
        );

    \I__13011\ : Span4Mux_v
    port map (
            O => \N__51954\,
            I => \N__51864\
        );

    \I__13010\ : LocalMux
    port map (
            O => \N__51951\,
            I => \N__51857\
        );

    \I__13009\ : LocalMux
    port map (
            O => \N__51948\,
            I => \N__51857\
        );

    \I__13008\ : LocalMux
    port map (
            O => \N__51939\,
            I => \N__51857\
        );

    \I__13007\ : InMux
    port map (
            O => \N__51938\,
            I => \N__51854\
        );

    \I__13006\ : LocalMux
    port map (
            O => \N__51935\,
            I => \N__51851\
        );

    \I__13005\ : Span4Mux_v
    port map (
            O => \N__51924\,
            I => \N__51846\
        );

    \I__13004\ : LocalMux
    port map (
            O => \N__51921\,
            I => \N__51846\
        );

    \I__13003\ : Span12Mux_h
    port map (
            O => \N__51918\,
            I => \N__51843\
        );

    \I__13002\ : Span4Mux_v
    port map (
            O => \N__51913\,
            I => \N__51836\
        );

    \I__13001\ : Span4Mux_h
    port map (
            O => \N__51910\,
            I => \N__51836\
        );

    \I__13000\ : LocalMux
    port map (
            O => \N__51905\,
            I => \N__51836\
        );

    \I__12999\ : LocalMux
    port map (
            O => \N__51898\,
            I => \N__51829\
        );

    \I__12998\ : Span4Mux_h
    port map (
            O => \N__51893\,
            I => \N__51829\
        );

    \I__12997\ : Span4Mux_v
    port map (
            O => \N__51888\,
            I => \N__51829\
        );

    \I__12996\ : CascadeMux
    port map (
            O => \N__51887\,
            I => \N__51826\
        );

    \I__12995\ : Span4Mux_h
    port map (
            O => \N__51882\,
            I => \N__51823\
        );

    \I__12994\ : LocalMux
    port map (
            O => \N__51879\,
            I => \N__51812\
        );

    \I__12993\ : LocalMux
    port map (
            O => \N__51874\,
            I => \N__51812\
        );

    \I__12992\ : Span4Mux_s1_v
    port map (
            O => \N__51871\,
            I => \N__51812\
        );

    \I__12991\ : Span4Mux_h
    port map (
            O => \N__51864\,
            I => \N__51812\
        );

    \I__12990\ : Span4Mux_v
    port map (
            O => \N__51857\,
            I => \N__51812\
        );

    \I__12989\ : LocalMux
    port map (
            O => \N__51854\,
            I => \N__51809\
        );

    \I__12988\ : Span12Mux_h
    port map (
            O => \N__51851\,
            I => \N__51802\
        );

    \I__12987\ : Sp12to4
    port map (
            O => \N__51846\,
            I => \N__51802\
        );

    \I__12986\ : Span12Mux_v
    port map (
            O => \N__51843\,
            I => \N__51802\
        );

    \I__12985\ : Span4Mux_h
    port map (
            O => \N__51836\,
            I => \N__51797\
        );

    \I__12984\ : Span4Mux_h
    port map (
            O => \N__51829\,
            I => \N__51797\
        );

    \I__12983\ : InMux
    port map (
            O => \N__51826\,
            I => \N__51794\
        );

    \I__12982\ : Odrv4
    port map (
            O => \N__51823\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__12981\ : Odrv4
    port map (
            O => \N__51812\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__12980\ : Odrv12
    port map (
            O => \N__51809\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__12979\ : Odrv12
    port map (
            O => \N__51802\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__12978\ : Odrv4
    port map (
            O => \N__51797\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__12977\ : LocalMux
    port map (
            O => \N__51794\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__12976\ : InMux
    port map (
            O => \N__51781\,
            I => \N__51778\
        );

    \I__12975\ : LocalMux
    port map (
            O => \N__51778\,
            I => \c0.n17632\
        );

    \I__12974\ : CascadeMux
    port map (
            O => \N__51775\,
            I => \N__51771\
        );

    \I__12973\ : CascadeMux
    port map (
            O => \N__51774\,
            I => \N__51767\
        );

    \I__12972\ : InMux
    port map (
            O => \N__51771\,
            I => \N__51764\
        );

    \I__12971\ : InMux
    port map (
            O => \N__51770\,
            I => \N__51758\
        );

    \I__12970\ : InMux
    port map (
            O => \N__51767\,
            I => \N__51755\
        );

    \I__12969\ : LocalMux
    port map (
            O => \N__51764\,
            I => \N__51752\
        );

    \I__12968\ : InMux
    port map (
            O => \N__51763\,
            I => \N__51749\
        );

    \I__12967\ : InMux
    port map (
            O => \N__51762\,
            I => \N__51746\
        );

    \I__12966\ : InMux
    port map (
            O => \N__51761\,
            I => \N__51743\
        );

    \I__12965\ : LocalMux
    port map (
            O => \N__51758\,
            I => \N__51740\
        );

    \I__12964\ : LocalMux
    port map (
            O => \N__51755\,
            I => \N__51733\
        );

    \I__12963\ : Span4Mux_v
    port map (
            O => \N__51752\,
            I => \N__51733\
        );

    \I__12962\ : LocalMux
    port map (
            O => \N__51749\,
            I => \N__51730\
        );

    \I__12961\ : LocalMux
    port map (
            O => \N__51746\,
            I => \N__51727\
        );

    \I__12960\ : LocalMux
    port map (
            O => \N__51743\,
            I => \N__51724\
        );

    \I__12959\ : Span4Mux_h
    port map (
            O => \N__51740\,
            I => \N__51721\
        );

    \I__12958\ : InMux
    port map (
            O => \N__51739\,
            I => \N__51718\
        );

    \I__12957\ : InMux
    port map (
            O => \N__51738\,
            I => \N__51715\
        );

    \I__12956\ : Span4Mux_v
    port map (
            O => \N__51733\,
            I => \N__51711\
        );

    \I__12955\ : Span4Mux_v
    port map (
            O => \N__51730\,
            I => \N__51702\
        );

    \I__12954\ : Span4Mux_v
    port map (
            O => \N__51727\,
            I => \N__51702\
        );

    \I__12953\ : Span4Mux_v
    port map (
            O => \N__51724\,
            I => \N__51702\
        );

    \I__12952\ : Span4Mux_h
    port map (
            O => \N__51721\,
            I => \N__51702\
        );

    \I__12951\ : LocalMux
    port map (
            O => \N__51718\,
            I => \N__51698\
        );

    \I__12950\ : LocalMux
    port map (
            O => \N__51715\,
            I => \N__51695\
        );

    \I__12949\ : InMux
    port map (
            O => \N__51714\,
            I => \N__51692\
        );

    \I__12948\ : Span4Mux_h
    port map (
            O => \N__51711\,
            I => \N__51689\
        );

    \I__12947\ : Span4Mux_v
    port map (
            O => \N__51702\,
            I => \N__51686\
        );

    \I__12946\ : InMux
    port map (
            O => \N__51701\,
            I => \N__51683\
        );

    \I__12945\ : Odrv4
    port map (
            O => \N__51698\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12944\ : Odrv4
    port map (
            O => \N__51695\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__51692\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12942\ : Odrv4
    port map (
            O => \N__51689\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12941\ : Odrv4
    port map (
            O => \N__51686\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12940\ : LocalMux
    port map (
            O => \N__51683\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12939\ : InMux
    port map (
            O => \N__51670\,
            I => \N__51667\
        );

    \I__12938\ : LocalMux
    port map (
            O => \N__51667\,
            I => \N__51664\
        );

    \I__12937\ : Span4Mux_h
    port map (
            O => \N__51664\,
            I => \N__51661\
        );

    \I__12936\ : Span4Mux_h
    port map (
            O => \N__51661\,
            I => \N__51658\
        );

    \I__12935\ : Odrv4
    port map (
            O => \N__51658\,
            I => \c0.n15_adj_2356\
        );

    \I__12934\ : CascadeMux
    port map (
            O => \N__51655\,
            I => \N__51652\
        );

    \I__12933\ : InMux
    port map (
            O => \N__51652\,
            I => \N__51648\
        );

    \I__12932\ : InMux
    port map (
            O => \N__51651\,
            I => \N__51640\
        );

    \I__12931\ : LocalMux
    port map (
            O => \N__51648\,
            I => \N__51637\
        );

    \I__12930\ : InMux
    port map (
            O => \N__51647\,
            I => \N__51634\
        );

    \I__12929\ : InMux
    port map (
            O => \N__51646\,
            I => \N__51626\
        );

    \I__12928\ : InMux
    port map (
            O => \N__51645\,
            I => \N__51626\
        );

    \I__12927\ : InMux
    port map (
            O => \N__51644\,
            I => \N__51623\
        );

    \I__12926\ : InMux
    port map (
            O => \N__51643\,
            I => \N__51610\
        );

    \I__12925\ : LocalMux
    port map (
            O => \N__51640\,
            I => \N__51601\
        );

    \I__12924\ : Span4Mux_v
    port map (
            O => \N__51637\,
            I => \N__51601\
        );

    \I__12923\ : LocalMux
    port map (
            O => \N__51634\,
            I => \N__51601\
        );

    \I__12922\ : InMux
    port map (
            O => \N__51633\,
            I => \N__51594\
        );

    \I__12921\ : InMux
    port map (
            O => \N__51632\,
            I => \N__51594\
        );

    \I__12920\ : InMux
    port map (
            O => \N__51631\,
            I => \N__51594\
        );

    \I__12919\ : LocalMux
    port map (
            O => \N__51626\,
            I => \N__51589\
        );

    \I__12918\ : LocalMux
    port map (
            O => \N__51623\,
            I => \N__51589\
        );

    \I__12917\ : InMux
    port map (
            O => \N__51622\,
            I => \N__51586\
        );

    \I__12916\ : InMux
    port map (
            O => \N__51621\,
            I => \N__51583\
        );

    \I__12915\ : InMux
    port map (
            O => \N__51620\,
            I => \N__51580\
        );

    \I__12914\ : InMux
    port map (
            O => \N__51619\,
            I => \N__51577\
        );

    \I__12913\ : InMux
    port map (
            O => \N__51618\,
            I => \N__51571\
        );

    \I__12912\ : InMux
    port map (
            O => \N__51617\,
            I => \N__51571\
        );

    \I__12911\ : InMux
    port map (
            O => \N__51616\,
            I => \N__51564\
        );

    \I__12910\ : InMux
    port map (
            O => \N__51615\,
            I => \N__51564\
        );

    \I__12909\ : InMux
    port map (
            O => \N__51614\,
            I => \N__51564\
        );

    \I__12908\ : InMux
    port map (
            O => \N__51613\,
            I => \N__51561\
        );

    \I__12907\ : LocalMux
    port map (
            O => \N__51610\,
            I => \N__51558\
        );

    \I__12906\ : InMux
    port map (
            O => \N__51609\,
            I => \N__51553\
        );

    \I__12905\ : InMux
    port map (
            O => \N__51608\,
            I => \N__51553\
        );

    \I__12904\ : Span4Mux_v
    port map (
            O => \N__51601\,
            I => \N__51550\
        );

    \I__12903\ : LocalMux
    port map (
            O => \N__51594\,
            I => \N__51545\
        );

    \I__12902\ : Span4Mux_v
    port map (
            O => \N__51589\,
            I => \N__51545\
        );

    \I__12901\ : LocalMux
    port map (
            O => \N__51586\,
            I => \N__51536\
        );

    \I__12900\ : LocalMux
    port map (
            O => \N__51583\,
            I => \N__51536\
        );

    \I__12899\ : LocalMux
    port map (
            O => \N__51580\,
            I => \N__51536\
        );

    \I__12898\ : LocalMux
    port map (
            O => \N__51577\,
            I => \N__51536\
        );

    \I__12897\ : InMux
    port map (
            O => \N__51576\,
            I => \N__51532\
        );

    \I__12896\ : LocalMux
    port map (
            O => \N__51571\,
            I => \N__51525\
        );

    \I__12895\ : LocalMux
    port map (
            O => \N__51564\,
            I => \N__51525\
        );

    \I__12894\ : LocalMux
    port map (
            O => \N__51561\,
            I => \N__51525\
        );

    \I__12893\ : Span4Mux_h
    port map (
            O => \N__51558\,
            I => \N__51522\
        );

    \I__12892\ : LocalMux
    port map (
            O => \N__51553\,
            I => \N__51515\
        );

    \I__12891\ : Span4Mux_h
    port map (
            O => \N__51550\,
            I => \N__51515\
        );

    \I__12890\ : Span4Mux_v
    port map (
            O => \N__51545\,
            I => \N__51515\
        );

    \I__12889\ : Span12Mux_v
    port map (
            O => \N__51536\,
            I => \N__51512\
        );

    \I__12888\ : InMux
    port map (
            O => \N__51535\,
            I => \N__51509\
        );

    \I__12887\ : LocalMux
    port map (
            O => \N__51532\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12886\ : Odrv12
    port map (
            O => \N__51525\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12885\ : Odrv4
    port map (
            O => \N__51522\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12884\ : Odrv4
    port map (
            O => \N__51515\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12883\ : Odrv12
    port map (
            O => \N__51512\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12882\ : LocalMux
    port map (
            O => \N__51509\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12881\ : InMux
    port map (
            O => \N__51496\,
            I => \N__51493\
        );

    \I__12880\ : LocalMux
    port map (
            O => \N__51493\,
            I => \N__51490\
        );

    \I__12879\ : Span4Mux_v
    port map (
            O => \N__51490\,
            I => \N__51487\
        );

    \I__12878\ : Odrv4
    port map (
            O => \N__51487\,
            I => \c0.n22_adj_2355\
        );

    \I__12877\ : CascadeMux
    port map (
            O => \N__51484\,
            I => \N__51481\
        );

    \I__12876\ : InMux
    port map (
            O => \N__51481\,
            I => \N__51478\
        );

    \I__12875\ : LocalMux
    port map (
            O => \N__51478\,
            I => \N__51475\
        );

    \I__12874\ : Span4Mux_h
    port map (
            O => \N__51475\,
            I => \N__51472\
        );

    \I__12873\ : Span4Mux_h
    port map (
            O => \N__51472\,
            I => \N__51469\
        );

    \I__12872\ : Span4Mux_v
    port map (
            O => \N__51469\,
            I => \N__51466\
        );

    \I__12871\ : Odrv4
    port map (
            O => \N__51466\,
            I => \c0.tx2.r_Tx_Data_4\
        );

    \I__12870\ : CEMux
    port map (
            O => \N__51463\,
            I => \N__51459\
        );

    \I__12869\ : CEMux
    port map (
            O => \N__51462\,
            I => \N__51456\
        );

    \I__12868\ : LocalMux
    port map (
            O => \N__51459\,
            I => \N__51453\
        );

    \I__12867\ : LocalMux
    port map (
            O => \N__51456\,
            I => \N__51448\
        );

    \I__12866\ : Span4Mux_v
    port map (
            O => \N__51453\,
            I => \N__51443\
        );

    \I__12865\ : CEMux
    port map (
            O => \N__51452\,
            I => \N__51440\
        );

    \I__12864\ : CEMux
    port map (
            O => \N__51451\,
            I => \N__51437\
        );

    \I__12863\ : Span4Mux_v
    port map (
            O => \N__51448\,
            I => \N__51434\
        );

    \I__12862\ : CEMux
    port map (
            O => \N__51447\,
            I => \N__51431\
        );

    \I__12861\ : CEMux
    port map (
            O => \N__51446\,
            I => \N__51428\
        );

    \I__12860\ : Span4Mux_h
    port map (
            O => \N__51443\,
            I => \N__51423\
        );

    \I__12859\ : LocalMux
    port map (
            O => \N__51440\,
            I => \N__51423\
        );

    \I__12858\ : LocalMux
    port map (
            O => \N__51437\,
            I => \N__51420\
        );

    \I__12857\ : Span4Mux_h
    port map (
            O => \N__51434\,
            I => \N__51415\
        );

    \I__12856\ : LocalMux
    port map (
            O => \N__51431\,
            I => \N__51415\
        );

    \I__12855\ : LocalMux
    port map (
            O => \N__51428\,
            I => \N__51412\
        );

    \I__12854\ : Span4Mux_h
    port map (
            O => \N__51423\,
            I => \N__51408\
        );

    \I__12853\ : Span4Mux_v
    port map (
            O => \N__51420\,
            I => \N__51405\
        );

    \I__12852\ : Span4Mux_v
    port map (
            O => \N__51415\,
            I => \N__51401\
        );

    \I__12851\ : Span4Mux_v
    port map (
            O => \N__51412\,
            I => \N__51398\
        );

    \I__12850\ : CEMux
    port map (
            O => \N__51411\,
            I => \N__51395\
        );

    \I__12849\ : Span4Mux_h
    port map (
            O => \N__51408\,
            I => \N__51390\
        );

    \I__12848\ : Span4Mux_h
    port map (
            O => \N__51405\,
            I => \N__51390\
        );

    \I__12847\ : CEMux
    port map (
            O => \N__51404\,
            I => \N__51387\
        );

    \I__12846\ : Sp12to4
    port map (
            O => \N__51401\,
            I => \N__51384\
        );

    \I__12845\ : Span4Mux_h
    port map (
            O => \N__51398\,
            I => \N__51381\
        );

    \I__12844\ : LocalMux
    port map (
            O => \N__51395\,
            I => \N__51378\
        );

    \I__12843\ : Span4Mux_v
    port map (
            O => \N__51390\,
            I => \N__51373\
        );

    \I__12842\ : LocalMux
    port map (
            O => \N__51387\,
            I => \N__51373\
        );

    \I__12841\ : Span12Mux_h
    port map (
            O => \N__51384\,
            I => \N__51370\
        );

    \I__12840\ : Span4Mux_h
    port map (
            O => \N__51381\,
            I => \N__51365\
        );

    \I__12839\ : Span4Mux_h
    port map (
            O => \N__51378\,
            I => \N__51365\
        );

    \I__12838\ : Span4Mux_h
    port map (
            O => \N__51373\,
            I => \N__51362\
        );

    \I__12837\ : Span12Mux_v
    port map (
            O => \N__51370\,
            I => \N__51359\
        );

    \I__12836\ : Span4Mux_h
    port map (
            O => \N__51365\,
            I => \N__51356\
        );

    \I__12835\ : Span4Mux_h
    port map (
            O => \N__51362\,
            I => \N__51353\
        );

    \I__12834\ : Odrv12
    port map (
            O => \N__51359\,
            I => \c0.tx2.n8737\
        );

    \I__12833\ : Odrv4
    port map (
            O => \N__51356\,
            I => \c0.tx2.n8737\
        );

    \I__12832\ : Odrv4
    port map (
            O => \N__51353\,
            I => \c0.tx2.n8737\
        );

    \I__12831\ : InMux
    port map (
            O => \N__51346\,
            I => \N__51343\
        );

    \I__12830\ : LocalMux
    port map (
            O => \N__51343\,
            I => \N__51340\
        );

    \I__12829\ : Span4Mux_v
    port map (
            O => \N__51340\,
            I => \N__51335\
        );

    \I__12828\ : InMux
    port map (
            O => \N__51339\,
            I => \N__51332\
        );

    \I__12827\ : InMux
    port map (
            O => \N__51338\,
            I => \N__51329\
        );

    \I__12826\ : Span4Mux_h
    port map (
            O => \N__51335\,
            I => \N__51322\
        );

    \I__12825\ : LocalMux
    port map (
            O => \N__51332\,
            I => \N__51322\
        );

    \I__12824\ : LocalMux
    port map (
            O => \N__51329\,
            I => \N__51319\
        );

    \I__12823\ : InMux
    port map (
            O => \N__51328\,
            I => \N__51316\
        );

    \I__12822\ : CascadeMux
    port map (
            O => \N__51327\,
            I => \N__51313\
        );

    \I__12821\ : Span4Mux_v
    port map (
            O => \N__51322\,
            I => \N__51310\
        );

    \I__12820\ : Span4Mux_h
    port map (
            O => \N__51319\,
            I => \N__51305\
        );

    \I__12819\ : LocalMux
    port map (
            O => \N__51316\,
            I => \N__51305\
        );

    \I__12818\ : InMux
    port map (
            O => \N__51313\,
            I => \N__51301\
        );

    \I__12817\ : Span4Mux_h
    port map (
            O => \N__51310\,
            I => \N__51298\
        );

    \I__12816\ : Span4Mux_h
    port map (
            O => \N__51305\,
            I => \N__51295\
        );

    \I__12815\ : InMux
    port map (
            O => \N__51304\,
            I => \N__51292\
        );

    \I__12814\ : LocalMux
    port map (
            O => \N__51301\,
            I => \N__51289\
        );

    \I__12813\ : Odrv4
    port map (
            O => \N__51298\,
            I => rand_data_7
        );

    \I__12812\ : Odrv4
    port map (
            O => \N__51295\,
            I => rand_data_7
        );

    \I__12811\ : LocalMux
    port map (
            O => \N__51292\,
            I => rand_data_7
        );

    \I__12810\ : Odrv12
    port map (
            O => \N__51289\,
            I => rand_data_7
        );

    \I__12809\ : InMux
    port map (
            O => \N__51280\,
            I => \N__51266\
        );

    \I__12808\ : InMux
    port map (
            O => \N__51279\,
            I => \N__51266\
        );

    \I__12807\ : InMux
    port map (
            O => \N__51278\,
            I => \N__51261\
        );

    \I__12806\ : InMux
    port map (
            O => \N__51277\,
            I => \N__51261\
        );

    \I__12805\ : InMux
    port map (
            O => \N__51276\,
            I => \N__51256\
        );

    \I__12804\ : InMux
    port map (
            O => \N__51275\,
            I => \N__51256\
        );

    \I__12803\ : InMux
    port map (
            O => \N__51274\,
            I => \N__51251\
        );

    \I__12802\ : InMux
    port map (
            O => \N__51273\,
            I => \N__51251\
        );

    \I__12801\ : InMux
    port map (
            O => \N__51272\,
            I => \N__51240\
        );

    \I__12800\ : InMux
    port map (
            O => \N__51271\,
            I => \N__51237\
        );

    \I__12799\ : LocalMux
    port map (
            O => \N__51266\,
            I => \N__51228\
        );

    \I__12798\ : LocalMux
    port map (
            O => \N__51261\,
            I => \N__51228\
        );

    \I__12797\ : LocalMux
    port map (
            O => \N__51256\,
            I => \N__51228\
        );

    \I__12796\ : LocalMux
    port map (
            O => \N__51251\,
            I => \N__51228\
        );

    \I__12795\ : InMux
    port map (
            O => \N__51250\,
            I => \N__51225\
        );

    \I__12794\ : InMux
    port map (
            O => \N__51249\,
            I => \N__51174\
        );

    \I__12793\ : CascadeMux
    port map (
            O => \N__51248\,
            I => \N__51171\
        );

    \I__12792\ : CascadeMux
    port map (
            O => \N__51247\,
            I => \N__51165\
        );

    \I__12791\ : CascadeMux
    port map (
            O => \N__51246\,
            I => \N__51162\
        );

    \I__12790\ : InMux
    port map (
            O => \N__51245\,
            I => \N__51154\
        );

    \I__12789\ : InMux
    port map (
            O => \N__51244\,
            I => \N__51154\
        );

    \I__12788\ : InMux
    port map (
            O => \N__51243\,
            I => \N__51154\
        );

    \I__12787\ : LocalMux
    port map (
            O => \N__51240\,
            I => \N__51151\
        );

    \I__12786\ : LocalMux
    port map (
            O => \N__51237\,
            I => \N__51148\
        );

    \I__12785\ : Span4Mux_v
    port map (
            O => \N__51228\,
            I => \N__51142\
        );

    \I__12784\ : LocalMux
    port map (
            O => \N__51225\,
            I => \N__51142\
        );

    \I__12783\ : InMux
    port map (
            O => \N__51224\,
            I => \N__51139\
        );

    \I__12782\ : InMux
    port map (
            O => \N__51223\,
            I => \N__51132\
        );

    \I__12781\ : InMux
    port map (
            O => \N__51222\,
            I => \N__51117\
        );

    \I__12780\ : InMux
    port map (
            O => \N__51221\,
            I => \N__51117\
        );

    \I__12779\ : InMux
    port map (
            O => \N__51220\,
            I => \N__51117\
        );

    \I__12778\ : InMux
    port map (
            O => \N__51219\,
            I => \N__51117\
        );

    \I__12777\ : InMux
    port map (
            O => \N__51218\,
            I => \N__51112\
        );

    \I__12776\ : InMux
    port map (
            O => \N__51217\,
            I => \N__51112\
        );

    \I__12775\ : CEMux
    port map (
            O => \N__51216\,
            I => \N__51109\
        );

    \I__12774\ : CEMux
    port map (
            O => \N__51215\,
            I => \N__51106\
        );

    \I__12773\ : InMux
    port map (
            O => \N__51214\,
            I => \N__51097\
        );

    \I__12772\ : InMux
    port map (
            O => \N__51213\,
            I => \N__51097\
        );

    \I__12771\ : InMux
    port map (
            O => \N__51212\,
            I => \N__51094\
        );

    \I__12770\ : InMux
    port map (
            O => \N__51211\,
            I => \N__51089\
        );

    \I__12769\ : InMux
    port map (
            O => \N__51210\,
            I => \N__51089\
        );

    \I__12768\ : InMux
    port map (
            O => \N__51209\,
            I => \N__51084\
        );

    \I__12767\ : InMux
    port map (
            O => \N__51208\,
            I => \N__51084\
        );

    \I__12766\ : InMux
    port map (
            O => \N__51207\,
            I => \N__51081\
        );

    \I__12765\ : InMux
    port map (
            O => \N__51206\,
            I => \N__51074\
        );

    \I__12764\ : InMux
    port map (
            O => \N__51205\,
            I => \N__51074\
        );

    \I__12763\ : InMux
    port map (
            O => \N__51204\,
            I => \N__51074\
        );

    \I__12762\ : InMux
    port map (
            O => \N__51203\,
            I => \N__51066\
        );

    \I__12761\ : InMux
    port map (
            O => \N__51202\,
            I => \N__51066\
        );

    \I__12760\ : InMux
    port map (
            O => \N__51201\,
            I => \N__51066\
        );

    \I__12759\ : InMux
    port map (
            O => \N__51200\,
            I => \N__51061\
        );

    \I__12758\ : InMux
    port map (
            O => \N__51199\,
            I => \N__51061\
        );

    \I__12757\ : InMux
    port map (
            O => \N__51198\,
            I => \N__51054\
        );

    \I__12756\ : InMux
    port map (
            O => \N__51197\,
            I => \N__51054\
        );

    \I__12755\ : InMux
    port map (
            O => \N__51196\,
            I => \N__51054\
        );

    \I__12754\ : InMux
    port map (
            O => \N__51195\,
            I => \N__51043\
        );

    \I__12753\ : InMux
    port map (
            O => \N__51194\,
            I => \N__51043\
        );

    \I__12752\ : InMux
    port map (
            O => \N__51193\,
            I => \N__51043\
        );

    \I__12751\ : InMux
    port map (
            O => \N__51192\,
            I => \N__51043\
        );

    \I__12750\ : InMux
    port map (
            O => \N__51191\,
            I => \N__51043\
        );

    \I__12749\ : InMux
    port map (
            O => \N__51190\,
            I => \N__51040\
        );

    \I__12748\ : InMux
    port map (
            O => \N__51189\,
            I => \N__51033\
        );

    \I__12747\ : InMux
    port map (
            O => \N__51188\,
            I => \N__51033\
        );

    \I__12746\ : InMux
    port map (
            O => \N__51187\,
            I => \N__51033\
        );

    \I__12745\ : InMux
    port map (
            O => \N__51186\,
            I => \N__51030\
        );

    \I__12744\ : CEMux
    port map (
            O => \N__51185\,
            I => \N__51027\
        );

    \I__12743\ : CEMux
    port map (
            O => \N__51184\,
            I => \N__51024\
        );

    \I__12742\ : InMux
    port map (
            O => \N__51183\,
            I => \N__51021\
        );

    \I__12741\ : CEMux
    port map (
            O => \N__51182\,
            I => \N__51018\
        );

    \I__12740\ : CEMux
    port map (
            O => \N__51181\,
            I => \N__51015\
        );

    \I__12739\ : InMux
    port map (
            O => \N__51180\,
            I => \N__51012\
        );

    \I__12738\ : InMux
    port map (
            O => \N__51179\,
            I => \N__51005\
        );

    \I__12737\ : InMux
    port map (
            O => \N__51178\,
            I => \N__51005\
        );

    \I__12736\ : InMux
    port map (
            O => \N__51177\,
            I => \N__51005\
        );

    \I__12735\ : LocalMux
    port map (
            O => \N__51174\,
            I => \N__51002\
        );

    \I__12734\ : InMux
    port map (
            O => \N__51171\,
            I => \N__50996\
        );

    \I__12733\ : InMux
    port map (
            O => \N__51170\,
            I => \N__50996\
        );

    \I__12732\ : CEMux
    port map (
            O => \N__51169\,
            I => \N__50992\
        );

    \I__12731\ : CEMux
    port map (
            O => \N__51168\,
            I => \N__50989\
        );

    \I__12730\ : InMux
    port map (
            O => \N__51165\,
            I => \N__50982\
        );

    \I__12729\ : InMux
    port map (
            O => \N__51162\,
            I => \N__50982\
        );

    \I__12728\ : InMux
    port map (
            O => \N__51161\,
            I => \N__50982\
        );

    \I__12727\ : LocalMux
    port map (
            O => \N__51154\,
            I => \N__50977\
        );

    \I__12726\ : Span4Mux_v
    port map (
            O => \N__51151\,
            I => \N__50977\
        );

    \I__12725\ : Span4Mux_h
    port map (
            O => \N__51148\,
            I => \N__50974\
        );

    \I__12724\ : InMux
    port map (
            O => \N__51147\,
            I => \N__50971\
        );

    \I__12723\ : Span4Mux_v
    port map (
            O => \N__51142\,
            I => \N__50966\
        );

    \I__12722\ : LocalMux
    port map (
            O => \N__51139\,
            I => \N__50966\
        );

    \I__12721\ : InMux
    port map (
            O => \N__51138\,
            I => \N__50956\
        );

    \I__12720\ : InMux
    port map (
            O => \N__51137\,
            I => \N__50956\
        );

    \I__12719\ : InMux
    port map (
            O => \N__51136\,
            I => \N__50956\
        );

    \I__12718\ : InMux
    port map (
            O => \N__51135\,
            I => \N__50956\
        );

    \I__12717\ : LocalMux
    port map (
            O => \N__51132\,
            I => \N__50953\
        );

    \I__12716\ : InMux
    port map (
            O => \N__51131\,
            I => \N__50908\
        );

    \I__12715\ : InMux
    port map (
            O => \N__51130\,
            I => \N__50908\
        );

    \I__12714\ : InMux
    port map (
            O => \N__51129\,
            I => \N__50908\
        );

    \I__12713\ : InMux
    port map (
            O => \N__51128\,
            I => \N__50908\
        );

    \I__12712\ : InMux
    port map (
            O => \N__51127\,
            I => \N__50908\
        );

    \I__12711\ : InMux
    port map (
            O => \N__51126\,
            I => \N__50908\
        );

    \I__12710\ : LocalMux
    port map (
            O => \N__51117\,
            I => \N__50901\
        );

    \I__12709\ : LocalMux
    port map (
            O => \N__51112\,
            I => \N__50901\
        );

    \I__12708\ : LocalMux
    port map (
            O => \N__51109\,
            I => \N__50901\
        );

    \I__12707\ : LocalMux
    port map (
            O => \N__51106\,
            I => \N__50898\
        );

    \I__12706\ : InMux
    port map (
            O => \N__51105\,
            I => \N__50889\
        );

    \I__12705\ : InMux
    port map (
            O => \N__51104\,
            I => \N__50889\
        );

    \I__12704\ : InMux
    port map (
            O => \N__51103\,
            I => \N__50889\
        );

    \I__12703\ : InMux
    port map (
            O => \N__51102\,
            I => \N__50889\
        );

    \I__12702\ : LocalMux
    port map (
            O => \N__51097\,
            I => \N__50882\
        );

    \I__12701\ : LocalMux
    port map (
            O => \N__51094\,
            I => \N__50882\
        );

    \I__12700\ : LocalMux
    port map (
            O => \N__51089\,
            I => \N__50882\
        );

    \I__12699\ : LocalMux
    port map (
            O => \N__51084\,
            I => \N__50879\
        );

    \I__12698\ : LocalMux
    port map (
            O => \N__51081\,
            I => \N__50874\
        );

    \I__12697\ : LocalMux
    port map (
            O => \N__51074\,
            I => \N__50874\
        );

    \I__12696\ : InMux
    port map (
            O => \N__51073\,
            I => \N__50871\
        );

    \I__12695\ : LocalMux
    port map (
            O => \N__51066\,
            I => \N__50866\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__51061\,
            I => \N__50866\
        );

    \I__12693\ : LocalMux
    port map (
            O => \N__51054\,
            I => \N__50863\
        );

    \I__12692\ : LocalMux
    port map (
            O => \N__51043\,
            I => \N__50854\
        );

    \I__12691\ : LocalMux
    port map (
            O => \N__51040\,
            I => \N__50854\
        );

    \I__12690\ : LocalMux
    port map (
            O => \N__51033\,
            I => \N__50854\
        );

    \I__12689\ : LocalMux
    port map (
            O => \N__51030\,
            I => \N__50854\
        );

    \I__12688\ : LocalMux
    port map (
            O => \N__51027\,
            I => \N__50849\
        );

    \I__12687\ : LocalMux
    port map (
            O => \N__51024\,
            I => \N__50849\
        );

    \I__12686\ : LocalMux
    port map (
            O => \N__51021\,
            I => \N__50844\
        );

    \I__12685\ : LocalMux
    port map (
            O => \N__51018\,
            I => \N__50844\
        );

    \I__12684\ : LocalMux
    port map (
            O => \N__51015\,
            I => \N__50841\
        );

    \I__12683\ : LocalMux
    port map (
            O => \N__51012\,
            I => \N__50834\
        );

    \I__12682\ : LocalMux
    port map (
            O => \N__51005\,
            I => \N__50834\
        );

    \I__12681\ : Span4Mux_h
    port map (
            O => \N__51002\,
            I => \N__50834\
        );

    \I__12680\ : InMux
    port map (
            O => \N__51001\,
            I => \N__50831\
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__50996\,
            I => \N__50828\
        );

    \I__12678\ : CEMux
    port map (
            O => \N__50995\,
            I => \N__50825\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__50992\,
            I => \N__50822\
        );

    \I__12676\ : LocalMux
    port map (
            O => \N__50989\,
            I => \N__50819\
        );

    \I__12675\ : LocalMux
    port map (
            O => \N__50982\,
            I => \N__50812\
        );

    \I__12674\ : Span4Mux_h
    port map (
            O => \N__50977\,
            I => \N__50812\
        );

    \I__12673\ : Span4Mux_h
    port map (
            O => \N__50974\,
            I => \N__50812\
        );

    \I__12672\ : LocalMux
    port map (
            O => \N__50971\,
            I => \N__50807\
        );

    \I__12671\ : Span4Mux_h
    port map (
            O => \N__50966\,
            I => \N__50807\
        );

    \I__12670\ : CEMux
    port map (
            O => \N__50965\,
            I => \N__50804\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__50956\,
            I => \N__50799\
        );

    \I__12668\ : Span4Mux_h
    port map (
            O => \N__50953\,
            I => \N__50799\
        );

    \I__12667\ : InMux
    port map (
            O => \N__50952\,
            I => \N__50790\
        );

    \I__12666\ : InMux
    port map (
            O => \N__50951\,
            I => \N__50790\
        );

    \I__12665\ : InMux
    port map (
            O => \N__50950\,
            I => \N__50790\
        );

    \I__12664\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50790\
        );

    \I__12663\ : InMux
    port map (
            O => \N__50948\,
            I => \N__50775\
        );

    \I__12662\ : InMux
    port map (
            O => \N__50947\,
            I => \N__50775\
        );

    \I__12661\ : InMux
    port map (
            O => \N__50946\,
            I => \N__50775\
        );

    \I__12660\ : InMux
    port map (
            O => \N__50945\,
            I => \N__50775\
        );

    \I__12659\ : InMux
    port map (
            O => \N__50944\,
            I => \N__50775\
        );

    \I__12658\ : InMux
    port map (
            O => \N__50943\,
            I => \N__50775\
        );

    \I__12657\ : InMux
    port map (
            O => \N__50942\,
            I => \N__50775\
        );

    \I__12656\ : InMux
    port map (
            O => \N__50941\,
            I => \N__50764\
        );

    \I__12655\ : InMux
    port map (
            O => \N__50940\,
            I => \N__50764\
        );

    \I__12654\ : InMux
    port map (
            O => \N__50939\,
            I => \N__50764\
        );

    \I__12653\ : InMux
    port map (
            O => \N__50938\,
            I => \N__50764\
        );

    \I__12652\ : InMux
    port map (
            O => \N__50937\,
            I => \N__50764\
        );

    \I__12651\ : InMux
    port map (
            O => \N__50936\,
            I => \N__50753\
        );

    \I__12650\ : InMux
    port map (
            O => \N__50935\,
            I => \N__50753\
        );

    \I__12649\ : InMux
    port map (
            O => \N__50934\,
            I => \N__50753\
        );

    \I__12648\ : InMux
    port map (
            O => \N__50933\,
            I => \N__50753\
        );

    \I__12647\ : InMux
    port map (
            O => \N__50932\,
            I => \N__50753\
        );

    \I__12646\ : InMux
    port map (
            O => \N__50931\,
            I => \N__50744\
        );

    \I__12645\ : InMux
    port map (
            O => \N__50930\,
            I => \N__50744\
        );

    \I__12644\ : InMux
    port map (
            O => \N__50929\,
            I => \N__50744\
        );

    \I__12643\ : InMux
    port map (
            O => \N__50928\,
            I => \N__50744\
        );

    \I__12642\ : InMux
    port map (
            O => \N__50927\,
            I => \N__50737\
        );

    \I__12641\ : InMux
    port map (
            O => \N__50926\,
            I => \N__50737\
        );

    \I__12640\ : InMux
    port map (
            O => \N__50925\,
            I => \N__50737\
        );

    \I__12639\ : InMux
    port map (
            O => \N__50924\,
            I => \N__50728\
        );

    \I__12638\ : InMux
    port map (
            O => \N__50923\,
            I => \N__50728\
        );

    \I__12637\ : InMux
    port map (
            O => \N__50922\,
            I => \N__50728\
        );

    \I__12636\ : InMux
    port map (
            O => \N__50921\,
            I => \N__50728\
        );

    \I__12635\ : LocalMux
    port map (
            O => \N__50908\,
            I => \N__50721\
        );

    \I__12634\ : Span4Mux_v
    port map (
            O => \N__50901\,
            I => \N__50721\
        );

    \I__12633\ : Span4Mux_v
    port map (
            O => \N__50898\,
            I => \N__50721\
        );

    \I__12632\ : LocalMux
    port map (
            O => \N__50889\,
            I => \N__50712\
        );

    \I__12631\ : Span4Mux_h
    port map (
            O => \N__50882\,
            I => \N__50712\
        );

    \I__12630\ : Span4Mux_v
    port map (
            O => \N__50879\,
            I => \N__50712\
        );

    \I__12629\ : Span4Mux_v
    port map (
            O => \N__50874\,
            I => \N__50712\
        );

    \I__12628\ : LocalMux
    port map (
            O => \N__50871\,
            I => \N__50703\
        );

    \I__12627\ : Span4Mux_v
    port map (
            O => \N__50866\,
            I => \N__50703\
        );

    \I__12626\ : Span4Mux_v
    port map (
            O => \N__50863\,
            I => \N__50703\
        );

    \I__12625\ : Span4Mux_v
    port map (
            O => \N__50854\,
            I => \N__50703\
        );

    \I__12624\ : Span4Mux_v
    port map (
            O => \N__50849\,
            I => \N__50694\
        );

    \I__12623\ : Span4Mux_v
    port map (
            O => \N__50844\,
            I => \N__50694\
        );

    \I__12622\ : Span4Mux_v
    port map (
            O => \N__50841\,
            I => \N__50694\
        );

    \I__12621\ : Span4Mux_h
    port map (
            O => \N__50834\,
            I => \N__50694\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__50831\,
            I => \N__50689\
        );

    \I__12619\ : Span4Mux_h
    port map (
            O => \N__50828\,
            I => \N__50689\
        );

    \I__12618\ : LocalMux
    port map (
            O => \N__50825\,
            I => \N__50678\
        );

    \I__12617\ : Span4Mux_h
    port map (
            O => \N__50822\,
            I => \N__50678\
        );

    \I__12616\ : Span4Mux_v
    port map (
            O => \N__50819\,
            I => \N__50678\
        );

    \I__12615\ : Span4Mux_v
    port map (
            O => \N__50812\,
            I => \N__50678\
        );

    \I__12614\ : Span4Mux_h
    port map (
            O => \N__50807\,
            I => \N__50678\
        );

    \I__12613\ : LocalMux
    port map (
            O => \N__50804\,
            I => \N__50673\
        );

    \I__12612\ : Span4Mux_v
    port map (
            O => \N__50799\,
            I => \N__50673\
        );

    \I__12611\ : LocalMux
    port map (
            O => \N__50790\,
            I => n10197
        );

    \I__12610\ : LocalMux
    port map (
            O => \N__50775\,
            I => n10197
        );

    \I__12609\ : LocalMux
    port map (
            O => \N__50764\,
            I => n10197
        );

    \I__12608\ : LocalMux
    port map (
            O => \N__50753\,
            I => n10197
        );

    \I__12607\ : LocalMux
    port map (
            O => \N__50744\,
            I => n10197
        );

    \I__12606\ : LocalMux
    port map (
            O => \N__50737\,
            I => n10197
        );

    \I__12605\ : LocalMux
    port map (
            O => \N__50728\,
            I => n10197
        );

    \I__12604\ : Odrv4
    port map (
            O => \N__50721\,
            I => n10197
        );

    \I__12603\ : Odrv4
    port map (
            O => \N__50712\,
            I => n10197
        );

    \I__12602\ : Odrv4
    port map (
            O => \N__50703\,
            I => n10197
        );

    \I__12601\ : Odrv4
    port map (
            O => \N__50694\,
            I => n10197
        );

    \I__12600\ : Odrv4
    port map (
            O => \N__50689\,
            I => n10197
        );

    \I__12599\ : Odrv4
    port map (
            O => \N__50678\,
            I => n10197
        );

    \I__12598\ : Odrv4
    port map (
            O => \N__50673\,
            I => n10197
        );

    \I__12597\ : CascadeMux
    port map (
            O => \N__50644\,
            I => \N__50641\
        );

    \I__12596\ : InMux
    port map (
            O => \N__50641\,
            I => \N__50638\
        );

    \I__12595\ : LocalMux
    port map (
            O => \N__50638\,
            I => \N__50631\
        );

    \I__12594\ : InMux
    port map (
            O => \N__50637\,
            I => \N__50628\
        );

    \I__12593\ : InMux
    port map (
            O => \N__50636\,
            I => \N__50623\
        );

    \I__12592\ : InMux
    port map (
            O => \N__50635\,
            I => \N__50623\
        );

    \I__12591\ : InMux
    port map (
            O => \N__50634\,
            I => \N__50620\
        );

    \I__12590\ : Span4Mux_h
    port map (
            O => \N__50631\,
            I => \N__50617\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__50628\,
            I => \N__50614\
        );

    \I__12588\ : LocalMux
    port map (
            O => \N__50623\,
            I => \N__50611\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__50620\,
            I => data_out_frame2_16_7
        );

    \I__12586\ : Odrv4
    port map (
            O => \N__50617\,
            I => data_out_frame2_16_7
        );

    \I__12585\ : Odrv12
    port map (
            O => \N__50614\,
            I => data_out_frame2_16_7
        );

    \I__12584\ : Odrv4
    port map (
            O => \N__50611\,
            I => data_out_frame2_16_7
        );

    \I__12583\ : ClkMux
    port map (
            O => \N__50602\,
            I => \N__49924\
        );

    \I__12582\ : ClkMux
    port map (
            O => \N__50601\,
            I => \N__49924\
        );

    \I__12581\ : ClkMux
    port map (
            O => \N__50600\,
            I => \N__49924\
        );

    \I__12580\ : ClkMux
    port map (
            O => \N__50599\,
            I => \N__49924\
        );

    \I__12579\ : ClkMux
    port map (
            O => \N__50598\,
            I => \N__49924\
        );

    \I__12578\ : ClkMux
    port map (
            O => \N__50597\,
            I => \N__49924\
        );

    \I__12577\ : ClkMux
    port map (
            O => \N__50596\,
            I => \N__49924\
        );

    \I__12576\ : ClkMux
    port map (
            O => \N__50595\,
            I => \N__49924\
        );

    \I__12575\ : ClkMux
    port map (
            O => \N__50594\,
            I => \N__49924\
        );

    \I__12574\ : ClkMux
    port map (
            O => \N__50593\,
            I => \N__49924\
        );

    \I__12573\ : ClkMux
    port map (
            O => \N__50592\,
            I => \N__49924\
        );

    \I__12572\ : ClkMux
    port map (
            O => \N__50591\,
            I => \N__49924\
        );

    \I__12571\ : ClkMux
    port map (
            O => \N__50590\,
            I => \N__49924\
        );

    \I__12570\ : ClkMux
    port map (
            O => \N__50589\,
            I => \N__49924\
        );

    \I__12569\ : ClkMux
    port map (
            O => \N__50588\,
            I => \N__49924\
        );

    \I__12568\ : ClkMux
    port map (
            O => \N__50587\,
            I => \N__49924\
        );

    \I__12567\ : ClkMux
    port map (
            O => \N__50586\,
            I => \N__49924\
        );

    \I__12566\ : ClkMux
    port map (
            O => \N__50585\,
            I => \N__49924\
        );

    \I__12565\ : ClkMux
    port map (
            O => \N__50584\,
            I => \N__49924\
        );

    \I__12564\ : ClkMux
    port map (
            O => \N__50583\,
            I => \N__49924\
        );

    \I__12563\ : ClkMux
    port map (
            O => \N__50582\,
            I => \N__49924\
        );

    \I__12562\ : ClkMux
    port map (
            O => \N__50581\,
            I => \N__49924\
        );

    \I__12561\ : ClkMux
    port map (
            O => \N__50580\,
            I => \N__49924\
        );

    \I__12560\ : ClkMux
    port map (
            O => \N__50579\,
            I => \N__49924\
        );

    \I__12559\ : ClkMux
    port map (
            O => \N__50578\,
            I => \N__49924\
        );

    \I__12558\ : ClkMux
    port map (
            O => \N__50577\,
            I => \N__49924\
        );

    \I__12557\ : ClkMux
    port map (
            O => \N__50576\,
            I => \N__49924\
        );

    \I__12556\ : ClkMux
    port map (
            O => \N__50575\,
            I => \N__49924\
        );

    \I__12555\ : ClkMux
    port map (
            O => \N__50574\,
            I => \N__49924\
        );

    \I__12554\ : ClkMux
    port map (
            O => \N__50573\,
            I => \N__49924\
        );

    \I__12553\ : ClkMux
    port map (
            O => \N__50572\,
            I => \N__49924\
        );

    \I__12552\ : ClkMux
    port map (
            O => \N__50571\,
            I => \N__49924\
        );

    \I__12551\ : ClkMux
    port map (
            O => \N__50570\,
            I => \N__49924\
        );

    \I__12550\ : ClkMux
    port map (
            O => \N__50569\,
            I => \N__49924\
        );

    \I__12549\ : ClkMux
    port map (
            O => \N__50568\,
            I => \N__49924\
        );

    \I__12548\ : ClkMux
    port map (
            O => \N__50567\,
            I => \N__49924\
        );

    \I__12547\ : ClkMux
    port map (
            O => \N__50566\,
            I => \N__49924\
        );

    \I__12546\ : ClkMux
    port map (
            O => \N__50565\,
            I => \N__49924\
        );

    \I__12545\ : ClkMux
    port map (
            O => \N__50564\,
            I => \N__49924\
        );

    \I__12544\ : ClkMux
    port map (
            O => \N__50563\,
            I => \N__49924\
        );

    \I__12543\ : ClkMux
    port map (
            O => \N__50562\,
            I => \N__49924\
        );

    \I__12542\ : ClkMux
    port map (
            O => \N__50561\,
            I => \N__49924\
        );

    \I__12541\ : ClkMux
    port map (
            O => \N__50560\,
            I => \N__49924\
        );

    \I__12540\ : ClkMux
    port map (
            O => \N__50559\,
            I => \N__49924\
        );

    \I__12539\ : ClkMux
    port map (
            O => \N__50558\,
            I => \N__49924\
        );

    \I__12538\ : ClkMux
    port map (
            O => \N__50557\,
            I => \N__49924\
        );

    \I__12537\ : ClkMux
    port map (
            O => \N__50556\,
            I => \N__49924\
        );

    \I__12536\ : ClkMux
    port map (
            O => \N__50555\,
            I => \N__49924\
        );

    \I__12535\ : ClkMux
    port map (
            O => \N__50554\,
            I => \N__49924\
        );

    \I__12534\ : ClkMux
    port map (
            O => \N__50553\,
            I => \N__49924\
        );

    \I__12533\ : ClkMux
    port map (
            O => \N__50552\,
            I => \N__49924\
        );

    \I__12532\ : ClkMux
    port map (
            O => \N__50551\,
            I => \N__49924\
        );

    \I__12531\ : ClkMux
    port map (
            O => \N__50550\,
            I => \N__49924\
        );

    \I__12530\ : ClkMux
    port map (
            O => \N__50549\,
            I => \N__49924\
        );

    \I__12529\ : ClkMux
    port map (
            O => \N__50548\,
            I => \N__49924\
        );

    \I__12528\ : ClkMux
    port map (
            O => \N__50547\,
            I => \N__49924\
        );

    \I__12527\ : ClkMux
    port map (
            O => \N__50546\,
            I => \N__49924\
        );

    \I__12526\ : ClkMux
    port map (
            O => \N__50545\,
            I => \N__49924\
        );

    \I__12525\ : ClkMux
    port map (
            O => \N__50544\,
            I => \N__49924\
        );

    \I__12524\ : ClkMux
    port map (
            O => \N__50543\,
            I => \N__49924\
        );

    \I__12523\ : ClkMux
    port map (
            O => \N__50542\,
            I => \N__49924\
        );

    \I__12522\ : ClkMux
    port map (
            O => \N__50541\,
            I => \N__49924\
        );

    \I__12521\ : ClkMux
    port map (
            O => \N__50540\,
            I => \N__49924\
        );

    \I__12520\ : ClkMux
    port map (
            O => \N__50539\,
            I => \N__49924\
        );

    \I__12519\ : ClkMux
    port map (
            O => \N__50538\,
            I => \N__49924\
        );

    \I__12518\ : ClkMux
    port map (
            O => \N__50537\,
            I => \N__49924\
        );

    \I__12517\ : ClkMux
    port map (
            O => \N__50536\,
            I => \N__49924\
        );

    \I__12516\ : ClkMux
    port map (
            O => \N__50535\,
            I => \N__49924\
        );

    \I__12515\ : ClkMux
    port map (
            O => \N__50534\,
            I => \N__49924\
        );

    \I__12514\ : ClkMux
    port map (
            O => \N__50533\,
            I => \N__49924\
        );

    \I__12513\ : ClkMux
    port map (
            O => \N__50532\,
            I => \N__49924\
        );

    \I__12512\ : ClkMux
    port map (
            O => \N__50531\,
            I => \N__49924\
        );

    \I__12511\ : ClkMux
    port map (
            O => \N__50530\,
            I => \N__49924\
        );

    \I__12510\ : ClkMux
    port map (
            O => \N__50529\,
            I => \N__49924\
        );

    \I__12509\ : ClkMux
    port map (
            O => \N__50528\,
            I => \N__49924\
        );

    \I__12508\ : ClkMux
    port map (
            O => \N__50527\,
            I => \N__49924\
        );

    \I__12507\ : ClkMux
    port map (
            O => \N__50526\,
            I => \N__49924\
        );

    \I__12506\ : ClkMux
    port map (
            O => \N__50525\,
            I => \N__49924\
        );

    \I__12505\ : ClkMux
    port map (
            O => \N__50524\,
            I => \N__49924\
        );

    \I__12504\ : ClkMux
    port map (
            O => \N__50523\,
            I => \N__49924\
        );

    \I__12503\ : ClkMux
    port map (
            O => \N__50522\,
            I => \N__49924\
        );

    \I__12502\ : ClkMux
    port map (
            O => \N__50521\,
            I => \N__49924\
        );

    \I__12501\ : ClkMux
    port map (
            O => \N__50520\,
            I => \N__49924\
        );

    \I__12500\ : ClkMux
    port map (
            O => \N__50519\,
            I => \N__49924\
        );

    \I__12499\ : ClkMux
    port map (
            O => \N__50518\,
            I => \N__49924\
        );

    \I__12498\ : ClkMux
    port map (
            O => \N__50517\,
            I => \N__49924\
        );

    \I__12497\ : ClkMux
    port map (
            O => \N__50516\,
            I => \N__49924\
        );

    \I__12496\ : ClkMux
    port map (
            O => \N__50515\,
            I => \N__49924\
        );

    \I__12495\ : ClkMux
    port map (
            O => \N__50514\,
            I => \N__49924\
        );

    \I__12494\ : ClkMux
    port map (
            O => \N__50513\,
            I => \N__49924\
        );

    \I__12493\ : ClkMux
    port map (
            O => \N__50512\,
            I => \N__49924\
        );

    \I__12492\ : ClkMux
    port map (
            O => \N__50511\,
            I => \N__49924\
        );

    \I__12491\ : ClkMux
    port map (
            O => \N__50510\,
            I => \N__49924\
        );

    \I__12490\ : ClkMux
    port map (
            O => \N__50509\,
            I => \N__49924\
        );

    \I__12489\ : ClkMux
    port map (
            O => \N__50508\,
            I => \N__49924\
        );

    \I__12488\ : ClkMux
    port map (
            O => \N__50507\,
            I => \N__49924\
        );

    \I__12487\ : ClkMux
    port map (
            O => \N__50506\,
            I => \N__49924\
        );

    \I__12486\ : ClkMux
    port map (
            O => \N__50505\,
            I => \N__49924\
        );

    \I__12485\ : ClkMux
    port map (
            O => \N__50504\,
            I => \N__49924\
        );

    \I__12484\ : ClkMux
    port map (
            O => \N__50503\,
            I => \N__49924\
        );

    \I__12483\ : ClkMux
    port map (
            O => \N__50502\,
            I => \N__49924\
        );

    \I__12482\ : ClkMux
    port map (
            O => \N__50501\,
            I => \N__49924\
        );

    \I__12481\ : ClkMux
    port map (
            O => \N__50500\,
            I => \N__49924\
        );

    \I__12480\ : ClkMux
    port map (
            O => \N__50499\,
            I => \N__49924\
        );

    \I__12479\ : ClkMux
    port map (
            O => \N__50498\,
            I => \N__49924\
        );

    \I__12478\ : ClkMux
    port map (
            O => \N__50497\,
            I => \N__49924\
        );

    \I__12477\ : ClkMux
    port map (
            O => \N__50496\,
            I => \N__49924\
        );

    \I__12476\ : ClkMux
    port map (
            O => \N__50495\,
            I => \N__49924\
        );

    \I__12475\ : ClkMux
    port map (
            O => \N__50494\,
            I => \N__49924\
        );

    \I__12474\ : ClkMux
    port map (
            O => \N__50493\,
            I => \N__49924\
        );

    \I__12473\ : ClkMux
    port map (
            O => \N__50492\,
            I => \N__49924\
        );

    \I__12472\ : ClkMux
    port map (
            O => \N__50491\,
            I => \N__49924\
        );

    \I__12471\ : ClkMux
    port map (
            O => \N__50490\,
            I => \N__49924\
        );

    \I__12470\ : ClkMux
    port map (
            O => \N__50489\,
            I => \N__49924\
        );

    \I__12469\ : ClkMux
    port map (
            O => \N__50488\,
            I => \N__49924\
        );

    \I__12468\ : ClkMux
    port map (
            O => \N__50487\,
            I => \N__49924\
        );

    \I__12467\ : ClkMux
    port map (
            O => \N__50486\,
            I => \N__49924\
        );

    \I__12466\ : ClkMux
    port map (
            O => \N__50485\,
            I => \N__49924\
        );

    \I__12465\ : ClkMux
    port map (
            O => \N__50484\,
            I => \N__49924\
        );

    \I__12464\ : ClkMux
    port map (
            O => \N__50483\,
            I => \N__49924\
        );

    \I__12463\ : ClkMux
    port map (
            O => \N__50482\,
            I => \N__49924\
        );

    \I__12462\ : ClkMux
    port map (
            O => \N__50481\,
            I => \N__49924\
        );

    \I__12461\ : ClkMux
    port map (
            O => \N__50480\,
            I => \N__49924\
        );

    \I__12460\ : ClkMux
    port map (
            O => \N__50479\,
            I => \N__49924\
        );

    \I__12459\ : ClkMux
    port map (
            O => \N__50478\,
            I => \N__49924\
        );

    \I__12458\ : ClkMux
    port map (
            O => \N__50477\,
            I => \N__49924\
        );

    \I__12457\ : ClkMux
    port map (
            O => \N__50476\,
            I => \N__49924\
        );

    \I__12456\ : ClkMux
    port map (
            O => \N__50475\,
            I => \N__49924\
        );

    \I__12455\ : ClkMux
    port map (
            O => \N__50474\,
            I => \N__49924\
        );

    \I__12454\ : ClkMux
    port map (
            O => \N__50473\,
            I => \N__49924\
        );

    \I__12453\ : ClkMux
    port map (
            O => \N__50472\,
            I => \N__49924\
        );

    \I__12452\ : ClkMux
    port map (
            O => \N__50471\,
            I => \N__49924\
        );

    \I__12451\ : ClkMux
    port map (
            O => \N__50470\,
            I => \N__49924\
        );

    \I__12450\ : ClkMux
    port map (
            O => \N__50469\,
            I => \N__49924\
        );

    \I__12449\ : ClkMux
    port map (
            O => \N__50468\,
            I => \N__49924\
        );

    \I__12448\ : ClkMux
    port map (
            O => \N__50467\,
            I => \N__49924\
        );

    \I__12447\ : ClkMux
    port map (
            O => \N__50466\,
            I => \N__49924\
        );

    \I__12446\ : ClkMux
    port map (
            O => \N__50465\,
            I => \N__49924\
        );

    \I__12445\ : ClkMux
    port map (
            O => \N__50464\,
            I => \N__49924\
        );

    \I__12444\ : ClkMux
    port map (
            O => \N__50463\,
            I => \N__49924\
        );

    \I__12443\ : ClkMux
    port map (
            O => \N__50462\,
            I => \N__49924\
        );

    \I__12442\ : ClkMux
    port map (
            O => \N__50461\,
            I => \N__49924\
        );

    \I__12441\ : ClkMux
    port map (
            O => \N__50460\,
            I => \N__49924\
        );

    \I__12440\ : ClkMux
    port map (
            O => \N__50459\,
            I => \N__49924\
        );

    \I__12439\ : ClkMux
    port map (
            O => \N__50458\,
            I => \N__49924\
        );

    \I__12438\ : ClkMux
    port map (
            O => \N__50457\,
            I => \N__49924\
        );

    \I__12437\ : ClkMux
    port map (
            O => \N__50456\,
            I => \N__49924\
        );

    \I__12436\ : ClkMux
    port map (
            O => \N__50455\,
            I => \N__49924\
        );

    \I__12435\ : ClkMux
    port map (
            O => \N__50454\,
            I => \N__49924\
        );

    \I__12434\ : ClkMux
    port map (
            O => \N__50453\,
            I => \N__49924\
        );

    \I__12433\ : ClkMux
    port map (
            O => \N__50452\,
            I => \N__49924\
        );

    \I__12432\ : ClkMux
    port map (
            O => \N__50451\,
            I => \N__49924\
        );

    \I__12431\ : ClkMux
    port map (
            O => \N__50450\,
            I => \N__49924\
        );

    \I__12430\ : ClkMux
    port map (
            O => \N__50449\,
            I => \N__49924\
        );

    \I__12429\ : ClkMux
    port map (
            O => \N__50448\,
            I => \N__49924\
        );

    \I__12428\ : ClkMux
    port map (
            O => \N__50447\,
            I => \N__49924\
        );

    \I__12427\ : ClkMux
    port map (
            O => \N__50446\,
            I => \N__49924\
        );

    \I__12426\ : ClkMux
    port map (
            O => \N__50445\,
            I => \N__49924\
        );

    \I__12425\ : ClkMux
    port map (
            O => \N__50444\,
            I => \N__49924\
        );

    \I__12424\ : ClkMux
    port map (
            O => \N__50443\,
            I => \N__49924\
        );

    \I__12423\ : ClkMux
    port map (
            O => \N__50442\,
            I => \N__49924\
        );

    \I__12422\ : ClkMux
    port map (
            O => \N__50441\,
            I => \N__49924\
        );

    \I__12421\ : ClkMux
    port map (
            O => \N__50440\,
            I => \N__49924\
        );

    \I__12420\ : ClkMux
    port map (
            O => \N__50439\,
            I => \N__49924\
        );

    \I__12419\ : ClkMux
    port map (
            O => \N__50438\,
            I => \N__49924\
        );

    \I__12418\ : ClkMux
    port map (
            O => \N__50437\,
            I => \N__49924\
        );

    \I__12417\ : ClkMux
    port map (
            O => \N__50436\,
            I => \N__49924\
        );

    \I__12416\ : ClkMux
    port map (
            O => \N__50435\,
            I => \N__49924\
        );

    \I__12415\ : ClkMux
    port map (
            O => \N__50434\,
            I => \N__49924\
        );

    \I__12414\ : ClkMux
    port map (
            O => \N__50433\,
            I => \N__49924\
        );

    \I__12413\ : ClkMux
    port map (
            O => \N__50432\,
            I => \N__49924\
        );

    \I__12412\ : ClkMux
    port map (
            O => \N__50431\,
            I => \N__49924\
        );

    \I__12411\ : ClkMux
    port map (
            O => \N__50430\,
            I => \N__49924\
        );

    \I__12410\ : ClkMux
    port map (
            O => \N__50429\,
            I => \N__49924\
        );

    \I__12409\ : ClkMux
    port map (
            O => \N__50428\,
            I => \N__49924\
        );

    \I__12408\ : ClkMux
    port map (
            O => \N__50427\,
            I => \N__49924\
        );

    \I__12407\ : ClkMux
    port map (
            O => \N__50426\,
            I => \N__49924\
        );

    \I__12406\ : ClkMux
    port map (
            O => \N__50425\,
            I => \N__49924\
        );

    \I__12405\ : ClkMux
    port map (
            O => \N__50424\,
            I => \N__49924\
        );

    \I__12404\ : ClkMux
    port map (
            O => \N__50423\,
            I => \N__49924\
        );

    \I__12403\ : ClkMux
    port map (
            O => \N__50422\,
            I => \N__49924\
        );

    \I__12402\ : ClkMux
    port map (
            O => \N__50421\,
            I => \N__49924\
        );

    \I__12401\ : ClkMux
    port map (
            O => \N__50420\,
            I => \N__49924\
        );

    \I__12400\ : ClkMux
    port map (
            O => \N__50419\,
            I => \N__49924\
        );

    \I__12399\ : ClkMux
    port map (
            O => \N__50418\,
            I => \N__49924\
        );

    \I__12398\ : ClkMux
    port map (
            O => \N__50417\,
            I => \N__49924\
        );

    \I__12397\ : ClkMux
    port map (
            O => \N__50416\,
            I => \N__49924\
        );

    \I__12396\ : ClkMux
    port map (
            O => \N__50415\,
            I => \N__49924\
        );

    \I__12395\ : ClkMux
    port map (
            O => \N__50414\,
            I => \N__49924\
        );

    \I__12394\ : ClkMux
    port map (
            O => \N__50413\,
            I => \N__49924\
        );

    \I__12393\ : ClkMux
    port map (
            O => \N__50412\,
            I => \N__49924\
        );

    \I__12392\ : ClkMux
    port map (
            O => \N__50411\,
            I => \N__49924\
        );

    \I__12391\ : ClkMux
    port map (
            O => \N__50410\,
            I => \N__49924\
        );

    \I__12390\ : ClkMux
    port map (
            O => \N__50409\,
            I => \N__49924\
        );

    \I__12389\ : ClkMux
    port map (
            O => \N__50408\,
            I => \N__49924\
        );

    \I__12388\ : ClkMux
    port map (
            O => \N__50407\,
            I => \N__49924\
        );

    \I__12387\ : ClkMux
    port map (
            O => \N__50406\,
            I => \N__49924\
        );

    \I__12386\ : ClkMux
    port map (
            O => \N__50405\,
            I => \N__49924\
        );

    \I__12385\ : ClkMux
    port map (
            O => \N__50404\,
            I => \N__49924\
        );

    \I__12384\ : ClkMux
    port map (
            O => \N__50403\,
            I => \N__49924\
        );

    \I__12383\ : ClkMux
    port map (
            O => \N__50402\,
            I => \N__49924\
        );

    \I__12382\ : ClkMux
    port map (
            O => \N__50401\,
            I => \N__49924\
        );

    \I__12381\ : ClkMux
    port map (
            O => \N__50400\,
            I => \N__49924\
        );

    \I__12380\ : ClkMux
    port map (
            O => \N__50399\,
            I => \N__49924\
        );

    \I__12379\ : ClkMux
    port map (
            O => \N__50398\,
            I => \N__49924\
        );

    \I__12378\ : ClkMux
    port map (
            O => \N__50397\,
            I => \N__49924\
        );

    \I__12377\ : ClkMux
    port map (
            O => \N__50396\,
            I => \N__49924\
        );

    \I__12376\ : ClkMux
    port map (
            O => \N__50395\,
            I => \N__49924\
        );

    \I__12375\ : ClkMux
    port map (
            O => \N__50394\,
            I => \N__49924\
        );

    \I__12374\ : ClkMux
    port map (
            O => \N__50393\,
            I => \N__49924\
        );

    \I__12373\ : ClkMux
    port map (
            O => \N__50392\,
            I => \N__49924\
        );

    \I__12372\ : ClkMux
    port map (
            O => \N__50391\,
            I => \N__49924\
        );

    \I__12371\ : ClkMux
    port map (
            O => \N__50390\,
            I => \N__49924\
        );

    \I__12370\ : ClkMux
    port map (
            O => \N__50389\,
            I => \N__49924\
        );

    \I__12369\ : ClkMux
    port map (
            O => \N__50388\,
            I => \N__49924\
        );

    \I__12368\ : ClkMux
    port map (
            O => \N__50387\,
            I => \N__49924\
        );

    \I__12367\ : ClkMux
    port map (
            O => \N__50386\,
            I => \N__49924\
        );

    \I__12366\ : ClkMux
    port map (
            O => \N__50385\,
            I => \N__49924\
        );

    \I__12365\ : ClkMux
    port map (
            O => \N__50384\,
            I => \N__49924\
        );

    \I__12364\ : ClkMux
    port map (
            O => \N__50383\,
            I => \N__49924\
        );

    \I__12363\ : ClkMux
    port map (
            O => \N__50382\,
            I => \N__49924\
        );

    \I__12362\ : ClkMux
    port map (
            O => \N__50381\,
            I => \N__49924\
        );

    \I__12361\ : ClkMux
    port map (
            O => \N__50380\,
            I => \N__49924\
        );

    \I__12360\ : ClkMux
    port map (
            O => \N__50379\,
            I => \N__49924\
        );

    \I__12359\ : ClkMux
    port map (
            O => \N__50378\,
            I => \N__49924\
        );

    \I__12358\ : ClkMux
    port map (
            O => \N__50377\,
            I => \N__49924\
        );

    \I__12357\ : GlobalMux
    port map (
            O => \N__49924\,
            I => \N__49921\
        );

    \I__12356\ : gio2CtrlBuf
    port map (
            O => \N__49921\,
            I => \CLK_c\
        );

    \I__12355\ : InMux
    port map (
            O => \N__49918\,
            I => \N__49913\
        );

    \I__12354\ : InMux
    port map (
            O => \N__49917\,
            I => \N__49910\
        );

    \I__12353\ : InMux
    port map (
            O => \N__49916\,
            I => \N__49907\
        );

    \I__12352\ : LocalMux
    port map (
            O => \N__49913\,
            I => \N__49901\
        );

    \I__12351\ : LocalMux
    port map (
            O => \N__49910\,
            I => \N__49901\
        );

    \I__12350\ : LocalMux
    port map (
            O => \N__49907\,
            I => \N__49898\
        );

    \I__12349\ : InMux
    port map (
            O => \N__49906\,
            I => \N__49894\
        );

    \I__12348\ : Span4Mux_v
    port map (
            O => \N__49901\,
            I => \N__49891\
        );

    \I__12347\ : Span4Mux_v
    port map (
            O => \N__49898\,
            I => \N__49888\
        );

    \I__12346\ : InMux
    port map (
            O => \N__49897\,
            I => \N__49885\
        );

    \I__12345\ : LocalMux
    port map (
            O => \N__49894\,
            I => \N__49882\
        );

    \I__12344\ : Span4Mux_h
    port map (
            O => \N__49891\,
            I => \N__49879\
        );

    \I__12343\ : Span4Mux_h
    port map (
            O => \N__49888\,
            I => \N__49873\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__49885\,
            I => \N__49873\
        );

    \I__12341\ : Span4Mux_h
    port map (
            O => \N__49882\,
            I => \N__49868\
        );

    \I__12340\ : Span4Mux_h
    port map (
            O => \N__49879\,
            I => \N__49868\
        );

    \I__12339\ : InMux
    port map (
            O => \N__49878\,
            I => \N__49865\
        );

    \I__12338\ : Span4Mux_v
    port map (
            O => \N__49873\,
            I => \N__49862\
        );

    \I__12337\ : Odrv4
    port map (
            O => \N__49868\,
            I => rand_data_6
        );

    \I__12336\ : LocalMux
    port map (
            O => \N__49865\,
            I => rand_data_6
        );

    \I__12335\ : Odrv4
    port map (
            O => \N__49862\,
            I => rand_data_6
        );

    \I__12334\ : CascadeMux
    port map (
            O => \N__49855\,
            I => \N__49851\
        );

    \I__12333\ : InMux
    port map (
            O => \N__49854\,
            I => \N__49848\
        );

    \I__12332\ : InMux
    port map (
            O => \N__49851\,
            I => \N__49844\
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__49848\,
            I => \N__49840\
        );

    \I__12330\ : InMux
    port map (
            O => \N__49847\,
            I => \N__49837\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__49844\,
            I => \N__49834\
        );

    \I__12328\ : InMux
    port map (
            O => \N__49843\,
            I => \N__49831\
        );

    \I__12327\ : Span4Mux_v
    port map (
            O => \N__49840\,
            I => \N__49828\
        );

    \I__12326\ : LocalMux
    port map (
            O => \N__49837\,
            I => \N__49825\
        );

    \I__12325\ : Span4Mux_h
    port map (
            O => \N__49834\,
            I => \N__49822\
        );

    \I__12324\ : LocalMux
    port map (
            O => \N__49831\,
            I => data_out_frame2_16_6
        );

    \I__12323\ : Odrv4
    port map (
            O => \N__49828\,
            I => data_out_frame2_16_6
        );

    \I__12322\ : Odrv12
    port map (
            O => \N__49825\,
            I => data_out_frame2_16_6
        );

    \I__12321\ : Odrv4
    port map (
            O => \N__49822\,
            I => data_out_frame2_16_6
        );

    \I__12320\ : InMux
    port map (
            O => \N__49813\,
            I => \N__49810\
        );

    \I__12319\ : LocalMux
    port map (
            O => \N__49810\,
            I => \N__49806\
        );

    \I__12318\ : InMux
    port map (
            O => \N__49809\,
            I => \N__49803\
        );

    \I__12317\ : Span4Mux_h
    port map (
            O => \N__49806\,
            I => \N__49796\
        );

    \I__12316\ : LocalMux
    port map (
            O => \N__49803\,
            I => \N__49796\
        );

    \I__12315\ : InMux
    port map (
            O => \N__49802\,
            I => \N__49793\
        );

    \I__12314\ : InMux
    port map (
            O => \N__49801\,
            I => \N__49790\
        );

    \I__12313\ : Span4Mux_v
    port map (
            O => \N__49796\,
            I => \N__49785\
        );

    \I__12312\ : LocalMux
    port map (
            O => \N__49793\,
            I => \N__49785\
        );

    \I__12311\ : LocalMux
    port map (
            O => \N__49790\,
            I => \N__49781\
        );

    \I__12310\ : Span4Mux_h
    port map (
            O => \N__49785\,
            I => \N__49777\
        );

    \I__12309\ : InMux
    port map (
            O => \N__49784\,
            I => \N__49774\
        );

    \I__12308\ : Span12Mux_v
    port map (
            O => \N__49781\,
            I => \N__49771\
        );

    \I__12307\ : InMux
    port map (
            O => \N__49780\,
            I => \N__49768\
        );

    \I__12306\ : Sp12to4
    port map (
            O => \N__49777\,
            I => \N__49763\
        );

    \I__12305\ : LocalMux
    port map (
            O => \N__49774\,
            I => \N__49763\
        );

    \I__12304\ : Odrv12
    port map (
            O => \N__49771\,
            I => rand_data_3
        );

    \I__12303\ : LocalMux
    port map (
            O => \N__49768\,
            I => rand_data_3
        );

    \I__12302\ : Odrv12
    port map (
            O => \N__49763\,
            I => rand_data_3
        );

    \I__12301\ : InMux
    port map (
            O => \N__49756\,
            I => \N__49752\
        );

    \I__12300\ : InMux
    port map (
            O => \N__49755\,
            I => \N__49749\
        );

    \I__12299\ : LocalMux
    port map (
            O => \N__49752\,
            I => data_out_frame2_18_3
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__49749\,
            I => data_out_frame2_18_3
        );

    \I__12297\ : CascadeMux
    port map (
            O => \N__49744\,
            I => \N__49739\
        );

    \I__12296\ : InMux
    port map (
            O => \N__49743\,
            I => \N__49736\
        );

    \I__12295\ : InMux
    port map (
            O => \N__49742\,
            I => \N__49732\
        );

    \I__12294\ : InMux
    port map (
            O => \N__49739\,
            I => \N__49729\
        );

    \I__12293\ : LocalMux
    port map (
            O => \N__49736\,
            I => \N__49726\
        );

    \I__12292\ : InMux
    port map (
            O => \N__49735\,
            I => \N__49723\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__49732\,
            I => \N__49720\
        );

    \I__12290\ : LocalMux
    port map (
            O => \N__49729\,
            I => \N__49717\
        );

    \I__12289\ : Span4Mux_v
    port map (
            O => \N__49726\,
            I => \N__49714\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__49723\,
            I => \N__49707\
        );

    \I__12287\ : Span4Mux_v
    port map (
            O => \N__49720\,
            I => \N__49707\
        );

    \I__12286\ : Span4Mux_h
    port map (
            O => \N__49717\,
            I => \N__49707\
        );

    \I__12285\ : Odrv4
    port map (
            O => \N__49714\,
            I => data_out_frame2_15_5
        );

    \I__12284\ : Odrv4
    port map (
            O => \N__49707\,
            I => data_out_frame2_15_5
        );

    \I__12283\ : InMux
    port map (
            O => \N__49702\,
            I => \N__49699\
        );

    \I__12282\ : LocalMux
    port map (
            O => \N__49699\,
            I => \N__49695\
        );

    \I__12281\ : InMux
    port map (
            O => \N__49698\,
            I => \N__49692\
        );

    \I__12280\ : Span4Mux_h
    port map (
            O => \N__49695\,
            I => \N__49687\
        );

    \I__12279\ : LocalMux
    port map (
            O => \N__49692\,
            I => \N__49687\
        );

    \I__12278\ : Span4Mux_v
    port map (
            O => \N__49687\,
            I => \N__49681\
        );

    \I__12277\ : InMux
    port map (
            O => \N__49686\,
            I => \N__49676\
        );

    \I__12276\ : InMux
    port map (
            O => \N__49685\,
            I => \N__49676\
        );

    \I__12275\ : InMux
    port map (
            O => \N__49684\,
            I => \N__49673\
        );

    \I__12274\ : Span4Mux_h
    port map (
            O => \N__49681\,
            I => \N__49670\
        );

    \I__12273\ : LocalMux
    port map (
            O => \N__49676\,
            I => data_out_frame2_11_0
        );

    \I__12272\ : LocalMux
    port map (
            O => \N__49673\,
            I => data_out_frame2_11_0
        );

    \I__12271\ : Odrv4
    port map (
            O => \N__49670\,
            I => data_out_frame2_11_0
        );

    \I__12270\ : InMux
    port map (
            O => \N__49663\,
            I => \N__49660\
        );

    \I__12269\ : LocalMux
    port map (
            O => \N__49660\,
            I => \N__49655\
        );

    \I__12268\ : InMux
    port map (
            O => \N__49659\,
            I => \N__49652\
        );

    \I__12267\ : CascadeMux
    port map (
            O => \N__49658\,
            I => \N__49648\
        );

    \I__12266\ : Span12Mux_s9_v
    port map (
            O => \N__49655\,
            I => \N__49643\
        );

    \I__12265\ : LocalMux
    port map (
            O => \N__49652\,
            I => \N__49643\
        );

    \I__12264\ : InMux
    port map (
            O => \N__49651\,
            I => \N__49638\
        );

    \I__12263\ : InMux
    port map (
            O => \N__49648\,
            I => \N__49638\
        );

    \I__12262\ : Odrv12
    port map (
            O => \N__49643\,
            I => data_out_frame2_13_6
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__49638\,
            I => data_out_frame2_13_6
        );

    \I__12260\ : InMux
    port map (
            O => \N__49633\,
            I => \N__49630\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__49630\,
            I => \N__49626\
        );

    \I__12258\ : InMux
    port map (
            O => \N__49629\,
            I => \N__49623\
        );

    \I__12257\ : Span4Mux_h
    port map (
            O => \N__49626\,
            I => \N__49620\
        );

    \I__12256\ : LocalMux
    port map (
            O => \N__49623\,
            I => \N__49617\
        );

    \I__12255\ : Span4Mux_h
    port map (
            O => \N__49620\,
            I => \N__49614\
        );

    \I__12254\ : Span4Mux_h
    port map (
            O => \N__49617\,
            I => \N__49611\
        );

    \I__12253\ : Span4Mux_h
    port map (
            O => \N__49614\,
            I => \N__49608\
        );

    \I__12252\ : Odrv4
    port map (
            O => \N__49611\,
            I => \c0.n16923\
        );

    \I__12251\ : Odrv4
    port map (
            O => \N__49608\,
            I => \c0.n16923\
        );

    \I__12250\ : CascadeMux
    port map (
            O => \N__49603\,
            I => \N__49600\
        );

    \I__12249\ : InMux
    port map (
            O => \N__49600\,
            I => \N__49597\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__49597\,
            I => \N__49592\
        );

    \I__12247\ : InMux
    port map (
            O => \N__49596\,
            I => \N__49589\
        );

    \I__12246\ : InMux
    port map (
            O => \N__49595\,
            I => \N__49586\
        );

    \I__12245\ : Span12Mux_h
    port map (
            O => \N__49592\,
            I => \N__49583\
        );

    \I__12244\ : LocalMux
    port map (
            O => \N__49589\,
            I => data_out_frame2_13_1
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__49586\,
            I => data_out_frame2_13_1
        );

    \I__12242\ : Odrv12
    port map (
            O => \N__49583\,
            I => data_out_frame2_13_1
        );

    \I__12241\ : InMux
    port map (
            O => \N__49576\,
            I => \N__49573\
        );

    \I__12240\ : LocalMux
    port map (
            O => \N__49573\,
            I => \N__49570\
        );

    \I__12239\ : Span4Mux_h
    port map (
            O => \N__49570\,
            I => \N__49567\
        );

    \I__12238\ : Odrv4
    port map (
            O => \N__49567\,
            I => \c0.n9910\
        );

    \I__12237\ : InMux
    port map (
            O => \N__49564\,
            I => \N__49561\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__49561\,
            I => \N__49558\
        );

    \I__12235\ : Span4Mux_v
    port map (
            O => \N__49558\,
            I => \N__49554\
        );

    \I__12234\ : InMux
    port map (
            O => \N__49557\,
            I => \N__49551\
        );

    \I__12233\ : Span4Mux_v
    port map (
            O => \N__49554\,
            I => \N__49548\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__49551\,
            I => \N__49545\
        );

    \I__12231\ : Odrv4
    port map (
            O => \N__49548\,
            I => \c0.n9826\
        );

    \I__12230\ : Odrv4
    port map (
            O => \N__49545\,
            I => \c0.n9826\
        );

    \I__12229\ : InMux
    port map (
            O => \N__49540\,
            I => \N__49537\
        );

    \I__12228\ : LocalMux
    port map (
            O => \N__49537\,
            I => \N__49532\
        );

    \I__12227\ : InMux
    port map (
            O => \N__49536\,
            I => \N__49529\
        );

    \I__12226\ : InMux
    port map (
            O => \N__49535\,
            I => \N__49526\
        );

    \I__12225\ : Span4Mux_h
    port map (
            O => \N__49532\,
            I => \N__49518\
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__49529\,
            I => \N__49518\
        );

    \I__12223\ : LocalMux
    port map (
            O => \N__49526\,
            I => \N__49518\
        );

    \I__12222\ : InMux
    port map (
            O => \N__49525\,
            I => \N__49515\
        );

    \I__12221\ : Span4Mux_h
    port map (
            O => \N__49518\,
            I => \N__49512\
        );

    \I__12220\ : LocalMux
    port map (
            O => \N__49515\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__12219\ : Odrv4
    port map (
            O => \N__49512\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__12218\ : CascadeMux
    port map (
            O => \N__49507\,
            I => \c0.n9910_cascade_\
        );

    \I__12217\ : InMux
    port map (
            O => \N__49504\,
            I => \N__49500\
        );

    \I__12216\ : InMux
    port map (
            O => \N__49503\,
            I => \N__49497\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__49500\,
            I => \N__49494\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__49497\,
            I => \N__49491\
        );

    \I__12213\ : Span4Mux_v
    port map (
            O => \N__49494\,
            I => \N__49488\
        );

    \I__12212\ : Span4Mux_v
    port map (
            O => \N__49491\,
            I => \N__49485\
        );

    \I__12211\ : Span4Mux_v
    port map (
            O => \N__49488\,
            I => \N__49480\
        );

    \I__12210\ : Span4Mux_v
    port map (
            O => \N__49485\,
            I => \N__49480\
        );

    \I__12209\ : Odrv4
    port map (
            O => \N__49480\,
            I => \c0.n9843\
        );

    \I__12208\ : InMux
    port map (
            O => \N__49477\,
            I => \N__49473\
        );

    \I__12207\ : CascadeMux
    port map (
            O => \N__49476\,
            I => \N__49470\
        );

    \I__12206\ : LocalMux
    port map (
            O => \N__49473\,
            I => \N__49466\
        );

    \I__12205\ : InMux
    port map (
            O => \N__49470\,
            I => \N__49463\
        );

    \I__12204\ : CascadeMux
    port map (
            O => \N__49469\,
            I => \N__49460\
        );

    \I__12203\ : Span4Mux_v
    port map (
            O => \N__49466\,
            I => \N__49456\
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__49463\,
            I => \N__49453\
        );

    \I__12201\ : InMux
    port map (
            O => \N__49460\,
            I => \N__49450\
        );

    \I__12200\ : InMux
    port map (
            O => \N__49459\,
            I => \N__49447\
        );

    \I__12199\ : Span4Mux_h
    port map (
            O => \N__49456\,
            I => \N__49442\
        );

    \I__12198\ : Span4Mux_v
    port map (
            O => \N__49453\,
            I => \N__49442\
        );

    \I__12197\ : LocalMux
    port map (
            O => \N__49450\,
            I => \N__49439\
        );

    \I__12196\ : LocalMux
    port map (
            O => \N__49447\,
            I => data_out_frame2_14_1
        );

    \I__12195\ : Odrv4
    port map (
            O => \N__49442\,
            I => data_out_frame2_14_1
        );

    \I__12194\ : Odrv12
    port map (
            O => \N__49439\,
            I => data_out_frame2_14_1
        );

    \I__12193\ : InMux
    port map (
            O => \N__49432\,
            I => \N__49428\
        );

    \I__12192\ : InMux
    port map (
            O => \N__49431\,
            I => \N__49424\
        );

    \I__12191\ : LocalMux
    port map (
            O => \N__49428\,
            I => \N__49420\
        );

    \I__12190\ : InMux
    port map (
            O => \N__49427\,
            I => \N__49417\
        );

    \I__12189\ : LocalMux
    port map (
            O => \N__49424\,
            I => \N__49412\
        );

    \I__12188\ : InMux
    port map (
            O => \N__49423\,
            I => \N__49409\
        );

    \I__12187\ : Span4Mux_h
    port map (
            O => \N__49420\,
            I => \N__49406\
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__49417\,
            I => \N__49403\
        );

    \I__12185\ : InMux
    port map (
            O => \N__49416\,
            I => \N__49398\
        );

    \I__12184\ : InMux
    port map (
            O => \N__49415\,
            I => \N__49398\
        );

    \I__12183\ : Span4Mux_h
    port map (
            O => \N__49412\,
            I => \N__49393\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__49409\,
            I => \N__49393\
        );

    \I__12181\ : Odrv4
    port map (
            O => \N__49406\,
            I => data_out_frame2_8_0
        );

    \I__12180\ : Odrv12
    port map (
            O => \N__49403\,
            I => data_out_frame2_8_0
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__49398\,
            I => data_out_frame2_8_0
        );

    \I__12178\ : Odrv4
    port map (
            O => \N__49393\,
            I => data_out_frame2_8_0
        );

    \I__12177\ : CascadeMux
    port map (
            O => \N__49384\,
            I => \N__49381\
        );

    \I__12176\ : InMux
    port map (
            O => \N__49381\,
            I => \N__49375\
        );

    \I__12175\ : InMux
    port map (
            O => \N__49380\,
            I => \N__49372\
        );

    \I__12174\ : InMux
    port map (
            O => \N__49379\,
            I => \N__49369\
        );

    \I__12173\ : CascadeMux
    port map (
            O => \N__49378\,
            I => \N__49366\
        );

    \I__12172\ : LocalMux
    port map (
            O => \N__49375\,
            I => \N__49362\
        );

    \I__12171\ : LocalMux
    port map (
            O => \N__49372\,
            I => \N__49357\
        );

    \I__12170\ : LocalMux
    port map (
            O => \N__49369\,
            I => \N__49357\
        );

    \I__12169\ : InMux
    port map (
            O => \N__49366\,
            I => \N__49352\
        );

    \I__12168\ : InMux
    port map (
            O => \N__49365\,
            I => \N__49352\
        );

    \I__12167\ : Odrv4
    port map (
            O => \N__49362\,
            I => data_out_frame2_15_0
        );

    \I__12166\ : Odrv12
    port map (
            O => \N__49357\,
            I => data_out_frame2_15_0
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__49352\,
            I => data_out_frame2_15_0
        );

    \I__12164\ : InMux
    port map (
            O => \N__49345\,
            I => \N__49340\
        );

    \I__12163\ : InMux
    port map (
            O => \N__49344\,
            I => \N__49337\
        );

    \I__12162\ : InMux
    port map (
            O => \N__49343\,
            I => \N__49334\
        );

    \I__12161\ : LocalMux
    port map (
            O => \N__49340\,
            I => \N__49331\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__49337\,
            I => \N__49328\
        );

    \I__12159\ : LocalMux
    port map (
            O => \N__49334\,
            I => \N__49325\
        );

    \I__12158\ : Span4Mux_h
    port map (
            O => \N__49331\,
            I => \N__49320\
        );

    \I__12157\ : Span4Mux_v
    port map (
            O => \N__49328\,
            I => \N__49317\
        );

    \I__12156\ : Span4Mux_h
    port map (
            O => \N__49325\,
            I => \N__49314\
        );

    \I__12155\ : InMux
    port map (
            O => \N__49324\,
            I => \N__49309\
        );

    \I__12154\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49309\
        );

    \I__12153\ : Odrv4
    port map (
            O => \N__49320\,
            I => data_out_frame2_8_4
        );

    \I__12152\ : Odrv4
    port map (
            O => \N__49317\,
            I => data_out_frame2_8_4
        );

    \I__12151\ : Odrv4
    port map (
            O => \N__49314\,
            I => data_out_frame2_8_4
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__49309\,
            I => data_out_frame2_8_4
        );

    \I__12149\ : InMux
    port map (
            O => \N__49300\,
            I => \N__49297\
        );

    \I__12148\ : LocalMux
    port map (
            O => \N__49297\,
            I => \c0.n16_adj_2327\
        );

    \I__12147\ : InMux
    port map (
            O => \N__49294\,
            I => \N__49291\
        );

    \I__12146\ : LocalMux
    port map (
            O => \N__49291\,
            I => \N__49287\
        );

    \I__12145\ : CascadeMux
    port map (
            O => \N__49290\,
            I => \N__49284\
        );

    \I__12144\ : Span4Mux_h
    port map (
            O => \N__49287\,
            I => \N__49280\
        );

    \I__12143\ : InMux
    port map (
            O => \N__49284\,
            I => \N__49277\
        );

    \I__12142\ : CascadeMux
    port map (
            O => \N__49283\,
            I => \N__49274\
        );

    \I__12141\ : Span4Mux_h
    port map (
            O => \N__49280\,
            I => \N__49266\
        );

    \I__12140\ : LocalMux
    port map (
            O => \N__49277\,
            I => \N__49266\
        );

    \I__12139\ : InMux
    port map (
            O => \N__49274\,
            I => \N__49263\
        );

    \I__12138\ : InMux
    port map (
            O => \N__49273\,
            I => \N__49260\
        );

    \I__12137\ : InMux
    port map (
            O => \N__49272\,
            I => \N__49257\
        );

    \I__12136\ : InMux
    port map (
            O => \N__49271\,
            I => \N__49254\
        );

    \I__12135\ : Span4Mux_v
    port map (
            O => \N__49266\,
            I => \N__49251\
        );

    \I__12134\ : LocalMux
    port map (
            O => \N__49263\,
            I => \N__49246\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__49260\,
            I => \N__49246\
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__49257\,
            I => data_out_frame2_12_2
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__49254\,
            I => data_out_frame2_12_2
        );

    \I__12130\ : Odrv4
    port map (
            O => \N__49251\,
            I => data_out_frame2_12_2
        );

    \I__12129\ : Odrv12
    port map (
            O => \N__49246\,
            I => data_out_frame2_12_2
        );

    \I__12128\ : CascadeMux
    port map (
            O => \N__49237\,
            I => \c0.n17_adj_2328_cascade_\
        );

    \I__12127\ : InMux
    port map (
            O => \N__49234\,
            I => \N__49231\
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__49231\,
            I => \N__49228\
        );

    \I__12125\ : Span4Mux_h
    port map (
            O => \N__49228\,
            I => \N__49224\
        );

    \I__12124\ : InMux
    port map (
            O => \N__49227\,
            I => \N__49221\
        );

    \I__12123\ : Odrv4
    port map (
            O => \N__49224\,
            I => \c0.n17010\
        );

    \I__12122\ : LocalMux
    port map (
            O => \N__49221\,
            I => \c0.n17010\
        );

    \I__12121\ : CascadeMux
    port map (
            O => \N__49216\,
            I => \N__49213\
        );

    \I__12120\ : InMux
    port map (
            O => \N__49213\,
            I => \N__49210\
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__49210\,
            I => \N__49207\
        );

    \I__12118\ : Span4Mux_h
    port map (
            O => \N__49207\,
            I => \N__49204\
        );

    \I__12117\ : Span4Mux_h
    port map (
            O => \N__49204\,
            I => \N__49201\
        );

    \I__12116\ : Odrv4
    port map (
            O => \N__49201\,
            I => \c0.data_out_frame2_19_1\
        );

    \I__12115\ : InMux
    port map (
            O => \N__49198\,
            I => \N__49195\
        );

    \I__12114\ : LocalMux
    port map (
            O => \N__49195\,
            I => \N__49191\
        );

    \I__12113\ : InMux
    port map (
            O => \N__49194\,
            I => \N__49188\
        );

    \I__12112\ : Span4Mux_h
    port map (
            O => \N__49191\,
            I => \N__49184\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__49188\,
            I => \N__49179\
        );

    \I__12110\ : InMux
    port map (
            O => \N__49187\,
            I => \N__49176\
        );

    \I__12109\ : Span4Mux_v
    port map (
            O => \N__49184\,
            I => \N__49173\
        );

    \I__12108\ : InMux
    port map (
            O => \N__49183\,
            I => \N__49168\
        );

    \I__12107\ : InMux
    port map (
            O => \N__49182\,
            I => \N__49168\
        );

    \I__12106\ : Span4Mux_h
    port map (
            O => \N__49179\,
            I => \N__49165\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__49176\,
            I => data_out_frame2_15_7
        );

    \I__12104\ : Odrv4
    port map (
            O => \N__49173\,
            I => data_out_frame2_15_7
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__49168\,
            I => data_out_frame2_15_7
        );

    \I__12102\ : Odrv4
    port map (
            O => \N__49165\,
            I => data_out_frame2_15_7
        );

    \I__12101\ : CascadeMux
    port map (
            O => \N__49156\,
            I => \N__49153\
        );

    \I__12100\ : InMux
    port map (
            O => \N__49153\,
            I => \N__49150\
        );

    \I__12099\ : LocalMux
    port map (
            O => \N__49150\,
            I => \N__49147\
        );

    \I__12098\ : Odrv4
    port map (
            O => \N__49147\,
            I => \c0.n16940\
        );

    \I__12097\ : InMux
    port map (
            O => \N__49144\,
            I => \N__49141\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__49141\,
            I => \c0.n26_adj_2314\
        );

    \I__12095\ : InMux
    port map (
            O => \N__49138\,
            I => \N__49135\
        );

    \I__12094\ : LocalMux
    port map (
            O => \N__49135\,
            I => \N__49132\
        );

    \I__12093\ : Span4Mux_h
    port map (
            O => \N__49132\,
            I => \N__49129\
        );

    \I__12092\ : Odrv4
    port map (
            O => \N__49129\,
            I => \c0.n25_adj_2316\
        );

    \I__12091\ : CascadeMux
    port map (
            O => \N__49126\,
            I => \c0.n23_adj_2318_cascade_\
        );

    \I__12090\ : InMux
    port map (
            O => \N__49123\,
            I => \N__49120\
        );

    \I__12089\ : LocalMux
    port map (
            O => \N__49120\,
            I => \N__49117\
        );

    \I__12088\ : Span4Mux_v
    port map (
            O => \N__49117\,
            I => \N__49114\
        );

    \I__12087\ : Odrv4
    port map (
            O => \N__49114\,
            I => \c0.n24_adj_2315\
        );

    \I__12086\ : CascadeMux
    port map (
            O => \N__49111\,
            I => \N__49107\
        );

    \I__12085\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49103\
        );

    \I__12084\ : InMux
    port map (
            O => \N__49107\,
            I => \N__49099\
        );

    \I__12083\ : InMux
    port map (
            O => \N__49106\,
            I => \N__49096\
        );

    \I__12082\ : LocalMux
    port map (
            O => \N__49103\,
            I => \N__49092\
        );

    \I__12081\ : InMux
    port map (
            O => \N__49102\,
            I => \N__49089\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__49099\,
            I => \N__49086\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__49096\,
            I => \N__49083\
        );

    \I__12078\ : InMux
    port map (
            O => \N__49095\,
            I => \N__49080\
        );

    \I__12077\ : Span4Mux_h
    port map (
            O => \N__49092\,
            I => \N__49077\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__49089\,
            I => \N__49074\
        );

    \I__12075\ : Span4Mux_v
    port map (
            O => \N__49086\,
            I => \N__49068\
        );

    \I__12074\ : Span4Mux_v
    port map (
            O => \N__49083\,
            I => \N__49068\
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__49080\,
            I => \N__49065\
        );

    \I__12072\ : Span4Mux_h
    port map (
            O => \N__49077\,
            I => \N__49062\
        );

    \I__12071\ : Span4Mux_h
    port map (
            O => \N__49074\,
            I => \N__49059\
        );

    \I__12070\ : InMux
    port map (
            O => \N__49073\,
            I => \N__49056\
        );

    \I__12069\ : Span4Mux_h
    port map (
            O => \N__49068\,
            I => \N__49051\
        );

    \I__12068\ : Span4Mux_s3_v
    port map (
            O => \N__49065\,
            I => \N__49051\
        );

    \I__12067\ : Odrv4
    port map (
            O => \N__49062\,
            I => rand_data_14
        );

    \I__12066\ : Odrv4
    port map (
            O => \N__49059\,
            I => rand_data_14
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__49056\,
            I => rand_data_14
        );

    \I__12064\ : Odrv4
    port map (
            O => \N__49051\,
            I => rand_data_14
        );

    \I__12063\ : CascadeMux
    port map (
            O => \N__49042\,
            I => \N__49039\
        );

    \I__12062\ : InMux
    port map (
            O => \N__49039\,
            I => \N__49035\
        );

    \I__12061\ : InMux
    port map (
            O => \N__49038\,
            I => \N__49032\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__49035\,
            I => \N__49029\
        );

    \I__12059\ : LocalMux
    port map (
            O => \N__49032\,
            I => data_out_frame2_17_6
        );

    \I__12058\ : Odrv12
    port map (
            O => \N__49029\,
            I => data_out_frame2_17_6
        );

    \I__12057\ : InMux
    port map (
            O => \N__49024\,
            I => \N__49021\
        );

    \I__12056\ : LocalMux
    port map (
            O => \N__49021\,
            I => \c0.data_out_frame2_19_3\
        );

    \I__12055\ : CascadeMux
    port map (
            O => \N__49018\,
            I => \c0.n17945_cascade_\
        );

    \I__12054\ : InMux
    port map (
            O => \N__49015\,
            I => \N__49012\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__49012\,
            I => \N__49008\
        );

    \I__12052\ : InMux
    port map (
            O => \N__49011\,
            I => \N__49004\
        );

    \I__12051\ : Span4Mux_v
    port map (
            O => \N__49008\,
            I => \N__49000\
        );

    \I__12050\ : InMux
    port map (
            O => \N__49007\,
            I => \N__48997\
        );

    \I__12049\ : LocalMux
    port map (
            O => \N__49004\,
            I => \N__48994\
        );

    \I__12048\ : InMux
    port map (
            O => \N__49003\,
            I => \N__48990\
        );

    \I__12047\ : Span4Mux_h
    port map (
            O => \N__49000\,
            I => \N__48986\
        );

    \I__12046\ : LocalMux
    port map (
            O => \N__48997\,
            I => \N__48981\
        );

    \I__12045\ : Span4Mux_h
    port map (
            O => \N__48994\,
            I => \N__48981\
        );

    \I__12044\ : InMux
    port map (
            O => \N__48993\,
            I => \N__48978\
        );

    \I__12043\ : LocalMux
    port map (
            O => \N__48990\,
            I => \N__48975\
        );

    \I__12042\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48972\
        );

    \I__12041\ : Span4Mux_h
    port map (
            O => \N__48986\,
            I => \N__48969\
        );

    \I__12040\ : Span4Mux_h
    port map (
            O => \N__48981\,
            I => \N__48966\
        );

    \I__12039\ : LocalMux
    port map (
            O => \N__48978\,
            I => data_out_frame2_16_3
        );

    \I__12038\ : Odrv4
    port map (
            O => \N__48975\,
            I => data_out_frame2_16_3
        );

    \I__12037\ : LocalMux
    port map (
            O => \N__48972\,
            I => data_out_frame2_16_3
        );

    \I__12036\ : Odrv4
    port map (
            O => \N__48969\,
            I => data_out_frame2_16_3
        );

    \I__12035\ : Odrv4
    port map (
            O => \N__48966\,
            I => data_out_frame2_16_3
        );

    \I__12034\ : InMux
    port map (
            O => \N__48955\,
            I => \N__48952\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__48952\,
            I => \N__48949\
        );

    \I__12032\ : Span4Mux_h
    port map (
            O => \N__48949\,
            I => \N__48946\
        );

    \I__12031\ : Span4Mux_v
    port map (
            O => \N__48946\,
            I => \N__48943\
        );

    \I__12030\ : Odrv4
    port map (
            O => \N__48943\,
            I => \c0.n17948\
        );

    \I__12029\ : InMux
    port map (
            O => \N__48940\,
            I => \N__48937\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__48937\,
            I => \N__48931\
        );

    \I__12027\ : InMux
    port map (
            O => \N__48936\,
            I => \N__48928\
        );

    \I__12026\ : InMux
    port map (
            O => \N__48935\,
            I => \N__48925\
        );

    \I__12025\ : InMux
    port map (
            O => \N__48934\,
            I => \N__48922\
        );

    \I__12024\ : Span4Mux_v
    port map (
            O => \N__48931\,
            I => \N__48919\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__48928\,
            I => \N__48916\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__48925\,
            I => \N__48913\
        );

    \I__12021\ : LocalMux
    port map (
            O => \N__48922\,
            I => \N__48909\
        );

    \I__12020\ : Span4Mux_h
    port map (
            O => \N__48919\,
            I => \N__48906\
        );

    \I__12019\ : Span12Mux_v
    port map (
            O => \N__48916\,
            I => \N__48903\
        );

    \I__12018\ : Span4Mux_v
    port map (
            O => \N__48913\,
            I => \N__48900\
        );

    \I__12017\ : InMux
    port map (
            O => \N__48912\,
            I => \N__48897\
        );

    \I__12016\ : Span4Mux_s1_v
    port map (
            O => \N__48909\,
            I => \N__48894\
        );

    \I__12015\ : Odrv4
    port map (
            O => \N__48906\,
            I => rand_data_30
        );

    \I__12014\ : Odrv12
    port map (
            O => \N__48903\,
            I => rand_data_30
        );

    \I__12013\ : Odrv4
    port map (
            O => \N__48900\,
            I => rand_data_30
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__48897\,
            I => rand_data_30
        );

    \I__12011\ : Odrv4
    port map (
            O => \N__48894\,
            I => rand_data_30
        );

    \I__12010\ : InMux
    port map (
            O => \N__48883\,
            I => \N__48877\
        );

    \I__12009\ : InMux
    port map (
            O => \N__48882\,
            I => \N__48877\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__48877\,
            I => \N__48873\
        );

    \I__12007\ : InMux
    port map (
            O => \N__48876\,
            I => \N__48869\
        );

    \I__12006\ : Span4Mux_v
    port map (
            O => \N__48873\,
            I => \N__48866\
        );

    \I__12005\ : InMux
    port map (
            O => \N__48872\,
            I => \N__48862\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__48869\,
            I => \N__48859\
        );

    \I__12003\ : Sp12to4
    port map (
            O => \N__48866\,
            I => \N__48856\
        );

    \I__12002\ : InMux
    port map (
            O => \N__48865\,
            I => \N__48853\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__48862\,
            I => data_out_frame2_5_6
        );

    \I__12000\ : Odrv4
    port map (
            O => \N__48859\,
            I => data_out_frame2_5_6
        );

    \I__11999\ : Odrv12
    port map (
            O => \N__48856\,
            I => data_out_frame2_5_6
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__48853\,
            I => data_out_frame2_5_6
        );

    \I__11997\ : InMux
    port map (
            O => \N__48844\,
            I => \N__48841\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__48841\,
            I => \N__48836\
        );

    \I__11995\ : InMux
    port map (
            O => \N__48840\,
            I => \N__48833\
        );

    \I__11994\ : InMux
    port map (
            O => \N__48839\,
            I => \N__48830\
        );

    \I__11993\ : Span4Mux_h
    port map (
            O => \N__48836\,
            I => \N__48825\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__48833\,
            I => \N__48822\
        );

    \I__11991\ : LocalMux
    port map (
            O => \N__48830\,
            I => \N__48819\
        );

    \I__11990\ : InMux
    port map (
            O => \N__48829\,
            I => \N__48816\
        );

    \I__11989\ : InMux
    port map (
            O => \N__48828\,
            I => \N__48812\
        );

    \I__11988\ : Span4Mux_v
    port map (
            O => \N__48825\,
            I => \N__48809\
        );

    \I__11987\ : Span12Mux_v
    port map (
            O => \N__48822\,
            I => \N__48806\
        );

    \I__11986\ : Span4Mux_v
    port map (
            O => \N__48819\,
            I => \N__48803\
        );

    \I__11985\ : LocalMux
    port map (
            O => \N__48816\,
            I => \N__48800\
        );

    \I__11984\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48797\
        );

    \I__11983\ : LocalMux
    port map (
            O => \N__48812\,
            I => \N__48794\
        );

    \I__11982\ : Odrv4
    port map (
            O => \N__48809\,
            I => rand_data_11
        );

    \I__11981\ : Odrv12
    port map (
            O => \N__48806\,
            I => rand_data_11
        );

    \I__11980\ : Odrv4
    port map (
            O => \N__48803\,
            I => rand_data_11
        );

    \I__11979\ : Odrv4
    port map (
            O => \N__48800\,
            I => rand_data_11
        );

    \I__11978\ : LocalMux
    port map (
            O => \N__48797\,
            I => rand_data_11
        );

    \I__11977\ : Odrv12
    port map (
            O => \N__48794\,
            I => rand_data_11
        );

    \I__11976\ : InMux
    port map (
            O => \N__48781\,
            I => \N__48777\
        );

    \I__11975\ : InMux
    port map (
            O => \N__48780\,
            I => \N__48774\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__48777\,
            I => data_out_frame2_17_3
        );

    \I__11973\ : LocalMux
    port map (
            O => \N__48774\,
            I => data_out_frame2_17_3
        );

    \I__11972\ : InMux
    port map (
            O => \N__48769\,
            I => \N__48763\
        );

    \I__11971\ : InMux
    port map (
            O => \N__48768\,
            I => \N__48760\
        );

    \I__11970\ : InMux
    port map (
            O => \N__48767\,
            I => \N__48757\
        );

    \I__11969\ : InMux
    port map (
            O => \N__48766\,
            I => \N__48754\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__48763\,
            I => \N__48751\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__48760\,
            I => \N__48748\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__48757\,
            I => \N__48745\
        );

    \I__11965\ : LocalMux
    port map (
            O => \N__48754\,
            I => \N__48741\
        );

    \I__11964\ : Span4Mux_h
    port map (
            O => \N__48751\,
            I => \N__48738\
        );

    \I__11963\ : Span4Mux_v
    port map (
            O => \N__48748\,
            I => \N__48733\
        );

    \I__11962\ : Span4Mux_v
    port map (
            O => \N__48745\,
            I => \N__48733\
        );

    \I__11961\ : InMux
    port map (
            O => \N__48744\,
            I => \N__48729\
        );

    \I__11960\ : Span4Mux_v
    port map (
            O => \N__48741\,
            I => \N__48724\
        );

    \I__11959\ : Span4Mux_h
    port map (
            O => \N__48738\,
            I => \N__48724\
        );

    \I__11958\ : Span4Mux_h
    port map (
            O => \N__48733\,
            I => \N__48721\
        );

    \I__11957\ : InMux
    port map (
            O => \N__48732\,
            I => \N__48718\
        );

    \I__11956\ : LocalMux
    port map (
            O => \N__48729\,
            I => \N__48715\
        );

    \I__11955\ : Odrv4
    port map (
            O => \N__48724\,
            I => rand_data_8
        );

    \I__11954\ : Odrv4
    port map (
            O => \N__48721\,
            I => rand_data_8
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__48718\,
            I => rand_data_8
        );

    \I__11952\ : Odrv12
    port map (
            O => \N__48715\,
            I => rand_data_8
        );

    \I__11951\ : InMux
    port map (
            O => \N__48706\,
            I => \N__48702\
        );

    \I__11950\ : InMux
    port map (
            O => \N__48705\,
            I => \N__48698\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__48702\,
            I => \N__48695\
        );

    \I__11948\ : InMux
    port map (
            O => \N__48701\,
            I => \N__48691\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__48698\,
            I => \N__48688\
        );

    \I__11946\ : Span4Mux_h
    port map (
            O => \N__48695\,
            I => \N__48685\
        );

    \I__11945\ : InMux
    port map (
            O => \N__48694\,
            I => \N__48682\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__48691\,
            I => \N__48679\
        );

    \I__11943\ : Span4Mux_h
    port map (
            O => \N__48688\,
            I => \N__48676\
        );

    \I__11942\ : Odrv4
    port map (
            O => \N__48685\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__48682\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__11940\ : Odrv12
    port map (
            O => \N__48679\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__11939\ : Odrv4
    port map (
            O => \N__48676\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__11938\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48662\
        );

    \I__11937\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48659\
        );

    \I__11936\ : InMux
    port map (
            O => \N__48665\,
            I => \N__48656\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__48662\,
            I => \N__48642\
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__48659\,
            I => \N__48642\
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__48656\,
            I => \N__48642\
        );

    \I__11932\ : InMux
    port map (
            O => \N__48655\,
            I => \N__48631\
        );

    \I__11931\ : InMux
    port map (
            O => \N__48654\,
            I => \N__48631\
        );

    \I__11930\ : CascadeMux
    port map (
            O => \N__48653\,
            I => \N__48626\
        );

    \I__11929\ : InMux
    port map (
            O => \N__48652\,
            I => \N__48618\
        );

    \I__11928\ : InMux
    port map (
            O => \N__48651\,
            I => \N__48618\
        );

    \I__11927\ : InMux
    port map (
            O => \N__48650\,
            I => \N__48615\
        );

    \I__11926\ : CascadeMux
    port map (
            O => \N__48649\,
            I => \N__48611\
        );

    \I__11925\ : Span4Mux_v
    port map (
            O => \N__48642\,
            I => \N__48608\
        );

    \I__11924\ : InMux
    port map (
            O => \N__48641\,
            I => \N__48605\
        );

    \I__11923\ : InMux
    port map (
            O => \N__48640\,
            I => \N__48601\
        );

    \I__11922\ : InMux
    port map (
            O => \N__48639\,
            I => \N__48596\
        );

    \I__11921\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48596\
        );

    \I__11920\ : CascadeMux
    port map (
            O => \N__48637\,
            I => \N__48590\
        );

    \I__11919\ : CascadeMux
    port map (
            O => \N__48636\,
            I => \N__48587\
        );

    \I__11918\ : LocalMux
    port map (
            O => \N__48631\,
            I => \N__48575\
        );

    \I__11917\ : InMux
    port map (
            O => \N__48630\,
            I => \N__48572\
        );

    \I__11916\ : CascadeMux
    port map (
            O => \N__48629\,
            I => \N__48569\
        );

    \I__11915\ : InMux
    port map (
            O => \N__48626\,
            I => \N__48565\
        );

    \I__11914\ : InMux
    port map (
            O => \N__48625\,
            I => \N__48561\
        );

    \I__11913\ : InMux
    port map (
            O => \N__48624\,
            I => \N__48558\
        );

    \I__11912\ : InMux
    port map (
            O => \N__48623\,
            I => \N__48555\
        );

    \I__11911\ : LocalMux
    port map (
            O => \N__48618\,
            I => \N__48552\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__48615\,
            I => \N__48549\
        );

    \I__11909\ : InMux
    port map (
            O => \N__48614\,
            I => \N__48546\
        );

    \I__11908\ : InMux
    port map (
            O => \N__48611\,
            I => \N__48543\
        );

    \I__11907\ : Span4Mux_h
    port map (
            O => \N__48608\,
            I => \N__48536\
        );

    \I__11906\ : LocalMux
    port map (
            O => \N__48605\,
            I => \N__48536\
        );

    \I__11905\ : InMux
    port map (
            O => \N__48604\,
            I => \N__48532\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__48601\,
            I => \N__48527\
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__48596\,
            I => \N__48527\
        );

    \I__11902\ : InMux
    port map (
            O => \N__48595\,
            I => \N__48524\
        );

    \I__11901\ : InMux
    port map (
            O => \N__48594\,
            I => \N__48517\
        );

    \I__11900\ : InMux
    port map (
            O => \N__48593\,
            I => \N__48517\
        );

    \I__11899\ : InMux
    port map (
            O => \N__48590\,
            I => \N__48517\
        );

    \I__11898\ : InMux
    port map (
            O => \N__48587\,
            I => \N__48514\
        );

    \I__11897\ : InMux
    port map (
            O => \N__48586\,
            I => \N__48509\
        );

    \I__11896\ : InMux
    port map (
            O => \N__48585\,
            I => \N__48506\
        );

    \I__11895\ : InMux
    port map (
            O => \N__48584\,
            I => \N__48503\
        );

    \I__11894\ : CascadeMux
    port map (
            O => \N__48583\,
            I => \N__48500\
        );

    \I__11893\ : CascadeMux
    port map (
            O => \N__48582\,
            I => \N__48497\
        );

    \I__11892\ : CascadeMux
    port map (
            O => \N__48581\,
            I => \N__48494\
        );

    \I__11891\ : CascadeMux
    port map (
            O => \N__48580\,
            I => \N__48486\
        );

    \I__11890\ : InMux
    port map (
            O => \N__48579\,
            I => \N__48481\
        );

    \I__11889\ : InMux
    port map (
            O => \N__48578\,
            I => \N__48481\
        );

    \I__11888\ : Span4Mux_v
    port map (
            O => \N__48575\,
            I => \N__48478\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__48572\,
            I => \N__48475\
        );

    \I__11886\ : InMux
    port map (
            O => \N__48569\,
            I => \N__48472\
        );

    \I__11885\ : InMux
    port map (
            O => \N__48568\,
            I => \N__48469\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__48565\,
            I => \N__48466\
        );

    \I__11883\ : CascadeMux
    port map (
            O => \N__48564\,
            I => \N__48462\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__48561\,
            I => \N__48453\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__48558\,
            I => \N__48450\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__48555\,
            I => \N__48447\
        );

    \I__11879\ : Span4Mux_v
    port map (
            O => \N__48552\,
            I => \N__48438\
        );

    \I__11878\ : Span4Mux_v
    port map (
            O => \N__48549\,
            I => \N__48438\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__48546\,
            I => \N__48438\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__48543\,
            I => \N__48438\
        );

    \I__11875\ : InMux
    port map (
            O => \N__48542\,
            I => \N__48433\
        );

    \I__11874\ : InMux
    port map (
            O => \N__48541\,
            I => \N__48433\
        );

    \I__11873\ : Span4Mux_v
    port map (
            O => \N__48536\,
            I => \N__48430\
        );

    \I__11872\ : InMux
    port map (
            O => \N__48535\,
            I => \N__48427\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__48532\,
            I => \N__48418\
        );

    \I__11870\ : Span4Mux_v
    port map (
            O => \N__48527\,
            I => \N__48418\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__48524\,
            I => \N__48418\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__48517\,
            I => \N__48418\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__48514\,
            I => \N__48415\
        );

    \I__11866\ : InMux
    port map (
            O => \N__48513\,
            I => \N__48412\
        );

    \I__11865\ : InMux
    port map (
            O => \N__48512\,
            I => \N__48409\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__48509\,
            I => \N__48402\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__48506\,
            I => \N__48402\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__48503\,
            I => \N__48402\
        );

    \I__11861\ : InMux
    port map (
            O => \N__48500\,
            I => \N__48397\
        );

    \I__11860\ : InMux
    port map (
            O => \N__48497\,
            I => \N__48397\
        );

    \I__11859\ : InMux
    port map (
            O => \N__48494\,
            I => \N__48394\
        );

    \I__11858\ : InMux
    port map (
            O => \N__48493\,
            I => \N__48388\
        );

    \I__11857\ : InMux
    port map (
            O => \N__48492\,
            I => \N__48381\
        );

    \I__11856\ : InMux
    port map (
            O => \N__48491\,
            I => \N__48381\
        );

    \I__11855\ : InMux
    port map (
            O => \N__48490\,
            I => \N__48381\
        );

    \I__11854\ : InMux
    port map (
            O => \N__48489\,
            I => \N__48378\
        );

    \I__11853\ : InMux
    port map (
            O => \N__48486\,
            I => \N__48375\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__48481\,
            I => \N__48372\
        );

    \I__11851\ : Span4Mux_h
    port map (
            O => \N__48478\,
            I => \N__48365\
        );

    \I__11850\ : Span4Mux_h
    port map (
            O => \N__48475\,
            I => \N__48365\
        );

    \I__11849\ : LocalMux
    port map (
            O => \N__48472\,
            I => \N__48365\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__48469\,
            I => \N__48360\
        );

    \I__11847\ : Span4Mux_h
    port map (
            O => \N__48466\,
            I => \N__48360\
        );

    \I__11846\ : InMux
    port map (
            O => \N__48465\,
            I => \N__48355\
        );

    \I__11845\ : InMux
    port map (
            O => \N__48462\,
            I => \N__48355\
        );

    \I__11844\ : InMux
    port map (
            O => \N__48461\,
            I => \N__48350\
        );

    \I__11843\ : InMux
    port map (
            O => \N__48460\,
            I => \N__48341\
        );

    \I__11842\ : InMux
    port map (
            O => \N__48459\,
            I => \N__48341\
        );

    \I__11841\ : InMux
    port map (
            O => \N__48458\,
            I => \N__48341\
        );

    \I__11840\ : InMux
    port map (
            O => \N__48457\,
            I => \N__48341\
        );

    \I__11839\ : InMux
    port map (
            O => \N__48456\,
            I => \N__48338\
        );

    \I__11838\ : Span4Mux_v
    port map (
            O => \N__48453\,
            I => \N__48331\
        );

    \I__11837\ : Span4Mux_v
    port map (
            O => \N__48450\,
            I => \N__48331\
        );

    \I__11836\ : Span4Mux_v
    port map (
            O => \N__48447\,
            I => \N__48331\
        );

    \I__11835\ : Span4Mux_v
    port map (
            O => \N__48438\,
            I => \N__48328\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__48433\,
            I => \N__48323\
        );

    \I__11833\ : Span4Mux_v
    port map (
            O => \N__48430\,
            I => \N__48323\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__48427\,
            I => \N__48318\
        );

    \I__11831\ : Span4Mux_v
    port map (
            O => \N__48418\,
            I => \N__48318\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__48415\,
            I => \N__48315\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__48412\,
            I => \N__48304\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__48409\,
            I => \N__48304\
        );

    \I__11827\ : Span4Mux_v
    port map (
            O => \N__48402\,
            I => \N__48304\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__48397\,
            I => \N__48304\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__48394\,
            I => \N__48304\
        );

    \I__11824\ : InMux
    port map (
            O => \N__48393\,
            I => \N__48299\
        );

    \I__11823\ : InMux
    port map (
            O => \N__48392\,
            I => \N__48299\
        );

    \I__11822\ : InMux
    port map (
            O => \N__48391\,
            I => \N__48296\
        );

    \I__11821\ : LocalMux
    port map (
            O => \N__48388\,
            I => \N__48279\
        );

    \I__11820\ : LocalMux
    port map (
            O => \N__48381\,
            I => \N__48279\
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48279\
        );

    \I__11818\ : LocalMux
    port map (
            O => \N__48375\,
            I => \N__48279\
        );

    \I__11817\ : Span4Mux_h
    port map (
            O => \N__48372\,
            I => \N__48279\
        );

    \I__11816\ : Span4Mux_v
    port map (
            O => \N__48365\,
            I => \N__48279\
        );

    \I__11815\ : Span4Mux_h
    port map (
            O => \N__48360\,
            I => \N__48279\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__48355\,
            I => \N__48279\
        );

    \I__11813\ : InMux
    port map (
            O => \N__48354\,
            I => \N__48276\
        );

    \I__11812\ : InMux
    port map (
            O => \N__48353\,
            I => \N__48273\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__48350\,
            I => \N__48270\
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__48341\,
            I => \N__48265\
        );

    \I__11809\ : LocalMux
    port map (
            O => \N__48338\,
            I => \N__48265\
        );

    \I__11808\ : Span4Mux_h
    port map (
            O => \N__48331\,
            I => \N__48260\
        );

    \I__11807\ : Span4Mux_h
    port map (
            O => \N__48328\,
            I => \N__48260\
        );

    \I__11806\ : Span4Mux_v
    port map (
            O => \N__48323\,
            I => \N__48251\
        );

    \I__11805\ : Span4Mux_h
    port map (
            O => \N__48318\,
            I => \N__48251\
        );

    \I__11804\ : Span4Mux_h
    port map (
            O => \N__48315\,
            I => \N__48251\
        );

    \I__11803\ : Span4Mux_v
    port map (
            O => \N__48304\,
            I => \N__48251\
        );

    \I__11802\ : LocalMux
    port map (
            O => \N__48299\,
            I => \N__48244\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__48296\,
            I => \N__48244\
        );

    \I__11800\ : Sp12to4
    port map (
            O => \N__48279\,
            I => \N__48244\
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__48276\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__48273\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11797\ : Odrv12
    port map (
            O => \N__48270\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11796\ : Odrv4
    port map (
            O => \N__48265\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11795\ : Odrv4
    port map (
            O => \N__48260\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11794\ : Odrv4
    port map (
            O => \N__48251\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11793\ : Odrv12
    port map (
            O => \N__48244\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11792\ : InMux
    port map (
            O => \N__48229\,
            I => \N__48216\
        );

    \I__11791\ : InMux
    port map (
            O => \N__48228\,
            I => \N__48216\
        );

    \I__11790\ : InMux
    port map (
            O => \N__48227\,
            I => \N__48202\
        );

    \I__11789\ : InMux
    port map (
            O => \N__48226\,
            I => \N__48202\
        );

    \I__11788\ : InMux
    port map (
            O => \N__48225\,
            I => \N__48195\
        );

    \I__11787\ : InMux
    port map (
            O => \N__48224\,
            I => \N__48195\
        );

    \I__11786\ : InMux
    port map (
            O => \N__48223\,
            I => \N__48195\
        );

    \I__11785\ : CascadeMux
    port map (
            O => \N__48222\,
            I => \N__48191\
        );

    \I__11784\ : InMux
    port map (
            O => \N__48221\,
            I => \N__48183\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__48216\,
            I => \N__48180\
        );

    \I__11782\ : InMux
    port map (
            O => \N__48215\,
            I => \N__48177\
        );

    \I__11781\ : InMux
    port map (
            O => \N__48214\,
            I => \N__48172\
        );

    \I__11780\ : InMux
    port map (
            O => \N__48213\,
            I => \N__48172\
        );

    \I__11779\ : InMux
    port map (
            O => \N__48212\,
            I => \N__48168\
        );

    \I__11778\ : InMux
    port map (
            O => \N__48211\,
            I => \N__48161\
        );

    \I__11777\ : InMux
    port map (
            O => \N__48210\,
            I => \N__48154\
        );

    \I__11776\ : InMux
    port map (
            O => \N__48209\,
            I => \N__48154\
        );

    \I__11775\ : InMux
    port map (
            O => \N__48208\,
            I => \N__48154\
        );

    \I__11774\ : InMux
    port map (
            O => \N__48207\,
            I => \N__48151\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__48202\,
            I => \N__48146\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__48195\,
            I => \N__48146\
        );

    \I__11771\ : InMux
    port map (
            O => \N__48194\,
            I => \N__48143\
        );

    \I__11770\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48137\
        );

    \I__11769\ : InMux
    port map (
            O => \N__48190\,
            I => \N__48134\
        );

    \I__11768\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48131\
        );

    \I__11767\ : InMux
    port map (
            O => \N__48188\,
            I => \N__48128\
        );

    \I__11766\ : InMux
    port map (
            O => \N__48187\,
            I => \N__48125\
        );

    \I__11765\ : InMux
    port map (
            O => \N__48186\,
            I => \N__48122\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__48183\,
            I => \N__48111\
        );

    \I__11763\ : Span4Mux_v
    port map (
            O => \N__48180\,
            I => \N__48111\
        );

    \I__11762\ : LocalMux
    port map (
            O => \N__48177\,
            I => \N__48111\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__48172\,
            I => \N__48111\
        );

    \I__11760\ : InMux
    port map (
            O => \N__48171\,
            I => \N__48108\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__48168\,
            I => \N__48101\
        );

    \I__11758\ : InMux
    port map (
            O => \N__48167\,
            I => \N__48098\
        );

    \I__11757\ : InMux
    port map (
            O => \N__48166\,
            I => \N__48093\
        );

    \I__11756\ : InMux
    port map (
            O => \N__48165\,
            I => \N__48089\
        );

    \I__11755\ : InMux
    port map (
            O => \N__48164\,
            I => \N__48086\
        );

    \I__11754\ : LocalMux
    port map (
            O => \N__48161\,
            I => \N__48081\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__48154\,
            I => \N__48081\
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__48151\,
            I => \N__48074\
        );

    \I__11751\ : Span4Mux_v
    port map (
            O => \N__48146\,
            I => \N__48074\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__48143\,
            I => \N__48074\
        );

    \I__11749\ : InMux
    port map (
            O => \N__48142\,
            I => \N__48067\
        );

    \I__11748\ : InMux
    port map (
            O => \N__48141\,
            I => \N__48067\
        );

    \I__11747\ : InMux
    port map (
            O => \N__48140\,
            I => \N__48067\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__48137\,
            I => \N__48060\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__48134\,
            I => \N__48060\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__48131\,
            I => \N__48053\
        );

    \I__11743\ : LocalMux
    port map (
            O => \N__48128\,
            I => \N__48053\
        );

    \I__11742\ : LocalMux
    port map (
            O => \N__48125\,
            I => \N__48053\
        );

    \I__11741\ : LocalMux
    port map (
            O => \N__48122\,
            I => \N__48048\
        );

    \I__11740\ : InMux
    port map (
            O => \N__48121\,
            I => \N__48045\
        );

    \I__11739\ : InMux
    port map (
            O => \N__48120\,
            I => \N__48039\
        );

    \I__11738\ : Span4Mux_v
    port map (
            O => \N__48111\,
            I => \N__48034\
        );

    \I__11737\ : LocalMux
    port map (
            O => \N__48108\,
            I => \N__48034\
        );

    \I__11736\ : InMux
    port map (
            O => \N__48107\,
            I => \N__48031\
        );

    \I__11735\ : InMux
    port map (
            O => \N__48106\,
            I => \N__48027\
        );

    \I__11734\ : InMux
    port map (
            O => \N__48105\,
            I => \N__48024\
        );

    \I__11733\ : InMux
    port map (
            O => \N__48104\,
            I => \N__48021\
        );

    \I__11732\ : Span4Mux_h
    port map (
            O => \N__48101\,
            I => \N__48016\
        );

    \I__11731\ : LocalMux
    port map (
            O => \N__48098\,
            I => \N__48016\
        );

    \I__11730\ : InMux
    port map (
            O => \N__48097\,
            I => \N__48013\
        );

    \I__11729\ : CascadeMux
    port map (
            O => \N__48096\,
            I => \N__48010\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__48093\,
            I => \N__48006\
        );

    \I__11727\ : InMux
    port map (
            O => \N__48092\,
            I => \N__48003\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__48089\,
            I => \N__47998\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__48086\,
            I => \N__47998\
        );

    \I__11724\ : Span4Mux_h
    port map (
            O => \N__48081\,
            I => \N__47991\
        );

    \I__11723\ : Span4Mux_v
    port map (
            O => \N__48074\,
            I => \N__47991\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__48067\,
            I => \N__47991\
        );

    \I__11721\ : InMux
    port map (
            O => \N__48066\,
            I => \N__47988\
        );

    \I__11720\ : InMux
    port map (
            O => \N__48065\,
            I => \N__47985\
        );

    \I__11719\ : Span4Mux_h
    port map (
            O => \N__48060\,
            I => \N__47980\
        );

    \I__11718\ : Span4Mux_v
    port map (
            O => \N__48053\,
            I => \N__47980\
        );

    \I__11717\ : InMux
    port map (
            O => \N__48052\,
            I => \N__47977\
        );

    \I__11716\ : InMux
    port map (
            O => \N__48051\,
            I => \N__47974\
        );

    \I__11715\ : Span4Mux_h
    port map (
            O => \N__48048\,
            I => \N__47969\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__48045\,
            I => \N__47969\
        );

    \I__11713\ : InMux
    port map (
            O => \N__48044\,
            I => \N__47964\
        );

    \I__11712\ : InMux
    port map (
            O => \N__48043\,
            I => \N__47964\
        );

    \I__11711\ : InMux
    port map (
            O => \N__48042\,
            I => \N__47957\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__48039\,
            I => \N__47954\
        );

    \I__11709\ : Span4Mux_h
    port map (
            O => \N__48034\,
            I => \N__47949\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__48031\,
            I => \N__47949\
        );

    \I__11707\ : InMux
    port map (
            O => \N__48030\,
            I => \N__47946\
        );

    \I__11706\ : LocalMux
    port map (
            O => \N__48027\,
            I => \N__47943\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__48024\,
            I => \N__47938\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__48021\,
            I => \N__47938\
        );

    \I__11703\ : Span4Mux_v
    port map (
            O => \N__48016\,
            I => \N__47933\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__48013\,
            I => \N__47933\
        );

    \I__11701\ : InMux
    port map (
            O => \N__48010\,
            I => \N__47930\
        );

    \I__11700\ : InMux
    port map (
            O => \N__48009\,
            I => \N__47927\
        );

    \I__11699\ : Span4Mux_v
    port map (
            O => \N__48006\,
            I => \N__47924\
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__48003\,
            I => \N__47917\
        );

    \I__11697\ : Span4Mux_v
    port map (
            O => \N__47998\,
            I => \N__47917\
        );

    \I__11696\ : Span4Mux_h
    port map (
            O => \N__47991\,
            I => \N__47917\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__47988\,
            I => \N__47910\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__47985\,
            I => \N__47910\
        );

    \I__11693\ : Span4Mux_h
    port map (
            O => \N__47980\,
            I => \N__47910\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__47977\,
            I => \N__47901\
        );

    \I__11691\ : LocalMux
    port map (
            O => \N__47974\,
            I => \N__47901\
        );

    \I__11690\ : Span4Mux_v
    port map (
            O => \N__47969\,
            I => \N__47901\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__47964\,
            I => \N__47901\
        );

    \I__11688\ : InMux
    port map (
            O => \N__47963\,
            I => \N__47898\
        );

    \I__11687\ : InMux
    port map (
            O => \N__47962\,
            I => \N__47895\
        );

    \I__11686\ : InMux
    port map (
            O => \N__47961\,
            I => \N__47890\
        );

    \I__11685\ : InMux
    port map (
            O => \N__47960\,
            I => \N__47890\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__47957\,
            I => \N__47881\
        );

    \I__11683\ : Span4Mux_h
    port map (
            O => \N__47954\,
            I => \N__47881\
        );

    \I__11682\ : Span4Mux_v
    port map (
            O => \N__47949\,
            I => \N__47881\
        );

    \I__11681\ : LocalMux
    port map (
            O => \N__47946\,
            I => \N__47881\
        );

    \I__11680\ : Span4Mux_v
    port map (
            O => \N__47943\,
            I => \N__47874\
        );

    \I__11679\ : Span4Mux_v
    port map (
            O => \N__47938\,
            I => \N__47874\
        );

    \I__11678\ : Span4Mux_h
    port map (
            O => \N__47933\,
            I => \N__47874\
        );

    \I__11677\ : LocalMux
    port map (
            O => \N__47930\,
            I => \N__47865\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__47927\,
            I => \N__47865\
        );

    \I__11675\ : Span4Mux_h
    port map (
            O => \N__47924\,
            I => \N__47865\
        );

    \I__11674\ : Span4Mux_v
    port map (
            O => \N__47917\,
            I => \N__47865\
        );

    \I__11673\ : Span4Mux_v
    port map (
            O => \N__47910\,
            I => \N__47860\
        );

    \I__11672\ : Span4Mux_v
    port map (
            O => \N__47901\,
            I => \N__47860\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__47898\,
            I => \N__47855\
        );

    \I__11670\ : LocalMux
    port map (
            O => \N__47895\,
            I => \N__47855\
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__47890\,
            I => \N__47848\
        );

    \I__11668\ : Span4Mux_v
    port map (
            O => \N__47881\,
            I => \N__47848\
        );

    \I__11667\ : Span4Mux_h
    port map (
            O => \N__47874\,
            I => \N__47848\
        );

    \I__11666\ : Odrv4
    port map (
            O => \N__47865\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11665\ : Odrv4
    port map (
            O => \N__47860\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11664\ : Odrv12
    port map (
            O => \N__47855\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11663\ : Odrv4
    port map (
            O => \N__47848\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11662\ : InMux
    port map (
            O => \N__47839\,
            I => \N__47836\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__47836\,
            I => \N__47833\
        );

    \I__11660\ : Odrv4
    port map (
            O => \N__47833\,
            I => \c0.n17563\
        );

    \I__11659\ : InMux
    port map (
            O => \N__47830\,
            I => \N__47827\
        );

    \I__11658\ : LocalMux
    port map (
            O => \N__47827\,
            I => \N__47824\
        );

    \I__11657\ : Odrv4
    port map (
            O => \N__47824\,
            I => \c0.n17999\
        );

    \I__11656\ : InMux
    port map (
            O => \N__47821\,
            I => \N__47818\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__47818\,
            I => \N__47811\
        );

    \I__11654\ : InMux
    port map (
            O => \N__47817\,
            I => \N__47808\
        );

    \I__11653\ : InMux
    port map (
            O => \N__47816\,
            I => \N__47805\
        );

    \I__11652\ : InMux
    port map (
            O => \N__47815\,
            I => \N__47801\
        );

    \I__11651\ : InMux
    port map (
            O => \N__47814\,
            I => \N__47798\
        );

    \I__11650\ : Span4Mux_h
    port map (
            O => \N__47811\,
            I => \N__47791\
        );

    \I__11649\ : LocalMux
    port map (
            O => \N__47808\,
            I => \N__47791\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__47805\,
            I => \N__47791\
        );

    \I__11647\ : InMux
    port map (
            O => \N__47804\,
            I => \N__47788\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__47801\,
            I => \N__47784\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__47798\,
            I => \N__47781\
        );

    \I__11644\ : Span4Mux_v
    port map (
            O => \N__47791\,
            I => \N__47776\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__47788\,
            I => \N__47776\
        );

    \I__11642\ : InMux
    port map (
            O => \N__47787\,
            I => \N__47773\
        );

    \I__11641\ : Span4Mux_h
    port map (
            O => \N__47784\,
            I => \N__47770\
        );

    \I__11640\ : Span4Mux_h
    port map (
            O => \N__47781\,
            I => \N__47767\
        );

    \I__11639\ : Span4Mux_v
    port map (
            O => \N__47776\,
            I => \N__47762\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__47773\,
            I => \N__47762\
        );

    \I__11637\ : Span4Mux_h
    port map (
            O => \N__47770\,
            I => \N__47758\
        );

    \I__11636\ : Span4Mux_v
    port map (
            O => \N__47767\,
            I => \N__47755\
        );

    \I__11635\ : Span4Mux_h
    port map (
            O => \N__47762\,
            I => \N__47752\
        );

    \I__11634\ : InMux
    port map (
            O => \N__47761\,
            I => \N__47749\
        );

    \I__11633\ : Odrv4
    port map (
            O => \N__47758\,
            I => \c0.n8621\
        );

    \I__11632\ : Odrv4
    port map (
            O => \N__47755\,
            I => \c0.n8621\
        );

    \I__11631\ : Odrv4
    port map (
            O => \N__47752\,
            I => \c0.n8621\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__47749\,
            I => \c0.n8621\
        );

    \I__11629\ : InMux
    port map (
            O => \N__47740\,
            I => \N__47737\
        );

    \I__11628\ : LocalMux
    port map (
            O => \N__47737\,
            I => \c0.n18002\
        );

    \I__11627\ : CascadeMux
    port map (
            O => \N__47734\,
            I => \N__47731\
        );

    \I__11626\ : InMux
    port map (
            O => \N__47731\,
            I => \N__47728\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__47728\,
            I => \N__47725\
        );

    \I__11624\ : Span4Mux_v
    port map (
            O => \N__47725\,
            I => \N__47722\
        );

    \I__11623\ : Sp12to4
    port map (
            O => \N__47722\,
            I => \N__47719\
        );

    \I__11622\ : Odrv12
    port map (
            O => \N__47719\,
            I => \c0.data_out_frame2_20_6\
        );

    \I__11621\ : InMux
    port map (
            O => \N__47716\,
            I => \N__47702\
        );

    \I__11620\ : InMux
    port map (
            O => \N__47715\,
            I => \N__47699\
        );

    \I__11619\ : InMux
    port map (
            O => \N__47714\,
            I => \N__47696\
        );

    \I__11618\ : InMux
    port map (
            O => \N__47713\,
            I => \N__47693\
        );

    \I__11617\ : InMux
    port map (
            O => \N__47712\,
            I => \N__47690\
        );

    \I__11616\ : InMux
    port map (
            O => \N__47711\,
            I => \N__47687\
        );

    \I__11615\ : InMux
    port map (
            O => \N__47710\,
            I => \N__47684\
        );

    \I__11614\ : InMux
    port map (
            O => \N__47709\,
            I => \N__47681\
        );

    \I__11613\ : InMux
    port map (
            O => \N__47708\,
            I => \N__47678\
        );

    \I__11612\ : InMux
    port map (
            O => \N__47707\,
            I => \N__47675\
        );

    \I__11611\ : InMux
    port map (
            O => \N__47706\,
            I => \N__47671\
        );

    \I__11610\ : InMux
    port map (
            O => \N__47705\,
            I => \N__47668\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__47702\,
            I => \N__47661\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__47699\,
            I => \N__47661\
        );

    \I__11607\ : LocalMux
    port map (
            O => \N__47696\,
            I => \N__47661\
        );

    \I__11606\ : LocalMux
    port map (
            O => \N__47693\,
            I => \N__47651\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__47690\,
            I => \N__47651\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__47687\,
            I => \N__47651\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__47684\,
            I => \N__47646\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__47681\,
            I => \N__47646\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__47678\,
            I => \N__47639\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__47675\,
            I => \N__47636\
        );

    \I__11599\ : InMux
    port map (
            O => \N__47674\,
            I => \N__47633\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__47671\,
            I => \N__47624\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__47668\,
            I => \N__47624\
        );

    \I__11596\ : Span4Mux_v
    port map (
            O => \N__47661\,
            I => \N__47624\
        );

    \I__11595\ : InMux
    port map (
            O => \N__47660\,
            I => \N__47621\
        );

    \I__11594\ : InMux
    port map (
            O => \N__47659\,
            I => \N__47618\
        );

    \I__11593\ : InMux
    port map (
            O => \N__47658\,
            I => \N__47615\
        );

    \I__11592\ : Span4Mux_v
    port map (
            O => \N__47651\,
            I => \N__47612\
        );

    \I__11591\ : Span4Mux_h
    port map (
            O => \N__47646\,
            I => \N__47609\
        );

    \I__11590\ : InMux
    port map (
            O => \N__47645\,
            I => \N__47606\
        );

    \I__11589\ : InMux
    port map (
            O => \N__47644\,
            I => \N__47601\
        );

    \I__11588\ : InMux
    port map (
            O => \N__47643\,
            I => \N__47601\
        );

    \I__11587\ : InMux
    port map (
            O => \N__47642\,
            I => \N__47598\
        );

    \I__11586\ : Span4Mux_h
    port map (
            O => \N__47639\,
            I => \N__47595\
        );

    \I__11585\ : Span4Mux_h
    port map (
            O => \N__47636\,
            I => \N__47590\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__47633\,
            I => \N__47590\
        );

    \I__11583\ : InMux
    port map (
            O => \N__47632\,
            I => \N__47587\
        );

    \I__11582\ : InMux
    port map (
            O => \N__47631\,
            I => \N__47584\
        );

    \I__11581\ : Span4Mux_h
    port map (
            O => \N__47624\,
            I => \N__47579\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__47621\,
            I => \N__47579\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__47618\,
            I => \N__47569\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__47615\,
            I => \N__47569\
        );

    \I__11577\ : Span4Mux_v
    port map (
            O => \N__47612\,
            I => \N__47569\
        );

    \I__11576\ : Span4Mux_v
    port map (
            O => \N__47609\,
            I => \N__47569\
        );

    \I__11575\ : LocalMux
    port map (
            O => \N__47606\,
            I => \N__47560\
        );

    \I__11574\ : LocalMux
    port map (
            O => \N__47601\,
            I => \N__47560\
        );

    \I__11573\ : LocalMux
    port map (
            O => \N__47598\,
            I => \N__47560\
        );

    \I__11572\ : Span4Mux_h
    port map (
            O => \N__47595\,
            I => \N__47560\
        );

    \I__11571\ : Span4Mux_h
    port map (
            O => \N__47590\,
            I => \N__47557\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__47587\,
            I => \N__47550\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__47584\,
            I => \N__47550\
        );

    \I__11568\ : Sp12to4
    port map (
            O => \N__47579\,
            I => \N__47550\
        );

    \I__11567\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47547\
        );

    \I__11566\ : Odrv4
    port map (
            O => \N__47569\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11565\ : Odrv4
    port map (
            O => \N__47560\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11564\ : Odrv4
    port map (
            O => \N__47557\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11563\ : Odrv12
    port map (
            O => \N__47550\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__47547\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11561\ : InMux
    port map (
            O => \N__47536\,
            I => \N__47533\
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__47533\,
            I => \c0.n22_adj_2353\
        );

    \I__11559\ : InMux
    port map (
            O => \N__47530\,
            I => \N__47527\
        );

    \I__11558\ : LocalMux
    port map (
            O => \N__47527\,
            I => \N__47524\
        );

    \I__11557\ : Span12Mux_h
    port map (
            O => \N__47524\,
            I => \N__47521\
        );

    \I__11556\ : Odrv12
    port map (
            O => \N__47521\,
            I => \c0.tx2.r_Tx_Data_6\
        );

    \I__11555\ : InMux
    port map (
            O => \N__47518\,
            I => \N__47515\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__47515\,
            I => \N__47512\
        );

    \I__11553\ : Odrv4
    port map (
            O => \N__47512\,
            I => \c0.n16915\
        );

    \I__11552\ : InMux
    port map (
            O => \N__47509\,
            I => \N__47506\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__47506\,
            I => \N__47502\
        );

    \I__11550\ : InMux
    port map (
            O => \N__47505\,
            I => \N__47499\
        );

    \I__11549\ : Span4Mux_h
    port map (
            O => \N__47502\,
            I => \N__47496\
        );

    \I__11548\ : LocalMux
    port map (
            O => \N__47499\,
            I => \N__47493\
        );

    \I__11547\ : Odrv4
    port map (
            O => \N__47496\,
            I => \c0.n17082\
        );

    \I__11546\ : Odrv4
    port map (
            O => \N__47493\,
            I => \c0.n17082\
        );

    \I__11545\ : CascadeMux
    port map (
            O => \N__47488\,
            I => \N__47485\
        );

    \I__11544\ : InMux
    port map (
            O => \N__47485\,
            I => \N__47481\
        );

    \I__11543\ : CascadeMux
    port map (
            O => \N__47484\,
            I => \N__47478\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__47481\,
            I => \N__47475\
        );

    \I__11541\ : InMux
    port map (
            O => \N__47478\,
            I => \N__47472\
        );

    \I__11540\ : Span4Mux_h
    port map (
            O => \N__47475\,
            I => \N__47467\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__47472\,
            I => \N__47467\
        );

    \I__11538\ : Span4Mux_h
    port map (
            O => \N__47467\,
            I => \N__47464\
        );

    \I__11537\ : Span4Mux_h
    port map (
            O => \N__47464\,
            I => \N__47461\
        );

    \I__11536\ : Odrv4
    port map (
            O => \N__47461\,
            I => \c0.n17118\
        );

    \I__11535\ : InMux
    port map (
            O => \N__47458\,
            I => \N__47455\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__47455\,
            I => \N__47452\
        );

    \I__11533\ : Span4Mux_v
    port map (
            O => \N__47452\,
            I => \N__47448\
        );

    \I__11532\ : InMux
    port map (
            O => \N__47451\,
            I => \N__47445\
        );

    \I__11531\ : Odrv4
    port map (
            O => \N__47448\,
            I => \c0.n17019\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__47445\,
            I => \c0.n17019\
        );

    \I__11529\ : CascadeMux
    port map (
            O => \N__47440\,
            I => \N__47437\
        );

    \I__11528\ : InMux
    port map (
            O => \N__47437\,
            I => \N__47434\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__47434\,
            I => \c0.n5_adj_2321\
        );

    \I__11526\ : InMux
    port map (
            O => \N__47431\,
            I => \N__47428\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__47428\,
            I => \c0.n18083\
        );

    \I__11524\ : CascadeMux
    port map (
            O => \N__47425\,
            I => \c0.n6_adj_2290_cascade_\
        );

    \I__11523\ : InMux
    port map (
            O => \N__47422\,
            I => \N__47419\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__47419\,
            I => \c0.n18086\
        );

    \I__11521\ : InMux
    port map (
            O => \N__47416\,
            I => \N__47412\
        );

    \I__11520\ : InMux
    port map (
            O => \N__47415\,
            I => \N__47406\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__47412\,
            I => \N__47403\
        );

    \I__11518\ : InMux
    port map (
            O => \N__47411\,
            I => \N__47398\
        );

    \I__11517\ : InMux
    port map (
            O => \N__47410\,
            I => \N__47398\
        );

    \I__11516\ : InMux
    port map (
            O => \N__47409\,
            I => \N__47395\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__47406\,
            I => \N__47392\
        );

    \I__11514\ : Span4Mux_v
    port map (
            O => \N__47403\,
            I => \N__47389\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__47398\,
            I => \N__47386\
        );

    \I__11512\ : LocalMux
    port map (
            O => \N__47395\,
            I => data_out_frame2_10_1
        );

    \I__11511\ : Odrv4
    port map (
            O => \N__47392\,
            I => data_out_frame2_10_1
        );

    \I__11510\ : Odrv4
    port map (
            O => \N__47389\,
            I => data_out_frame2_10_1
        );

    \I__11509\ : Odrv4
    port map (
            O => \N__47386\,
            I => data_out_frame2_10_1
        );

    \I__11508\ : InMux
    port map (
            O => \N__47377\,
            I => \N__47373\
        );

    \I__11507\ : InMux
    port map (
            O => \N__47376\,
            I => \N__47368\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__47373\,
            I => \N__47365\
        );

    \I__11505\ : InMux
    port map (
            O => \N__47372\,
            I => \N__47362\
        );

    \I__11504\ : InMux
    port map (
            O => \N__47371\,
            I => \N__47357\
        );

    \I__11503\ : LocalMux
    port map (
            O => \N__47368\,
            I => \N__47354\
        );

    \I__11502\ : Span4Mux_v
    port map (
            O => \N__47365\,
            I => \N__47351\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__47362\,
            I => \N__47348\
        );

    \I__11500\ : InMux
    port map (
            O => \N__47361\,
            I => \N__47345\
        );

    \I__11499\ : InMux
    port map (
            O => \N__47360\,
            I => \N__47342\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__47357\,
            I => \N__47339\
        );

    \I__11497\ : Span4Mux_v
    port map (
            O => \N__47354\,
            I => \N__47332\
        );

    \I__11496\ : Span4Mux_h
    port map (
            O => \N__47351\,
            I => \N__47332\
        );

    \I__11495\ : Span4Mux_v
    port map (
            O => \N__47348\,
            I => \N__47332\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__47345\,
            I => \N__47329\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__47342\,
            I => data_out_frame2_12_0
        );

    \I__11492\ : Odrv4
    port map (
            O => \N__47339\,
            I => data_out_frame2_12_0
        );

    \I__11491\ : Odrv4
    port map (
            O => \N__47332\,
            I => data_out_frame2_12_0
        );

    \I__11490\ : Odrv12
    port map (
            O => \N__47329\,
            I => data_out_frame2_12_0
        );

    \I__11489\ : CascadeMux
    port map (
            O => \N__47320\,
            I => \N__47317\
        );

    \I__11488\ : InMux
    port map (
            O => \N__47317\,
            I => \N__47314\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__47314\,
            I => \N__47309\
        );

    \I__11486\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47306\
        );

    \I__11485\ : CascadeMux
    port map (
            O => \N__47312\,
            I => \N__47303\
        );

    \I__11484\ : Span4Mux_h
    port map (
            O => \N__47309\,
            I => \N__47296\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__47306\,
            I => \N__47296\
        );

    \I__11482\ : InMux
    port map (
            O => \N__47303\,
            I => \N__47293\
        );

    \I__11481\ : CascadeMux
    port map (
            O => \N__47302\,
            I => \N__47290\
        );

    \I__11480\ : InMux
    port map (
            O => \N__47301\,
            I => \N__47287\
        );

    \I__11479\ : Span4Mux_v
    port map (
            O => \N__47296\,
            I => \N__47282\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__47293\,
            I => \N__47282\
        );

    \I__11477\ : InMux
    port map (
            O => \N__47290\,
            I => \N__47279\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__47287\,
            I => \N__47276\
        );

    \I__11475\ : Span4Mux_h
    port map (
            O => \N__47282\,
            I => \N__47271\
        );

    \I__11474\ : LocalMux
    port map (
            O => \N__47279\,
            I => \N__47271\
        );

    \I__11473\ : Span4Mux_h
    port map (
            O => \N__47276\,
            I => \N__47267\
        );

    \I__11472\ : Span4Mux_v
    port map (
            O => \N__47271\,
            I => \N__47264\
        );

    \I__11471\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47261\
        );

    \I__11470\ : Span4Mux_h
    port map (
            O => \N__47267\,
            I => \N__47258\
        );

    \I__11469\ : Span4Mux_h
    port map (
            O => \N__47264\,
            I => \N__47255\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__47261\,
            I => data_out_frame2_8_1
        );

    \I__11467\ : Odrv4
    port map (
            O => \N__47258\,
            I => data_out_frame2_8_1
        );

    \I__11466\ : Odrv4
    port map (
            O => \N__47255\,
            I => data_out_frame2_8_1
        );

    \I__11465\ : CascadeMux
    port map (
            O => \N__47248\,
            I => \N__47244\
        );

    \I__11464\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47241\
        );

    \I__11463\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47238\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__47241\,
            I => \N__47232\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__47238\,
            I => \N__47232\
        );

    \I__11460\ : InMux
    port map (
            O => \N__47237\,
            I => \N__47228\
        );

    \I__11459\ : Span4Mux_h
    port map (
            O => \N__47232\,
            I => \N__47225\
        );

    \I__11458\ : InMux
    port map (
            O => \N__47231\,
            I => \N__47221\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__47228\,
            I => \N__47216\
        );

    \I__11456\ : Span4Mux_h
    port map (
            O => \N__47225\,
            I => \N__47216\
        );

    \I__11455\ : InMux
    port map (
            O => \N__47224\,
            I => \N__47213\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__47221\,
            I => \N__47210\
        );

    \I__11453\ : Odrv4
    port map (
            O => \N__47216\,
            I => data_out_frame2_14_3
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__47213\,
            I => data_out_frame2_14_3
        );

    \I__11451\ : Odrv4
    port map (
            O => \N__47210\,
            I => data_out_frame2_14_3
        );

    \I__11450\ : CascadeMux
    port map (
            O => \N__47203\,
            I => \c0.n9895_cascade_\
        );

    \I__11449\ : InMux
    port map (
            O => \N__47200\,
            I => \N__47195\
        );

    \I__11448\ : InMux
    port map (
            O => \N__47199\,
            I => \N__47192\
        );

    \I__11447\ : InMux
    port map (
            O => \N__47198\,
            I => \N__47189\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__47195\,
            I => \N__47185\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__47192\,
            I => \N__47182\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__47189\,
            I => \N__47178\
        );

    \I__11443\ : InMux
    port map (
            O => \N__47188\,
            I => \N__47175\
        );

    \I__11442\ : Span4Mux_h
    port map (
            O => \N__47185\,
            I => \N__47172\
        );

    \I__11441\ : Span12Mux_h
    port map (
            O => \N__47182\,
            I => \N__47169\
        );

    \I__11440\ : InMux
    port map (
            O => \N__47181\,
            I => \N__47166\
        );

    \I__11439\ : Span12Mux_s9_v
    port map (
            O => \N__47178\,
            I => \N__47163\
        );

    \I__11438\ : LocalMux
    port map (
            O => \N__47175\,
            I => data_out_frame2_15_1
        );

    \I__11437\ : Odrv4
    port map (
            O => \N__47172\,
            I => data_out_frame2_15_1
        );

    \I__11436\ : Odrv12
    port map (
            O => \N__47169\,
            I => data_out_frame2_15_1
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__47166\,
            I => data_out_frame2_15_1
        );

    \I__11434\ : Odrv12
    port map (
            O => \N__47163\,
            I => data_out_frame2_15_1
        );

    \I__11433\ : CascadeMux
    port map (
            O => \N__47152\,
            I => \N__47149\
        );

    \I__11432\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47146\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__47146\,
            I => \N__47143\
        );

    \I__11430\ : Odrv4
    port map (
            O => \N__47143\,
            I => \c0.n6_adj_2274\
        );

    \I__11429\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47135\
        );

    \I__11428\ : InMux
    port map (
            O => \N__47139\,
            I => \N__47132\
        );

    \I__11427\ : InMux
    port map (
            O => \N__47138\,
            I => \N__47129\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__47135\,
            I => \N__47126\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__47132\,
            I => \N__47123\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__47129\,
            I => \N__47120\
        );

    \I__11423\ : Span4Mux_v
    port map (
            O => \N__47126\,
            I => \N__47117\
        );

    \I__11422\ : Span4Mux_v
    port map (
            O => \N__47123\,
            I => \N__47112\
        );

    \I__11421\ : Span4Mux_h
    port map (
            O => \N__47120\,
            I => \N__47112\
        );

    \I__11420\ : Span4Mux_h
    port map (
            O => \N__47117\,
            I => \N__47109\
        );

    \I__11419\ : Span4Mux_h
    port map (
            O => \N__47112\,
            I => \N__47106\
        );

    \I__11418\ : Odrv4
    port map (
            O => \N__47109\,
            I => \c0.data_out_9_4\
        );

    \I__11417\ : Odrv4
    port map (
            O => \N__47106\,
            I => \c0.data_out_9_4\
        );

    \I__11416\ : CascadeMux
    port map (
            O => \N__47101\,
            I => \N__47098\
        );

    \I__11415\ : InMux
    port map (
            O => \N__47098\,
            I => \N__47093\
        );

    \I__11414\ : InMux
    port map (
            O => \N__47097\,
            I => \N__47090\
        );

    \I__11413\ : InMux
    port map (
            O => \N__47096\,
            I => \N__47087\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__47093\,
            I => \N__47084\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__47090\,
            I => \N__47081\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__47087\,
            I => \N__47078\
        );

    \I__11409\ : Span4Mux_h
    port map (
            O => \N__47084\,
            I => \N__47075\
        );

    \I__11408\ : Span4Mux_v
    port map (
            O => \N__47081\,
            I => \N__47072\
        );

    \I__11407\ : Span4Mux_v
    port map (
            O => \N__47078\,
            I => \N__47069\
        );

    \I__11406\ : Span4Mux_v
    port map (
            O => \N__47075\,
            I => \N__47064\
        );

    \I__11405\ : Span4Mux_h
    port map (
            O => \N__47072\,
            I => \N__47064\
        );

    \I__11404\ : Span4Mux_h
    port map (
            O => \N__47069\,
            I => \N__47061\
        );

    \I__11403\ : Odrv4
    port map (
            O => \N__47064\,
            I => \c0.data_out_10_4\
        );

    \I__11402\ : Odrv4
    port map (
            O => \N__47061\,
            I => \c0.data_out_10_4\
        );

    \I__11401\ : InMux
    port map (
            O => \N__47056\,
            I => \N__47053\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__47053\,
            I => \N__47050\
        );

    \I__11399\ : Span4Mux_h
    port map (
            O => \N__47050\,
            I => \N__47046\
        );

    \I__11398\ : CascadeMux
    port map (
            O => \N__47049\,
            I => \N__47042\
        );

    \I__11397\ : Span4Mux_h
    port map (
            O => \N__47046\,
            I => \N__47039\
        );

    \I__11396\ : InMux
    port map (
            O => \N__47045\,
            I => \N__47034\
        );

    \I__11395\ : InMux
    port map (
            O => \N__47042\,
            I => \N__47034\
        );

    \I__11394\ : Odrv4
    port map (
            O => \N__47039\,
            I => \c0.data_out_7_2\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__47034\,
            I => \c0.data_out_7_2\
        );

    \I__11392\ : InMux
    port map (
            O => \N__47029\,
            I => \N__47026\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__47026\,
            I => \c0.n17058\
        );

    \I__11390\ : InMux
    port map (
            O => \N__47023\,
            I => \N__47019\
        );

    \I__11389\ : InMux
    port map (
            O => \N__47022\,
            I => \N__47016\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__47019\,
            I => \c0.n17028\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__47016\,
            I => \c0.n17028\
        );

    \I__11386\ : CascadeMux
    port map (
            O => \N__47011\,
            I => \c0.n17058_cascade_\
        );

    \I__11385\ : InMux
    port map (
            O => \N__47008\,
            I => \N__47005\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__47005\,
            I => \N__47001\
        );

    \I__11383\ : InMux
    port map (
            O => \N__47004\,
            I => \N__46998\
        );

    \I__11382\ : Odrv4
    port map (
            O => \N__47001\,
            I => \c0.n17094\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__46998\,
            I => \c0.n17094\
        );

    \I__11380\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46990\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__46990\,
            I => \N__46987\
        );

    \I__11378\ : Odrv4
    port map (
            O => \N__46987\,
            I => \c0.n19_adj_2283\
        );

    \I__11377\ : CascadeMux
    port map (
            O => \N__46984\,
            I => \c0.n21_adj_2284_cascade_\
        );

    \I__11376\ : InMux
    port map (
            O => \N__46981\,
            I => \N__46978\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__46978\,
            I => \N__46975\
        );

    \I__11374\ : Span4Mux_h
    port map (
            O => \N__46975\,
            I => \N__46972\
        );

    \I__11373\ : Odrv4
    port map (
            O => \N__46972\,
            I => \c0.n20_adj_2282\
        );

    \I__11372\ : InMux
    port map (
            O => \N__46969\,
            I => \N__46963\
        );

    \I__11371\ : InMux
    port map (
            O => \N__46968\,
            I => \N__46960\
        );

    \I__11370\ : InMux
    port map (
            O => \N__46967\,
            I => \N__46955\
        );

    \I__11369\ : InMux
    port map (
            O => \N__46966\,
            I => \N__46955\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__46963\,
            I => \N__46952\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__46960\,
            I => \N__46949\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__46955\,
            I => \N__46946\
        );

    \I__11365\ : Span4Mux_s3_v
    port map (
            O => \N__46952\,
            I => \N__46943\
        );

    \I__11364\ : Span4Mux_h
    port map (
            O => \N__46949\,
            I => \N__46940\
        );

    \I__11363\ : Span4Mux_h
    port map (
            O => \N__46946\,
            I => \N__46937\
        );

    \I__11362\ : Span4Mux_h
    port map (
            O => \N__46943\,
            I => \N__46934\
        );

    \I__11361\ : Odrv4
    port map (
            O => \N__46940\,
            I => \c0.data_out_9_7\
        );

    \I__11360\ : Odrv4
    port map (
            O => \N__46937\,
            I => \c0.data_out_9_7\
        );

    \I__11359\ : Odrv4
    port map (
            O => \N__46934\,
            I => \c0.data_out_9_7\
        );

    \I__11358\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46921\
        );

    \I__11357\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46921\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__46921\,
            I => \N__46918\
        );

    \I__11355\ : Span4Mux_h
    port map (
            O => \N__46918\,
            I => \N__46915\
        );

    \I__11354\ : Odrv4
    port map (
            O => \N__46915\,
            I => \c0.n17007\
        );

    \I__11353\ : InMux
    port map (
            O => \N__46912\,
            I => \N__46908\
        );

    \I__11352\ : InMux
    port map (
            O => \N__46911\,
            I => \N__46905\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__46908\,
            I => \N__46902\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__46905\,
            I => \N__46899\
        );

    \I__11349\ : Span4Mux_h
    port map (
            O => \N__46902\,
            I => \N__46895\
        );

    \I__11348\ : Span4Mux_h
    port map (
            O => \N__46899\,
            I => \N__46892\
        );

    \I__11347\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46889\
        );

    \I__11346\ : Odrv4
    port map (
            O => \N__46895\,
            I => \c0.n9505\
        );

    \I__11345\ : Odrv4
    port map (
            O => \N__46892\,
            I => \c0.n9505\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__46889\,
            I => \c0.n9505\
        );

    \I__11343\ : CascadeMux
    port map (
            O => \N__46882\,
            I => \N__46879\
        );

    \I__11342\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46875\
        );

    \I__11341\ : InMux
    port map (
            O => \N__46878\,
            I => \N__46872\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__46875\,
            I => \c0.n17076\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__46872\,
            I => \c0.n17076\
        );

    \I__11338\ : InMux
    port map (
            O => \N__46867\,
            I => \N__46864\
        );

    \I__11337\ : LocalMux
    port map (
            O => \N__46864\,
            I => \N__46860\
        );

    \I__11336\ : InMux
    port map (
            O => \N__46863\,
            I => \N__46857\
        );

    \I__11335\ : Span4Mux_h
    port map (
            O => \N__46860\,
            I => \N__46848\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__46857\,
            I => \N__46848\
        );

    \I__11333\ : InMux
    port map (
            O => \N__46856\,
            I => \N__46845\
        );

    \I__11332\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46842\
        );

    \I__11331\ : InMux
    port map (
            O => \N__46854\,
            I => \N__46839\
        );

    \I__11330\ : InMux
    port map (
            O => \N__46853\,
            I => \N__46836\
        );

    \I__11329\ : Span4Mux_h
    port map (
            O => \N__46848\,
            I => \N__46831\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__46845\,
            I => \N__46831\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__46842\,
            I => data_out_8_0
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__46839\,
            I => data_out_8_0
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__46836\,
            I => data_out_8_0
        );

    \I__11324\ : Odrv4
    port map (
            O => \N__46831\,
            I => data_out_8_0
        );

    \I__11323\ : InMux
    port map (
            O => \N__46822\,
            I => \N__46817\
        );

    \I__11322\ : InMux
    port map (
            O => \N__46821\,
            I => \N__46812\
        );

    \I__11321\ : InMux
    port map (
            O => \N__46820\,
            I => \N__46812\
        );

    \I__11320\ : LocalMux
    port map (
            O => \N__46817\,
            I => \N__46809\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__46812\,
            I => \c0.data_out_10_3\
        );

    \I__11318\ : Odrv12
    port map (
            O => \N__46809\,
            I => \c0.data_out_10_3\
        );

    \I__11317\ : InMux
    port map (
            O => \N__46804\,
            I => \N__46800\
        );

    \I__11316\ : InMux
    port map (
            O => \N__46803\,
            I => \N__46795\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__46800\,
            I => \N__46792\
        );

    \I__11314\ : InMux
    port map (
            O => \N__46799\,
            I => \N__46788\
        );

    \I__11313\ : InMux
    port map (
            O => \N__46798\,
            I => \N__46785\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__46795\,
            I => \N__46780\
        );

    \I__11311\ : Span4Mux_v
    port map (
            O => \N__46792\,
            I => \N__46780\
        );

    \I__11310\ : InMux
    port map (
            O => \N__46791\,
            I => \N__46777\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__46788\,
            I => \N__46772\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__46785\,
            I => \N__46772\
        );

    \I__11307\ : Span4Mux_h
    port map (
            O => \N__46780\,
            I => \N__46769\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__46777\,
            I => \N__46766\
        );

    \I__11305\ : Span4Mux_h
    port map (
            O => \N__46772\,
            I => \N__46763\
        );

    \I__11304\ : Odrv4
    port map (
            O => \N__46769\,
            I => \c0.data_out_9_6\
        );

    \I__11303\ : Odrv4
    port map (
            O => \N__46766\,
            I => \c0.data_out_9_6\
        );

    \I__11302\ : Odrv4
    port map (
            O => \N__46763\,
            I => \c0.data_out_9_6\
        );

    \I__11301\ : InMux
    port map (
            O => \N__46756\,
            I => \N__46752\
        );

    \I__11300\ : InMux
    port map (
            O => \N__46755\,
            I => \N__46749\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__46752\,
            I => \N__46746\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__46749\,
            I => \N__46743\
        );

    \I__11297\ : Span4Mux_s2_v
    port map (
            O => \N__46746\,
            I => \N__46740\
        );

    \I__11296\ : Span4Mux_h
    port map (
            O => \N__46743\,
            I => \N__46734\
        );

    \I__11295\ : Span4Mux_h
    port map (
            O => \N__46740\,
            I => \N__46734\
        );

    \I__11294\ : InMux
    port map (
            O => \N__46739\,
            I => \N__46731\
        );

    \I__11293\ : Odrv4
    port map (
            O => \N__46734\,
            I => \c0.data_out_10_2\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__46731\,
            I => \c0.data_out_10_2\
        );

    \I__11291\ : CascadeMux
    port map (
            O => \N__46726\,
            I => \N__46723\
        );

    \I__11290\ : InMux
    port map (
            O => \N__46723\,
            I => \N__46720\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__46720\,
            I => \N__46716\
        );

    \I__11288\ : InMux
    port map (
            O => \N__46719\,
            I => \N__46713\
        );

    \I__11287\ : Span4Mux_h
    port map (
            O => \N__46716\,
            I => \N__46710\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__46713\,
            I => \N__46707\
        );

    \I__11285\ : Odrv4
    port map (
            O => \N__46710\,
            I => \c0.n16998\
        );

    \I__11284\ : Odrv4
    port map (
            O => \N__46707\,
            I => \c0.n16998\
        );

    \I__11283\ : CascadeMux
    port map (
            O => \N__46702\,
            I => \N__46698\
        );

    \I__11282\ : InMux
    port map (
            O => \N__46701\,
            I => \N__46694\
        );

    \I__11281\ : InMux
    port map (
            O => \N__46698\,
            I => \N__46691\
        );

    \I__11280\ : InMux
    port map (
            O => \N__46697\,
            I => \N__46686\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__46694\,
            I => \N__46683\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__46691\,
            I => \N__46680\
        );

    \I__11277\ : InMux
    port map (
            O => \N__46690\,
            I => \N__46677\
        );

    \I__11276\ : InMux
    port map (
            O => \N__46689\,
            I => \N__46674\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__46686\,
            I => \N__46671\
        );

    \I__11274\ : Span4Mux_v
    port map (
            O => \N__46683\,
            I => \N__46664\
        );

    \I__11273\ : Span4Mux_v
    port map (
            O => \N__46680\,
            I => \N__46664\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__46677\,
            I => \N__46664\
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__46674\,
            I => \N__46661\
        );

    \I__11270\ : Odrv4
    port map (
            O => \N__46671\,
            I => \c0.data_out_6_2\
        );

    \I__11269\ : Odrv4
    port map (
            O => \N__46664\,
            I => \c0.data_out_6_2\
        );

    \I__11268\ : Odrv4
    port map (
            O => \N__46661\,
            I => \c0.data_out_6_2\
        );

    \I__11267\ : InMux
    port map (
            O => \N__46654\,
            I => \N__46651\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__46651\,
            I => \N__46648\
        );

    \I__11265\ : Span4Mux_v
    port map (
            O => \N__46648\,
            I => \N__46643\
        );

    \I__11264\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46640\
        );

    \I__11263\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46637\
        );

    \I__11262\ : Span4Mux_h
    port map (
            O => \N__46643\,
            I => \N__46630\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__46640\,
            I => \N__46630\
        );

    \I__11260\ : LocalMux
    port map (
            O => \N__46637\,
            I => \N__46630\
        );

    \I__11259\ : Span4Mux_v
    port map (
            O => \N__46630\,
            I => \N__46627\
        );

    \I__11258\ : Odrv4
    port map (
            O => \N__46627\,
            I => \c0.data_out_10_6\
        );

    \I__11257\ : CEMux
    port map (
            O => \N__46624\,
            I => \N__46617\
        );

    \I__11256\ : CEMux
    port map (
            O => \N__46623\,
            I => \N__46613\
        );

    \I__11255\ : CEMux
    port map (
            O => \N__46622\,
            I => \N__46610\
        );

    \I__11254\ : CEMux
    port map (
            O => \N__46621\,
            I => \N__46607\
        );

    \I__11253\ : CEMux
    port map (
            O => \N__46620\,
            I => \N__46603\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46600\
        );

    \I__11251\ : CEMux
    port map (
            O => \N__46616\,
            I => \N__46597\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__46613\,
            I => \N__46590\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__46610\,
            I => \N__46590\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__46607\,
            I => \N__46590\
        );

    \I__11247\ : CEMux
    port map (
            O => \N__46606\,
            I => \N__46586\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__46603\,
            I => \N__46583\
        );

    \I__11245\ : Span4Mux_v
    port map (
            O => \N__46600\,
            I => \N__46580\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__46597\,
            I => \N__46577\
        );

    \I__11243\ : Span4Mux_v
    port map (
            O => \N__46590\,
            I => \N__46574\
        );

    \I__11242\ : CEMux
    port map (
            O => \N__46589\,
            I => \N__46571\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__46586\,
            I => \N__46568\
        );

    \I__11240\ : Span4Mux_h
    port map (
            O => \N__46583\,
            I => \N__46564\
        );

    \I__11239\ : Span4Mux_h
    port map (
            O => \N__46580\,
            I => \N__46555\
        );

    \I__11238\ : Span4Mux_h
    port map (
            O => \N__46577\,
            I => \N__46555\
        );

    \I__11237\ : Span4Mux_h
    port map (
            O => \N__46574\,
            I => \N__46555\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__46571\,
            I => \N__46555\
        );

    \I__11235\ : IoSpan4Mux
    port map (
            O => \N__46568\,
            I => \N__46552\
        );

    \I__11234\ : InMux
    port map (
            O => \N__46567\,
            I => \N__46549\
        );

    \I__11233\ : Span4Mux_h
    port map (
            O => \N__46564\,
            I => \N__46546\
        );

    \I__11232\ : Span4Mux_h
    port map (
            O => \N__46555\,
            I => \N__46543\
        );

    \I__11231\ : IoSpan4Mux
    port map (
            O => \N__46552\,
            I => \N__46540\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__46549\,
            I => \N__46537\
        );

    \I__11229\ : Span4Mux_h
    port map (
            O => \N__46546\,
            I => \N__46534\
        );

    \I__11228\ : Span4Mux_v
    port map (
            O => \N__46543\,
            I => \N__46531\
        );

    \I__11227\ : IoSpan4Mux
    port map (
            O => \N__46540\,
            I => \N__46526\
        );

    \I__11226\ : Span4Mux_h
    port map (
            O => \N__46537\,
            I => \N__46526\
        );

    \I__11225\ : Odrv4
    port map (
            O => \N__46534\,
            I => \data_out_10__7__N_110\
        );

    \I__11224\ : Odrv4
    port map (
            O => \N__46531\,
            I => \data_out_10__7__N_110\
        );

    \I__11223\ : Odrv4
    port map (
            O => \N__46526\,
            I => \data_out_10__7__N_110\
        );

    \I__11222\ : InMux
    port map (
            O => \N__46519\,
            I => \N__46515\
        );

    \I__11221\ : CascadeMux
    port map (
            O => \N__46518\,
            I => \N__46512\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__46515\,
            I => \N__46509\
        );

    \I__11219\ : InMux
    port map (
            O => \N__46512\,
            I => \N__46506\
        );

    \I__11218\ : Odrv12
    port map (
            O => \N__46509\,
            I => rand_setpoint_21
        );

    \I__11217\ : LocalMux
    port map (
            O => \N__46506\,
            I => rand_setpoint_21
        );

    \I__11216\ : CascadeMux
    port map (
            O => \N__46501\,
            I => \N__46498\
        );

    \I__11215\ : InMux
    port map (
            O => \N__46498\,
            I => \N__46495\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__46495\,
            I => \c0.n17522\
        );

    \I__11213\ : InMux
    port map (
            O => \N__46492\,
            I => \N__46482\
        );

    \I__11212\ : InMux
    port map (
            O => \N__46491\,
            I => \N__46476\
        );

    \I__11211\ : InMux
    port map (
            O => \N__46490\,
            I => \N__46472\
        );

    \I__11210\ : InMux
    port map (
            O => \N__46489\,
            I => \N__46467\
        );

    \I__11209\ : InMux
    port map (
            O => \N__46488\,
            I => \N__46467\
        );

    \I__11208\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46459\
        );

    \I__11207\ : InMux
    port map (
            O => \N__46486\,
            I => \N__46459\
        );

    \I__11206\ : InMux
    port map (
            O => \N__46485\,
            I => \N__46459\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__46482\,
            I => \N__46456\
        );

    \I__11204\ : InMux
    port map (
            O => \N__46481\,
            I => \N__46453\
        );

    \I__11203\ : InMux
    port map (
            O => \N__46480\,
            I => \N__46450\
        );

    \I__11202\ : InMux
    port map (
            O => \N__46479\,
            I => \N__46444\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__46476\,
            I => \N__46441\
        );

    \I__11200\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46438\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__46472\,
            I => \N__46427\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__46467\,
            I => \N__46427\
        );

    \I__11197\ : InMux
    port map (
            O => \N__46466\,
            I => \N__46424\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__46459\,
            I => \N__46408\
        );

    \I__11195\ : Span4Mux_v
    port map (
            O => \N__46456\,
            I => \N__46408\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__46453\,
            I => \N__46408\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46405\
        );

    \I__11192\ : InMux
    port map (
            O => \N__46449\,
            I => \N__46396\
        );

    \I__11191\ : InMux
    port map (
            O => \N__46448\,
            I => \N__46390\
        );

    \I__11190\ : InMux
    port map (
            O => \N__46447\,
            I => \N__46390\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__46444\,
            I => \N__46383\
        );

    \I__11188\ : Span4Mux_v
    port map (
            O => \N__46441\,
            I => \N__46383\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__46438\,
            I => \N__46383\
        );

    \I__11186\ : InMux
    port map (
            O => \N__46437\,
            I => \N__46380\
        );

    \I__11185\ : InMux
    port map (
            O => \N__46436\,
            I => \N__46369\
        );

    \I__11184\ : InMux
    port map (
            O => \N__46435\,
            I => \N__46369\
        );

    \I__11183\ : InMux
    port map (
            O => \N__46434\,
            I => \N__46369\
        );

    \I__11182\ : InMux
    port map (
            O => \N__46433\,
            I => \N__46369\
        );

    \I__11181\ : InMux
    port map (
            O => \N__46432\,
            I => \N__46369\
        );

    \I__11180\ : Span4Mux_v
    port map (
            O => \N__46427\,
            I => \N__46366\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__46424\,
            I => \N__46363\
        );

    \I__11178\ : InMux
    port map (
            O => \N__46423\,
            I => \N__46359\
        );

    \I__11177\ : InMux
    port map (
            O => \N__46422\,
            I => \N__46356\
        );

    \I__11176\ : InMux
    port map (
            O => \N__46421\,
            I => \N__46353\
        );

    \I__11175\ : InMux
    port map (
            O => \N__46420\,
            I => \N__46344\
        );

    \I__11174\ : InMux
    port map (
            O => \N__46419\,
            I => \N__46344\
        );

    \I__11173\ : InMux
    port map (
            O => \N__46418\,
            I => \N__46344\
        );

    \I__11172\ : InMux
    port map (
            O => \N__46417\,
            I => \N__46344\
        );

    \I__11171\ : InMux
    port map (
            O => \N__46416\,
            I => \N__46339\
        );

    \I__11170\ : InMux
    port map (
            O => \N__46415\,
            I => \N__46339\
        );

    \I__11169\ : Span4Mux_v
    port map (
            O => \N__46408\,
            I => \N__46336\
        );

    \I__11168\ : Span4Mux_v
    port map (
            O => \N__46405\,
            I => \N__46333\
        );

    \I__11167\ : InMux
    port map (
            O => \N__46404\,
            I => \N__46322\
        );

    \I__11166\ : InMux
    port map (
            O => \N__46403\,
            I => \N__46322\
        );

    \I__11165\ : InMux
    port map (
            O => \N__46402\,
            I => \N__46322\
        );

    \I__11164\ : InMux
    port map (
            O => \N__46401\,
            I => \N__46322\
        );

    \I__11163\ : InMux
    port map (
            O => \N__46400\,
            I => \N__46322\
        );

    \I__11162\ : CascadeMux
    port map (
            O => \N__46399\,
            I => \N__46318\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__46396\,
            I => \N__46315\
        );

    \I__11160\ : InMux
    port map (
            O => \N__46395\,
            I => \N__46312\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__46390\,
            I => \N__46307\
        );

    \I__11158\ : Span4Mux_h
    port map (
            O => \N__46383\,
            I => \N__46307\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__46380\,
            I => \N__46293\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__46369\,
            I => \N__46293\
        );

    \I__11155\ : Span4Mux_h
    port map (
            O => \N__46366\,
            I => \N__46288\
        );

    \I__11154\ : Span4Mux_v
    port map (
            O => \N__46363\,
            I => \N__46288\
        );

    \I__11153\ : InMux
    port map (
            O => \N__46362\,
            I => \N__46285\
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__46359\,
            I => \N__46268\
        );

    \I__11151\ : LocalMux
    port map (
            O => \N__46356\,
            I => \N__46268\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__46353\,
            I => \N__46268\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__46344\,
            I => \N__46268\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__46339\,
            I => \N__46268\
        );

    \I__11147\ : Sp12to4
    port map (
            O => \N__46336\,
            I => \N__46268\
        );

    \I__11146\ : Sp12to4
    port map (
            O => \N__46333\,
            I => \N__46268\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__46322\,
            I => \N__46268\
        );

    \I__11144\ : InMux
    port map (
            O => \N__46321\,
            I => \N__46263\
        );

    \I__11143\ : InMux
    port map (
            O => \N__46318\,
            I => \N__46263\
        );

    \I__11142\ : Span4Mux_v
    port map (
            O => \N__46315\,
            I => \N__46256\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__46312\,
            I => \N__46256\
        );

    \I__11140\ : Span4Mux_h
    port map (
            O => \N__46307\,
            I => \N__46256\
        );

    \I__11139\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46253\
        );

    \I__11138\ : InMux
    port map (
            O => \N__46305\,
            I => \N__46242\
        );

    \I__11137\ : InMux
    port map (
            O => \N__46304\,
            I => \N__46242\
        );

    \I__11136\ : InMux
    port map (
            O => \N__46303\,
            I => \N__46242\
        );

    \I__11135\ : InMux
    port map (
            O => \N__46302\,
            I => \N__46242\
        );

    \I__11134\ : InMux
    port map (
            O => \N__46301\,
            I => \N__46242\
        );

    \I__11133\ : InMux
    port map (
            O => \N__46300\,
            I => \N__46235\
        );

    \I__11132\ : InMux
    port map (
            O => \N__46299\,
            I => \N__46235\
        );

    \I__11131\ : InMux
    port map (
            O => \N__46298\,
            I => \N__46235\
        );

    \I__11130\ : Span4Mux_h
    port map (
            O => \N__46293\,
            I => \N__46232\
        );

    \I__11129\ : Span4Mux_h
    port map (
            O => \N__46288\,
            I => \N__46227\
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__46285\,
            I => \N__46227\
        );

    \I__11127\ : Span12Mux_h
    port map (
            O => \N__46268\,
            I => \N__46224\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__46263\,
            I => \N__46221\
        );

    \I__11125\ : Span4Mux_h
    port map (
            O => \N__46256\,
            I => \N__46218\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__46253\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__46242\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__46235\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11121\ : Odrv4
    port map (
            O => \N__46232\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11120\ : Odrv4
    port map (
            O => \N__46227\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11119\ : Odrv12
    port map (
            O => \N__46224\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11118\ : Odrv4
    port map (
            O => \N__46221\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11117\ : Odrv4
    port map (
            O => \N__46218\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11116\ : InMux
    port map (
            O => \N__46201\,
            I => \N__46196\
        );

    \I__11115\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46193\
        );

    \I__11114\ : InMux
    port map (
            O => \N__46199\,
            I => \N__46189\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__46196\,
            I => \N__46186\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__46193\,
            I => \N__46183\
        );

    \I__11111\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46180\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__46189\,
            I => \N__46177\
        );

    \I__11109\ : Span4Mux_v
    port map (
            O => \N__46186\,
            I => \N__46174\
        );

    \I__11108\ : Span4Mux_v
    port map (
            O => \N__46183\,
            I => \N__46171\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__46180\,
            I => \N__46166\
        );

    \I__11106\ : Span4Mux_v
    port map (
            O => \N__46177\,
            I => \N__46166\
        );

    \I__11105\ : Span4Mux_v
    port map (
            O => \N__46174\,
            I => \N__46163\
        );

    \I__11104\ : Span4Mux_s1_v
    port map (
            O => \N__46171\,
            I => \N__46160\
        );

    \I__11103\ : Span4Mux_v
    port map (
            O => \N__46166\,
            I => \N__46155\
        );

    \I__11102\ : Span4Mux_h
    port map (
            O => \N__46163\,
            I => \N__46155\
        );

    \I__11101\ : Odrv4
    port map (
            O => \N__46160\,
            I => \c0.data_out_6_5\
        );

    \I__11100\ : Odrv4
    port map (
            O => \N__46155\,
            I => \c0.data_out_6_5\
        );

    \I__11099\ : CascadeMux
    port map (
            O => \N__46150\,
            I => \N__46146\
        );

    \I__11098\ : CascadeMux
    port map (
            O => \N__46149\,
            I => \N__46143\
        );

    \I__11097\ : InMux
    port map (
            O => \N__46146\,
            I => \N__46140\
        );

    \I__11096\ : InMux
    port map (
            O => \N__46143\,
            I => \N__46134\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__46140\,
            I => \N__46125\
        );

    \I__11094\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46122\
        );

    \I__11093\ : CascadeMux
    port map (
            O => \N__46138\,
            I => \N__46119\
        );

    \I__11092\ : CEMux
    port map (
            O => \N__46137\,
            I => \N__46116\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__46134\,
            I => \N__46113\
        );

    \I__11090\ : CascadeMux
    port map (
            O => \N__46133\,
            I => \N__46110\
        );

    \I__11089\ : CascadeMux
    port map (
            O => \N__46132\,
            I => \N__46107\
        );

    \I__11088\ : CEMux
    port map (
            O => \N__46131\,
            I => \N__46103\
        );

    \I__11087\ : CEMux
    port map (
            O => \N__46130\,
            I => \N__46100\
        );

    \I__11086\ : CEMux
    port map (
            O => \N__46129\,
            I => \N__46097\
        );

    \I__11085\ : CEMux
    port map (
            O => \N__46128\,
            I => \N__46094\
        );

    \I__11084\ : Span4Mux_h
    port map (
            O => \N__46125\,
            I => \N__46089\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__46122\,
            I => \N__46089\
        );

    \I__11082\ : InMux
    port map (
            O => \N__46119\,
            I => \N__46086\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__46116\,
            I => \N__46083\
        );

    \I__11080\ : Span4Mux_h
    port map (
            O => \N__46113\,
            I => \N__46080\
        );

    \I__11079\ : InMux
    port map (
            O => \N__46110\,
            I => \N__46077\
        );

    \I__11078\ : InMux
    port map (
            O => \N__46107\,
            I => \N__46074\
        );

    \I__11077\ : CEMux
    port map (
            O => \N__46106\,
            I => \N__46071\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__46103\,
            I => \N__46066\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__46100\,
            I => \N__46066\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__46097\,
            I => \N__46063\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__46094\,
            I => \N__46058\
        );

    \I__11072\ : Span4Mux_h
    port map (
            O => \N__46089\,
            I => \N__46058\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__46086\,
            I => \N__46051\
        );

    \I__11070\ : Span4Mux_s2_v
    port map (
            O => \N__46083\,
            I => \N__46051\
        );

    \I__11069\ : Span4Mux_h
    port map (
            O => \N__46080\,
            I => \N__46051\
        );

    \I__11068\ : LocalMux
    port map (
            O => \N__46077\,
            I => \N__46048\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__46074\,
            I => \N__46041\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__46071\,
            I => \N__46041\
        );

    \I__11065\ : Span4Mux_h
    port map (
            O => \N__46066\,
            I => \N__46041\
        );

    \I__11064\ : Span4Mux_h
    port map (
            O => \N__46063\,
            I => \N__46036\
        );

    \I__11063\ : Span4Mux_h
    port map (
            O => \N__46058\,
            I => \N__46036\
        );

    \I__11062\ : Span4Mux_h
    port map (
            O => \N__46051\,
            I => \N__46033\
        );

    \I__11061\ : Odrv12
    port map (
            O => \N__46048\,
            I => n10055
        );

    \I__11060\ : Odrv4
    port map (
            O => \N__46041\,
            I => n10055
        );

    \I__11059\ : Odrv4
    port map (
            O => \N__46036\,
            I => n10055
        );

    \I__11058\ : Odrv4
    port map (
            O => \N__46033\,
            I => n10055
        );

    \I__11057\ : InMux
    port map (
            O => \N__46024\,
            I => \N__46021\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__46021\,
            I => \N__46018\
        );

    \I__11055\ : Span4Mux_s1_v
    port map (
            O => \N__46018\,
            I => \N__46014\
        );

    \I__11054\ : CascadeMux
    port map (
            O => \N__46017\,
            I => \N__46011\
        );

    \I__11053\ : Span4Mux_h
    port map (
            O => \N__46014\,
            I => \N__46008\
        );

    \I__11052\ : InMux
    port map (
            O => \N__46011\,
            I => \N__46005\
        );

    \I__11051\ : Odrv4
    port map (
            O => \N__46008\,
            I => rand_setpoint_10
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__46005\,
            I => rand_setpoint_10
        );

    \I__11049\ : CascadeMux
    port map (
            O => \N__46000\,
            I => \N__45983\
        );

    \I__11048\ : CascadeMux
    port map (
            O => \N__45999\,
            I => \N__45979\
        );

    \I__11047\ : InMux
    port map (
            O => \N__45998\,
            I => \N__45971\
        );

    \I__11046\ : InMux
    port map (
            O => \N__45997\,
            I => \N__45971\
        );

    \I__11045\ : InMux
    port map (
            O => \N__45996\,
            I => \N__45968\
        );

    \I__11044\ : InMux
    port map (
            O => \N__45995\,
            I => \N__45957\
        );

    \I__11043\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45957\
        );

    \I__11042\ : InMux
    port map (
            O => \N__45993\,
            I => \N__45957\
        );

    \I__11041\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45957\
        );

    \I__11040\ : InMux
    port map (
            O => \N__45991\,
            I => \N__45957\
        );

    \I__11039\ : CascadeMux
    port map (
            O => \N__45990\,
            I => \N__45948\
        );

    \I__11038\ : CascadeMux
    port map (
            O => \N__45989\,
            I => \N__45944\
        );

    \I__11037\ : CascadeMux
    port map (
            O => \N__45988\,
            I => \N__45940\
        );

    \I__11036\ : CascadeMux
    port map (
            O => \N__45987\,
            I => \N__45937\
        );

    \I__11035\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45932\
        );

    \I__11034\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45925\
        );

    \I__11033\ : CascadeMux
    port map (
            O => \N__45982\,
            I => \N__45921\
        );

    \I__11032\ : InMux
    port map (
            O => \N__45979\,
            I => \N__45915\
        );

    \I__11031\ : InMux
    port map (
            O => \N__45978\,
            I => \N__45915\
        );

    \I__11030\ : InMux
    port map (
            O => \N__45977\,
            I => \N__45912\
        );

    \I__11029\ : CascadeMux
    port map (
            O => \N__45976\,
            I => \N__45908\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__45971\,
            I => \N__45898\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__45968\,
            I => \N__45898\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__45957\,
            I => \N__45898\
        );

    \I__11025\ : InMux
    port map (
            O => \N__45956\,
            I => \N__45889\
        );

    \I__11024\ : InMux
    port map (
            O => \N__45955\,
            I => \N__45889\
        );

    \I__11023\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45889\
        );

    \I__11022\ : InMux
    port map (
            O => \N__45953\,
            I => \N__45889\
        );

    \I__11021\ : CascadeMux
    port map (
            O => \N__45952\,
            I => \N__45886\
        );

    \I__11020\ : CascadeMux
    port map (
            O => \N__45951\,
            I => \N__45883\
        );

    \I__11019\ : InMux
    port map (
            O => \N__45948\,
            I => \N__45880\
        );

    \I__11018\ : InMux
    port map (
            O => \N__45947\,
            I => \N__45876\
        );

    \I__11017\ : InMux
    port map (
            O => \N__45944\,
            I => \N__45869\
        );

    \I__11016\ : InMux
    port map (
            O => \N__45943\,
            I => \N__45869\
        );

    \I__11015\ : InMux
    port map (
            O => \N__45940\,
            I => \N__45864\
        );

    \I__11014\ : InMux
    port map (
            O => \N__45937\,
            I => \N__45864\
        );

    \I__11013\ : InMux
    port map (
            O => \N__45936\,
            I => \N__45861\
        );

    \I__11012\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45858\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__45932\,
            I => \N__45855\
        );

    \I__11010\ : InMux
    port map (
            O => \N__45931\,
            I => \N__45852\
        );

    \I__11009\ : InMux
    port map (
            O => \N__45930\,
            I => \N__45849\
        );

    \I__11008\ : CascadeMux
    port map (
            O => \N__45929\,
            I => \N__45845\
        );

    \I__11007\ : CascadeMux
    port map (
            O => \N__45928\,
            I => \N__45841\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__45925\,
            I => \N__45838\
        );

    \I__11005\ : InMux
    port map (
            O => \N__45924\,
            I => \N__45835\
        );

    \I__11004\ : InMux
    port map (
            O => \N__45921\,
            I => \N__45830\
        );

    \I__11003\ : InMux
    port map (
            O => \N__45920\,
            I => \N__45830\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__45915\,
            I => \N__45825\
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__45912\,
            I => \N__45825\
        );

    \I__11000\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45820\
        );

    \I__10999\ : InMux
    port map (
            O => \N__45908\,
            I => \N__45820\
        );

    \I__10998\ : InMux
    port map (
            O => \N__45907\,
            I => \N__45817\
        );

    \I__10997\ : InMux
    port map (
            O => \N__45906\,
            I => \N__45812\
        );

    \I__10996\ : InMux
    port map (
            O => \N__45905\,
            I => \N__45812\
        );

    \I__10995\ : Span4Mux_h
    port map (
            O => \N__45898\,
            I => \N__45807\
        );

    \I__10994\ : LocalMux
    port map (
            O => \N__45889\,
            I => \N__45807\
        );

    \I__10993\ : InMux
    port map (
            O => \N__45886\,
            I => \N__45804\
        );

    \I__10992\ : InMux
    port map (
            O => \N__45883\,
            I => \N__45798\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__45880\,
            I => \N__45795\
        );

    \I__10990\ : InMux
    port map (
            O => \N__45879\,
            I => \N__45792\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__45876\,
            I => \N__45789\
        );

    \I__10988\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45786\
        );

    \I__10987\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45778\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__45869\,
            I => \N__45771\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__45864\,
            I => \N__45771\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__45861\,
            I => \N__45771\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__45858\,
            I => \N__45762\
        );

    \I__10982\ : Span4Mux_h
    port map (
            O => \N__45855\,
            I => \N__45762\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__45852\,
            I => \N__45762\
        );

    \I__10980\ : LocalMux
    port map (
            O => \N__45849\,
            I => \N__45762\
        );

    \I__10979\ : CascadeMux
    port map (
            O => \N__45848\,
            I => \N__45757\
        );

    \I__10978\ : InMux
    port map (
            O => \N__45845\,
            I => \N__45754\
        );

    \I__10977\ : InMux
    port map (
            O => \N__45844\,
            I => \N__45751\
        );

    \I__10976\ : InMux
    port map (
            O => \N__45841\,
            I => \N__45748\
        );

    \I__10975\ : Span4Mux_v
    port map (
            O => \N__45838\,
            I => \N__45745\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__45835\,
            I => \N__45742\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__45830\,
            I => \N__45739\
        );

    \I__10972\ : Span4Mux_v
    port map (
            O => \N__45825\,
            I => \N__45734\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__45820\,
            I => \N__45734\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__45817\,
            I => \N__45725\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__45812\,
            I => \N__45725\
        );

    \I__10968\ : Span4Mux_h
    port map (
            O => \N__45807\,
            I => \N__45725\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__45804\,
            I => \N__45725\
        );

    \I__10966\ : InMux
    port map (
            O => \N__45803\,
            I => \N__45718\
        );

    \I__10965\ : InMux
    port map (
            O => \N__45802\,
            I => \N__45718\
        );

    \I__10964\ : InMux
    port map (
            O => \N__45801\,
            I => \N__45718\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__45798\,
            I => \N__45713\
        );

    \I__10962\ : Span4Mux_v
    port map (
            O => \N__45795\,
            I => \N__45713\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__45792\,
            I => \N__45706\
        );

    \I__10960\ : Span4Mux_s1_v
    port map (
            O => \N__45789\,
            I => \N__45706\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__45786\,
            I => \N__45706\
        );

    \I__10958\ : InMux
    port map (
            O => \N__45785\,
            I => \N__45695\
        );

    \I__10957\ : InMux
    port map (
            O => \N__45784\,
            I => \N__45695\
        );

    \I__10956\ : InMux
    port map (
            O => \N__45783\,
            I => \N__45695\
        );

    \I__10955\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45695\
        );

    \I__10954\ : InMux
    port map (
            O => \N__45781\,
            I => \N__45695\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__45778\,
            I => \N__45688\
        );

    \I__10952\ : Span4Mux_v
    port map (
            O => \N__45771\,
            I => \N__45688\
        );

    \I__10951\ : Span4Mux_v
    port map (
            O => \N__45762\,
            I => \N__45688\
        );

    \I__10950\ : InMux
    port map (
            O => \N__45761\,
            I => \N__45683\
        );

    \I__10949\ : InMux
    port map (
            O => \N__45760\,
            I => \N__45683\
        );

    \I__10948\ : InMux
    port map (
            O => \N__45757\,
            I => \N__45680\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__45754\,
            I => \N__45667\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__45751\,
            I => \N__45667\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__45748\,
            I => \N__45667\
        );

    \I__10944\ : Span4Mux_h
    port map (
            O => \N__45745\,
            I => \N__45667\
        );

    \I__10943\ : Span4Mux_v
    port map (
            O => \N__45742\,
            I => \N__45667\
        );

    \I__10942\ : Span4Mux_v
    port map (
            O => \N__45739\,
            I => \N__45667\
        );

    \I__10941\ : Span4Mux_h
    port map (
            O => \N__45734\,
            I => \N__45662\
        );

    \I__10940\ : Span4Mux_h
    port map (
            O => \N__45725\,
            I => \N__45662\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__45718\,
            I => \N__45651\
        );

    \I__10938\ : Sp12to4
    port map (
            O => \N__45713\,
            I => \N__45651\
        );

    \I__10937\ : Sp12to4
    port map (
            O => \N__45706\,
            I => \N__45651\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__45695\,
            I => \N__45651\
        );

    \I__10935\ : Sp12to4
    port map (
            O => \N__45688\,
            I => \N__45651\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__45683\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__45680\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__10932\ : Odrv4
    port map (
            O => \N__45667\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__10931\ : Odrv4
    port map (
            O => \N__45662\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__10930\ : Odrv12
    port map (
            O => \N__45651\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__10929\ : CascadeMux
    port map (
            O => \N__45640\,
            I => \N__45637\
        );

    \I__10928\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45634\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__45634\,
            I => \N__45631\
        );

    \I__10926\ : Odrv12
    port map (
            O => \N__45631\,
            I => \c0.n17450\
        );

    \I__10925\ : InMux
    port map (
            O => \N__45628\,
            I => \N__45625\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__45625\,
            I => \N__45621\
        );

    \I__10923\ : CascadeMux
    port map (
            O => \N__45624\,
            I => \N__45618\
        );

    \I__10922\ : Span4Mux_v
    port map (
            O => \N__45621\,
            I => \N__45613\
        );

    \I__10921\ : InMux
    port map (
            O => \N__45618\,
            I => \N__45606\
        );

    \I__10920\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45606\
        );

    \I__10919\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45606\
        );

    \I__10918\ : Odrv4
    port map (
            O => \N__45613\,
            I => data_out_frame2_7_5
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__45606\,
            I => data_out_frame2_7_5
        );

    \I__10916\ : CascadeMux
    port map (
            O => \N__45601\,
            I => \N__45598\
        );

    \I__10915\ : InMux
    port map (
            O => \N__45598\,
            I => \N__45593\
        );

    \I__10914\ : InMux
    port map (
            O => \N__45597\,
            I => \N__45590\
        );

    \I__10913\ : InMux
    port map (
            O => \N__45596\,
            I => \N__45587\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__45593\,
            I => \N__45582\
        );

    \I__10911\ : LocalMux
    port map (
            O => \N__45590\,
            I => \N__45582\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__45587\,
            I => \c0.n9678\
        );

    \I__10909\ : Odrv12
    port map (
            O => \N__45582\,
            I => \c0.n9678\
        );

    \I__10908\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45574\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__45574\,
            I => \c0.n18092\
        );

    \I__10906\ : InMux
    port map (
            O => \N__45571\,
            I => \N__45568\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__45568\,
            I => \c0.n22_adj_2352\
        );

    \I__10904\ : InMux
    port map (
            O => \N__45565\,
            I => \N__45562\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__45562\,
            I => \N__45559\
        );

    \I__10902\ : Span4Mux_v
    port map (
            O => \N__45559\,
            I => \N__45556\
        );

    \I__10901\ : Span4Mux_h
    port map (
            O => \N__45556\,
            I => \N__45553\
        );

    \I__10900\ : Odrv4
    port map (
            O => \N__45553\,
            I => \c0.tx2.r_Tx_Data_7\
        );

    \I__10899\ : SRMux
    port map (
            O => \N__45550\,
            I => \N__45541\
        );

    \I__10898\ : CascadeMux
    port map (
            O => \N__45549\,
            I => \N__45538\
        );

    \I__10897\ : InMux
    port map (
            O => \N__45548\,
            I => \N__45533\
        );

    \I__10896\ : InMux
    port map (
            O => \N__45547\,
            I => \N__45526\
        );

    \I__10895\ : InMux
    port map (
            O => \N__45546\,
            I => \N__45526\
        );

    \I__10894\ : InMux
    port map (
            O => \N__45545\,
            I => \N__45526\
        );

    \I__10893\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45523\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__45541\,
            I => \N__45520\
        );

    \I__10891\ : InMux
    port map (
            O => \N__45538\,
            I => \N__45517\
        );

    \I__10890\ : CascadeMux
    port map (
            O => \N__45537\,
            I => \N__45511\
        );

    \I__10889\ : InMux
    port map (
            O => \N__45536\,
            I => \N__45507\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__45533\,
            I => \N__45504\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__45526\,
            I => \N__45499\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__45523\,
            I => \N__45499\
        );

    \I__10885\ : Span4Mux_s2_v
    port map (
            O => \N__45520\,
            I => \N__45496\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__45517\,
            I => \N__45493\
        );

    \I__10883\ : InMux
    port map (
            O => \N__45516\,
            I => \N__45488\
        );

    \I__10882\ : InMux
    port map (
            O => \N__45515\,
            I => \N__45483\
        );

    \I__10881\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45480\
        );

    \I__10880\ : InMux
    port map (
            O => \N__45511\,
            I => \N__45477\
        );

    \I__10879\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45474\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__45507\,
            I => \N__45471\
        );

    \I__10877\ : Span4Mux_s2_v
    port map (
            O => \N__45504\,
            I => \N__45462\
        );

    \I__10876\ : Span4Mux_v
    port map (
            O => \N__45499\,
            I => \N__45462\
        );

    \I__10875\ : Span4Mux_h
    port map (
            O => \N__45496\,
            I => \N__45462\
        );

    \I__10874\ : Span4Mux_s2_v
    port map (
            O => \N__45493\,
            I => \N__45462\
        );

    \I__10873\ : InMux
    port map (
            O => \N__45492\,
            I => \N__45457\
        );

    \I__10872\ : InMux
    port map (
            O => \N__45491\,
            I => \N__45457\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__45488\,
            I => \N__45451\
        );

    \I__10870\ : InMux
    port map (
            O => \N__45487\,
            I => \N__45446\
        );

    \I__10869\ : InMux
    port map (
            O => \N__45486\,
            I => \N__45446\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__45483\,
            I => \N__45443\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__45480\,
            I => \N__45436\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__45477\,
            I => \N__45436\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__45474\,
            I => \N__45436\
        );

    \I__10864\ : Span4Mux_s2_v
    port map (
            O => \N__45471\,
            I => \N__45428\
        );

    \I__10863\ : Span4Mux_h
    port map (
            O => \N__45462\,
            I => \N__45428\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__45457\,
            I => \N__45428\
        );

    \I__10861\ : InMux
    port map (
            O => \N__45456\,
            I => \N__45425\
        );

    \I__10860\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45422\
        );

    \I__10859\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45419\
        );

    \I__10858\ : Span4Mux_v
    port map (
            O => \N__45451\,
            I => \N__45416\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__45446\,
            I => \N__45411\
        );

    \I__10856\ : Span12Mux_s3_v
    port map (
            O => \N__45443\,
            I => \N__45411\
        );

    \I__10855\ : Span4Mux_v
    port map (
            O => \N__45436\,
            I => \N__45408\
        );

    \I__10854\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45405\
        );

    \I__10853\ : Span4Mux_h
    port map (
            O => \N__45428\,
            I => \N__45402\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__45425\,
            I => \N__45399\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__45422\,
            I => n4445
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__45419\,
            I => n4445
        );

    \I__10849\ : Odrv4
    port map (
            O => \N__45416\,
            I => n4445
        );

    \I__10848\ : Odrv12
    port map (
            O => \N__45411\,
            I => n4445
        );

    \I__10847\ : Odrv4
    port map (
            O => \N__45408\,
            I => n4445
        );

    \I__10846\ : LocalMux
    port map (
            O => \N__45405\,
            I => n4445
        );

    \I__10845\ : Odrv4
    port map (
            O => \N__45402\,
            I => n4445
        );

    \I__10844\ : Odrv4
    port map (
            O => \N__45399\,
            I => n4445
        );

    \I__10843\ : CascadeMux
    port map (
            O => \N__45382\,
            I => \N__45379\
        );

    \I__10842\ : InMux
    port map (
            O => \N__45379\,
            I => \N__45375\
        );

    \I__10841\ : InMux
    port map (
            O => \N__45378\,
            I => \N__45372\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__45375\,
            I => data_out_0_0
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__45372\,
            I => data_out_0_0
        );

    \I__10838\ : InMux
    port map (
            O => \N__45367\,
            I => \N__45364\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__45364\,
            I => \N__45358\
        );

    \I__10836\ : InMux
    port map (
            O => \N__45363\,
            I => \N__45355\
        );

    \I__10835\ : InMux
    port map (
            O => \N__45362\,
            I => \N__45352\
        );

    \I__10834\ : CascadeMux
    port map (
            O => \N__45361\,
            I => \N__45349\
        );

    \I__10833\ : Span4Mux_h
    port map (
            O => \N__45358\,
            I => \N__45343\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__45355\,
            I => \N__45343\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__45352\,
            I => \N__45340\
        );

    \I__10830\ : InMux
    port map (
            O => \N__45349\,
            I => \N__45337\
        );

    \I__10829\ : InMux
    port map (
            O => \N__45348\,
            I => \N__45333\
        );

    \I__10828\ : Span4Mux_h
    port map (
            O => \N__45343\,
            I => \N__45330\
        );

    \I__10827\ : Span4Mux_h
    port map (
            O => \N__45340\,
            I => \N__45327\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__45337\,
            I => \N__45324\
        );

    \I__10825\ : InMux
    port map (
            O => \N__45336\,
            I => \N__45321\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__45333\,
            I => \N__45318\
        );

    \I__10823\ : Span4Mux_v
    port map (
            O => \N__45330\,
            I => \N__45315\
        );

    \I__10822\ : Span4Mux_v
    port map (
            O => \N__45327\,
            I => \N__45310\
        );

    \I__10821\ : Span4Mux_v
    port map (
            O => \N__45324\,
            I => \N__45310\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__45321\,
            I => data_out_frame2_12_3
        );

    \I__10819\ : Odrv4
    port map (
            O => \N__45318\,
            I => data_out_frame2_12_3
        );

    \I__10818\ : Odrv4
    port map (
            O => \N__45315\,
            I => data_out_frame2_12_3
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__45310\,
            I => data_out_frame2_12_3
        );

    \I__10816\ : InMux
    port map (
            O => \N__45301\,
            I => \N__45297\
        );

    \I__10815\ : InMux
    port map (
            O => \N__45300\,
            I => \N__45294\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__45297\,
            I => \N__45289\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__45294\,
            I => \N__45286\
        );

    \I__10812\ : InMux
    port map (
            O => \N__45293\,
            I => \N__45283\
        );

    \I__10811\ : InMux
    port map (
            O => \N__45292\,
            I => \N__45280\
        );

    \I__10810\ : Span4Mux_v
    port map (
            O => \N__45289\,
            I => \N__45272\
        );

    \I__10809\ : Span4Mux_v
    port map (
            O => \N__45286\,
            I => \N__45272\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__45283\,
            I => \N__45272\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__45280\,
            I => \N__45269\
        );

    \I__10806\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45266\
        );

    \I__10805\ : Span4Mux_h
    port map (
            O => \N__45272\,
            I => \N__45261\
        );

    \I__10804\ : Span4Mux_s2_v
    port map (
            O => \N__45269\,
            I => \N__45261\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__45266\,
            I => rand_data_29
        );

    \I__10802\ : Odrv4
    port map (
            O => \N__45261\,
            I => rand_data_29
        );

    \I__10801\ : CascadeMux
    port map (
            O => \N__45256\,
            I => \N__45253\
        );

    \I__10800\ : InMux
    port map (
            O => \N__45253\,
            I => \N__45249\
        );

    \I__10799\ : InMux
    port map (
            O => \N__45252\,
            I => \N__45245\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__45249\,
            I => \N__45242\
        );

    \I__10797\ : InMux
    port map (
            O => \N__45248\,
            I => \N__45239\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__45245\,
            I => \N__45235\
        );

    \I__10795\ : Span4Mux_v
    port map (
            O => \N__45242\,
            I => \N__45230\
        );

    \I__10794\ : LocalMux
    port map (
            O => \N__45239\,
            I => \N__45230\
        );

    \I__10793\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45227\
        );

    \I__10792\ : Span4Mux_h
    port map (
            O => \N__45235\,
            I => \N__45224\
        );

    \I__10791\ : Span4Mux_h
    port map (
            O => \N__45230\,
            I => \N__45221\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__45227\,
            I => data_out_frame2_13_5
        );

    \I__10789\ : Odrv4
    port map (
            O => \N__45224\,
            I => data_out_frame2_13_5
        );

    \I__10788\ : Odrv4
    port map (
            O => \N__45221\,
            I => data_out_frame2_13_5
        );

    \I__10787\ : CascadeMux
    port map (
            O => \N__45214\,
            I => \N__45210\
        );

    \I__10786\ : InMux
    port map (
            O => \N__45213\,
            I => \N__45207\
        );

    \I__10785\ : InMux
    port map (
            O => \N__45210\,
            I => \N__45202\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__45207\,
            I => \N__45198\
        );

    \I__10783\ : InMux
    port map (
            O => \N__45206\,
            I => \N__45195\
        );

    \I__10782\ : InMux
    port map (
            O => \N__45205\,
            I => \N__45192\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__45202\,
            I => \N__45188\
        );

    \I__10780\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45185\
        );

    \I__10779\ : Span4Mux_v
    port map (
            O => \N__45198\,
            I => \N__45182\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__45195\,
            I => \N__45177\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__45192\,
            I => \N__45177\
        );

    \I__10776\ : InMux
    port map (
            O => \N__45191\,
            I => \N__45174\
        );

    \I__10775\ : Span4Mux_s3_v
    port map (
            O => \N__45188\,
            I => \N__45169\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__45185\,
            I => \N__45169\
        );

    \I__10773\ : Span4Mux_h
    port map (
            O => \N__45182\,
            I => \N__45166\
        );

    \I__10772\ : Span4Mux_h
    port map (
            O => \N__45177\,
            I => \N__45161\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__45174\,
            I => \N__45161\
        );

    \I__10770\ : Span4Mux_h
    port map (
            O => \N__45169\,
            I => \N__45158\
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__45166\,
            I => \c0.data_out_5_1\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__45161\,
            I => \c0.data_out_5_1\
        );

    \I__10767\ : Odrv4
    port map (
            O => \N__45158\,
            I => \c0.data_out_5_1\
        );

    \I__10766\ : InMux
    port map (
            O => \N__45151\,
            I => \N__45148\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__45148\,
            I => \N__45145\
        );

    \I__10764\ : Span4Mux_h
    port map (
            O => \N__45145\,
            I => \N__45141\
        );

    \I__10763\ : InMux
    port map (
            O => \N__45144\,
            I => \N__45138\
        );

    \I__10762\ : Odrv4
    port map (
            O => \N__45141\,
            I => \c0.n17043\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__45138\,
            I => \c0.n17043\
        );

    \I__10760\ : CascadeMux
    port map (
            O => \N__45133\,
            I => \N__45130\
        );

    \I__10759\ : InMux
    port map (
            O => \N__45130\,
            I => \N__45127\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__45127\,
            I => \N__45124\
        );

    \I__10757\ : Span4Mux_v
    port map (
            O => \N__45124\,
            I => \N__45121\
        );

    \I__10756\ : Odrv4
    port map (
            O => \N__45121\,
            I => \c0.n16949\
        );

    \I__10755\ : InMux
    port map (
            O => \N__45118\,
            I => \N__45115\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__45115\,
            I => \N__45111\
        );

    \I__10753\ : InMux
    port map (
            O => \N__45114\,
            I => \N__45108\
        );

    \I__10752\ : Span4Mux_v
    port map (
            O => \N__45111\,
            I => \N__45103\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__45108\,
            I => \N__45100\
        );

    \I__10750\ : InMux
    port map (
            O => \N__45107\,
            I => \N__45094\
        );

    \I__10749\ : InMux
    port map (
            O => \N__45106\,
            I => \N__45094\
        );

    \I__10748\ : Span4Mux_h
    port map (
            O => \N__45103\,
            I => \N__45089\
        );

    \I__10747\ : Span4Mux_h
    port map (
            O => \N__45100\,
            I => \N__45089\
        );

    \I__10746\ : InMux
    port map (
            O => \N__45099\,
            I => \N__45086\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__45094\,
            I => data_out_8_7
        );

    \I__10744\ : Odrv4
    port map (
            O => \N__45089\,
            I => data_out_8_7
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__45086\,
            I => data_out_8_7
        );

    \I__10742\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45076\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__45076\,
            I => \N__45071\
        );

    \I__10740\ : InMux
    port map (
            O => \N__45075\,
            I => \N__45064\
        );

    \I__10739\ : InMux
    port map (
            O => \N__45074\,
            I => \N__45064\
        );

    \I__10738\ : Span4Mux_h
    port map (
            O => \N__45071\,
            I => \N__45061\
        );

    \I__10737\ : InMux
    port map (
            O => \N__45070\,
            I => \N__45058\
        );

    \I__10736\ : InMux
    port map (
            O => \N__45069\,
            I => \N__45054\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__45064\,
            I => \N__45051\
        );

    \I__10734\ : Span4Mux_h
    port map (
            O => \N__45061\,
            I => \N__45046\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__45058\,
            I => \N__45046\
        );

    \I__10732\ : InMux
    port map (
            O => \N__45057\,
            I => \N__45043\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__45054\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__10730\ : Odrv4
    port map (
            O => \N__45051\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__10729\ : Odrv4
    port map (
            O => \N__45046\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__45043\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__10727\ : InMux
    port map (
            O => \N__45034\,
            I => \N__45031\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__45031\,
            I => \N__45028\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__45028\,
            I => \N__45025\
        );

    \I__10724\ : Odrv4
    port map (
            O => \N__45025\,
            I => \c0.n10_adj_2276\
        );

    \I__10723\ : InMux
    port map (
            O => \N__45022\,
            I => \N__45017\
        );

    \I__10722\ : InMux
    port map (
            O => \N__45021\,
            I => \N__45012\
        );

    \I__10721\ : InMux
    port map (
            O => \N__45020\,
            I => \N__45012\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__45017\,
            I => \N__45009\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__45012\,
            I => \c0.data_out_9_3\
        );

    \I__10718\ : Odrv4
    port map (
            O => \N__45009\,
            I => \c0.data_out_9_3\
        );

    \I__10717\ : InMux
    port map (
            O => \N__45004\,
            I => \N__45001\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__45001\,
            I => \N__44997\
        );

    \I__10715\ : InMux
    port map (
            O => \N__45000\,
            I => \N__44994\
        );

    \I__10714\ : Span4Mux_v
    port map (
            O => \N__44997\,
            I => \N__44991\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__44994\,
            I => \N__44988\
        );

    \I__10712\ : Span4Mux_h
    port map (
            O => \N__44991\,
            I => \N__44985\
        );

    \I__10711\ : Span4Mux_v
    port map (
            O => \N__44988\,
            I => \N__44982\
        );

    \I__10710\ : Odrv4
    port map (
            O => \N__44985\,
            I => \c0.n16981\
        );

    \I__10709\ : Odrv4
    port map (
            O => \N__44982\,
            I => \c0.n16981\
        );

    \I__10708\ : InMux
    port map (
            O => \N__44977\,
            I => \N__44974\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__44974\,
            I => \N__44970\
        );

    \I__10706\ : CascadeMux
    port map (
            O => \N__44973\,
            I => \N__44967\
        );

    \I__10705\ : Span4Mux_v
    port map (
            O => \N__44970\,
            I => \N__44964\
        );

    \I__10704\ : InMux
    port map (
            O => \N__44967\,
            I => \N__44961\
        );

    \I__10703\ : Span4Mux_h
    port map (
            O => \N__44964\,
            I => \N__44958\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__44961\,
            I => \N__44955\
        );

    \I__10701\ : Odrv4
    port map (
            O => \N__44958\,
            I => \c0.n16969\
        );

    \I__10700\ : Odrv4
    port map (
            O => \N__44955\,
            I => \c0.n16969\
        );

    \I__10699\ : InMux
    port map (
            O => \N__44950\,
            I => \N__44947\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__44947\,
            I => \N__44940\
        );

    \I__10697\ : InMux
    port map (
            O => \N__44946\,
            I => \N__44937\
        );

    \I__10696\ : InMux
    port map (
            O => \N__44945\,
            I => \N__44934\
        );

    \I__10695\ : InMux
    port map (
            O => \N__44944\,
            I => \N__44931\
        );

    \I__10694\ : CascadeMux
    port map (
            O => \N__44943\,
            I => \N__44928\
        );

    \I__10693\ : Span4Mux_v
    port map (
            O => \N__44940\,
            I => \N__44925\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__44937\,
            I => \N__44922\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__44934\,
            I => \N__44919\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__44931\,
            I => \N__44915\
        );

    \I__10689\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44912\
        );

    \I__10688\ : Span4Mux_h
    port map (
            O => \N__44925\,
            I => \N__44907\
        );

    \I__10687\ : Span4Mux_h
    port map (
            O => \N__44922\,
            I => \N__44907\
        );

    \I__10686\ : Span4Mux_h
    port map (
            O => \N__44919\,
            I => \N__44904\
        );

    \I__10685\ : InMux
    port map (
            O => \N__44918\,
            I => \N__44901\
        );

    \I__10684\ : Span12Mux_h
    port map (
            O => \N__44915\,
            I => \N__44896\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__44912\,
            I => \N__44896\
        );

    \I__10682\ : Odrv4
    port map (
            O => \N__44907\,
            I => rand_data_15
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__44904\,
            I => rand_data_15
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__44901\,
            I => rand_data_15
        );

    \I__10679\ : Odrv12
    port map (
            O => \N__44896\,
            I => rand_data_15
        );

    \I__10678\ : InMux
    port map (
            O => \N__44887\,
            I => \N__44883\
        );

    \I__10677\ : InMux
    port map (
            O => \N__44886\,
            I => \N__44879\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__44883\,
            I => \N__44874\
        );

    \I__10675\ : InMux
    port map (
            O => \N__44882\,
            I => \N__44871\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__44879\,
            I => \N__44868\
        );

    \I__10673\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44863\
        );

    \I__10672\ : InMux
    port map (
            O => \N__44877\,
            I => \N__44863\
        );

    \I__10671\ : Odrv12
    port map (
            O => \N__44874\,
            I => data_out_frame2_9_7
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__44871\,
            I => data_out_frame2_9_7
        );

    \I__10669\ : Odrv4
    port map (
            O => \N__44868\,
            I => data_out_frame2_9_7
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__44863\,
            I => data_out_frame2_9_7
        );

    \I__10667\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44849\
        );

    \I__10666\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44846\
        );

    \I__10665\ : CascadeMux
    port map (
            O => \N__44852\,
            I => \N__44843\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__44849\,
            I => \N__44838\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__44846\,
            I => \N__44835\
        );

    \I__10662\ : InMux
    port map (
            O => \N__44843\,
            I => \N__44832\
        );

    \I__10661\ : InMux
    port map (
            O => \N__44842\,
            I => \N__44829\
        );

    \I__10660\ : InMux
    port map (
            O => \N__44841\,
            I => \N__44826\
        );

    \I__10659\ : Span4Mux_h
    port map (
            O => \N__44838\,
            I => \N__44823\
        );

    \I__10658\ : Span4Mux_h
    port map (
            O => \N__44835\,
            I => \N__44820\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__44832\,
            I => \N__44817\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__44829\,
            I => data_out_frame2_9_5
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__44826\,
            I => data_out_frame2_9_5
        );

    \I__10654\ : Odrv4
    port map (
            O => \N__44823\,
            I => data_out_frame2_9_5
        );

    \I__10653\ : Odrv4
    port map (
            O => \N__44820\,
            I => data_out_frame2_9_5
        );

    \I__10652\ : Odrv4
    port map (
            O => \N__44817\,
            I => data_out_frame2_9_5
        );

    \I__10651\ : CascadeMux
    port map (
            O => \N__44806\,
            I => \N__44803\
        );

    \I__10650\ : InMux
    port map (
            O => \N__44803\,
            I => \N__44800\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__44800\,
            I => \N__44797\
        );

    \I__10648\ : Span4Mux_h
    port map (
            O => \N__44797\,
            I => \N__44794\
        );

    \I__10647\ : Span4Mux_h
    port map (
            O => \N__44794\,
            I => \N__44791\
        );

    \I__10646\ : Odrv4
    port map (
            O => \N__44791\,
            I => \c0.n16926\
        );

    \I__10645\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44785\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__44785\,
            I => \N__44779\
        );

    \I__10643\ : InMux
    port map (
            O => \N__44784\,
            I => \N__44776\
        );

    \I__10642\ : InMux
    port map (
            O => \N__44783\,
            I => \N__44773\
        );

    \I__10641\ : InMux
    port map (
            O => \N__44782\,
            I => \N__44770\
        );

    \I__10640\ : Span4Mux_h
    port map (
            O => \N__44779\,
            I => \N__44765\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__44776\,
            I => \N__44765\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__44773\,
            I => \N__44762\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__44770\,
            I => \N__44758\
        );

    \I__10636\ : Span4Mux_h
    port map (
            O => \N__44765\,
            I => \N__44755\
        );

    \I__10635\ : Span4Mux_h
    port map (
            O => \N__44762\,
            I => \N__44752\
        );

    \I__10634\ : InMux
    port map (
            O => \N__44761\,
            I => \N__44749\
        );

    \I__10633\ : Span4Mux_s2_v
    port map (
            O => \N__44758\,
            I => \N__44746\
        );

    \I__10632\ : Odrv4
    port map (
            O => \N__44755\,
            I => rand_data_24
        );

    \I__10631\ : Odrv4
    port map (
            O => \N__44752\,
            I => rand_data_24
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__44749\,
            I => rand_data_24
        );

    \I__10629\ : Odrv4
    port map (
            O => \N__44746\,
            I => rand_data_24
        );

    \I__10628\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44731\
        );

    \I__10627\ : CascadeMux
    port map (
            O => \N__44736\,
            I => \N__44728\
        );

    \I__10626\ : InMux
    port map (
            O => \N__44735\,
            I => \N__44723\
        );

    \I__10625\ : InMux
    port map (
            O => \N__44734\,
            I => \N__44723\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__44731\,
            I => \N__44720\
        );

    \I__10623\ : InMux
    port map (
            O => \N__44728\,
            I => \N__44717\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__44723\,
            I => \N__44713\
        );

    \I__10621\ : Span4Mux_v
    port map (
            O => \N__44720\,
            I => \N__44708\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__44717\,
            I => \N__44708\
        );

    \I__10619\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44705\
        );

    \I__10618\ : Span4Mux_v
    port map (
            O => \N__44713\,
            I => \N__44700\
        );

    \I__10617\ : Span4Mux_h
    port map (
            O => \N__44708\,
            I => \N__44700\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__44705\,
            I => data_out_frame2_5_0
        );

    \I__10615\ : Odrv4
    port map (
            O => \N__44700\,
            I => data_out_frame2_5_0
        );

    \I__10614\ : InMux
    port map (
            O => \N__44695\,
            I => \N__44691\
        );

    \I__10613\ : CascadeMux
    port map (
            O => \N__44694\,
            I => \N__44688\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__44691\,
            I => \N__44683\
        );

    \I__10611\ : InMux
    port map (
            O => \N__44688\,
            I => \N__44680\
        );

    \I__10610\ : InMux
    port map (
            O => \N__44687\,
            I => \N__44677\
        );

    \I__10609\ : InMux
    port map (
            O => \N__44686\,
            I => \N__44674\
        );

    \I__10608\ : Span4Mux_h
    port map (
            O => \N__44683\,
            I => \N__44667\
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__44680\,
            I => \N__44667\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__44677\,
            I => \N__44667\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__44674\,
            I => \N__44663\
        );

    \I__10604\ : Span4Mux_h
    port map (
            O => \N__44667\,
            I => \N__44660\
        );

    \I__10603\ : InMux
    port map (
            O => \N__44666\,
            I => \N__44657\
        );

    \I__10602\ : Span4Mux_s2_v
    port map (
            O => \N__44663\,
            I => \N__44654\
        );

    \I__10601\ : Odrv4
    port map (
            O => \N__44660\,
            I => rand_data_25
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__44657\,
            I => rand_data_25
        );

    \I__10599\ : Odrv4
    port map (
            O => \N__44654\,
            I => rand_data_25
        );

    \I__10598\ : InMux
    port map (
            O => \N__44647\,
            I => \N__44643\
        );

    \I__10597\ : InMux
    port map (
            O => \N__44646\,
            I => \N__44639\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__44643\,
            I => \N__44636\
        );

    \I__10595\ : CascadeMux
    port map (
            O => \N__44642\,
            I => \N__44633\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__44639\,
            I => \N__44629\
        );

    \I__10593\ : Span4Mux_v
    port map (
            O => \N__44636\,
            I => \N__44626\
        );

    \I__10592\ : InMux
    port map (
            O => \N__44633\,
            I => \N__44621\
        );

    \I__10591\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44621\
        );

    \I__10590\ : Odrv12
    port map (
            O => \N__44629\,
            I => data_out_frame2_6_5
        );

    \I__10589\ : Odrv4
    port map (
            O => \N__44626\,
            I => data_out_frame2_6_5
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__44621\,
            I => data_out_frame2_6_5
        );

    \I__10587\ : CascadeMux
    port map (
            O => \N__44614\,
            I => \N__44611\
        );

    \I__10586\ : InMux
    port map (
            O => \N__44611\,
            I => \N__44607\
        );

    \I__10585\ : InMux
    port map (
            O => \N__44610\,
            I => \N__44602\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__44607\,
            I => \N__44599\
        );

    \I__10583\ : InMux
    port map (
            O => \N__44606\,
            I => \N__44596\
        );

    \I__10582\ : InMux
    port map (
            O => \N__44605\,
            I => \N__44593\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__44602\,
            I => data_out_frame2_5_5
        );

    \I__10580\ : Odrv4
    port map (
            O => \N__44599\,
            I => data_out_frame2_5_5
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__44596\,
            I => data_out_frame2_5_5
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__44593\,
            I => data_out_frame2_5_5
        );

    \I__10577\ : CascadeMux
    port map (
            O => \N__44584\,
            I => \c0.n5_adj_2349_cascade_\
        );

    \I__10576\ : InMux
    port map (
            O => \N__44581\,
            I => \N__44578\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__44578\,
            I => \N__44575\
        );

    \I__10574\ : Span4Mux_h
    port map (
            O => \N__44575\,
            I => \N__44572\
        );

    \I__10573\ : Odrv4
    port map (
            O => \N__44572\,
            I => \c0.n6_adj_2280\
        );

    \I__10572\ : InMux
    port map (
            O => \N__44569\,
            I => \N__44563\
        );

    \I__10571\ : InMux
    port map (
            O => \N__44568\,
            I => \N__44558\
        );

    \I__10570\ : InMux
    port map (
            O => \N__44567\,
            I => \N__44558\
        );

    \I__10569\ : CascadeMux
    port map (
            O => \N__44566\,
            I => \N__44554\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__44563\,
            I => \N__44551\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__44558\,
            I => \N__44548\
        );

    \I__10566\ : InMux
    port map (
            O => \N__44557\,
            I => \N__44544\
        );

    \I__10565\ : InMux
    port map (
            O => \N__44554\,
            I => \N__44541\
        );

    \I__10564\ : Span4Mux_h
    port map (
            O => \N__44551\,
            I => \N__44538\
        );

    \I__10563\ : Span4Mux_v
    port map (
            O => \N__44548\,
            I => \N__44535\
        );

    \I__10562\ : InMux
    port map (
            O => \N__44547\,
            I => \N__44532\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__44544\,
            I => \N__44527\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__44541\,
            I => \N__44527\
        );

    \I__10559\ : Odrv4
    port map (
            O => \N__44538\,
            I => rand_data_13
        );

    \I__10558\ : Odrv4
    port map (
            O => \N__44535\,
            I => rand_data_13
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__44532\,
            I => rand_data_13
        );

    \I__10556\ : Odrv12
    port map (
            O => \N__44527\,
            I => rand_data_13
        );

    \I__10555\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44515\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__44515\,
            I => \N__44512\
        );

    \I__10553\ : Odrv12
    port map (
            O => \N__44512\,
            I => \c0.n6_adj_2278\
        );

    \I__10552\ : InMux
    port map (
            O => \N__44509\,
            I => \N__44506\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__44506\,
            I => \N__44503\
        );

    \I__10550\ : Odrv4
    port map (
            O => \N__44503\,
            I => \c0.n18089\
        );

    \I__10549\ : CascadeMux
    port map (
            O => \N__44500\,
            I => \N__44497\
        );

    \I__10548\ : InMux
    port map (
            O => \N__44497\,
            I => \N__44494\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__44494\,
            I => \N__44491\
        );

    \I__10546\ : Odrv12
    port map (
            O => \N__44491\,
            I => \c0.n17561\
        );

    \I__10545\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44484\
        );

    \I__10544\ : InMux
    port map (
            O => \N__44487\,
            I => \N__44481\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__44484\,
            I => \N__44477\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__44481\,
            I => \N__44474\
        );

    \I__10541\ : InMux
    port map (
            O => \N__44480\,
            I => \N__44471\
        );

    \I__10540\ : Span4Mux_v
    port map (
            O => \N__44477\,
            I => \N__44463\
        );

    \I__10539\ : Span4Mux_v
    port map (
            O => \N__44474\,
            I => \N__44463\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__44471\,
            I => \N__44463\
        );

    \I__10537\ : InMux
    port map (
            O => \N__44470\,
            I => \N__44459\
        );

    \I__10536\ : Span4Mux_h
    port map (
            O => \N__44463\,
            I => \N__44456\
        );

    \I__10535\ : InMux
    port map (
            O => \N__44462\,
            I => \N__44453\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__44459\,
            I => \N__44450\
        );

    \I__10533\ : Odrv4
    port map (
            O => \N__44456\,
            I => rand_data_18
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__44453\,
            I => rand_data_18
        );

    \I__10531\ : Odrv12
    port map (
            O => \N__44450\,
            I => rand_data_18
        );

    \I__10530\ : CascadeMux
    port map (
            O => \N__44443\,
            I => \N__44438\
        );

    \I__10529\ : InMux
    port map (
            O => \N__44442\,
            I => \N__44435\
        );

    \I__10528\ : InMux
    port map (
            O => \N__44441\,
            I => \N__44431\
        );

    \I__10527\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44428\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__44435\,
            I => \N__44425\
        );

    \I__10525\ : InMux
    port map (
            O => \N__44434\,
            I => \N__44422\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__44431\,
            I => \N__44418\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__44428\,
            I => \N__44411\
        );

    \I__10522\ : Span4Mux_v
    port map (
            O => \N__44425\,
            I => \N__44411\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__44422\,
            I => \N__44411\
        );

    \I__10520\ : InMux
    port map (
            O => \N__44421\,
            I => \N__44408\
        );

    \I__10519\ : Span4Mux_v
    port map (
            O => \N__44418\,
            I => \N__44405\
        );

    \I__10518\ : Span4Mux_h
    port map (
            O => \N__44411\,
            I => \N__44402\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__44408\,
            I => data_out_frame2_6_2
        );

    \I__10516\ : Odrv4
    port map (
            O => \N__44405\,
            I => data_out_frame2_6_2
        );

    \I__10515\ : Odrv4
    port map (
            O => \N__44402\,
            I => data_out_frame2_6_2
        );

    \I__10514\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44390\
        );

    \I__10513\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44385\
        );

    \I__10512\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44385\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__44390\,
            I => \N__44382\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__44385\,
            I => \N__44379\
        );

    \I__10509\ : Span4Mux_h
    port map (
            O => \N__44382\,
            I => \N__44375\
        );

    \I__10508\ : Span4Mux_h
    port map (
            O => \N__44379\,
            I => \N__44372\
        );

    \I__10507\ : InMux
    port map (
            O => \N__44378\,
            I => \N__44369\
        );

    \I__10506\ : Span4Mux_h
    port map (
            O => \N__44375\,
            I => \N__44366\
        );

    \I__10505\ : Span4Mux_h
    port map (
            O => \N__44372\,
            I => \N__44363\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__44369\,
            I => data_out_frame2_15_6
        );

    \I__10503\ : Odrv4
    port map (
            O => \N__44366\,
            I => data_out_frame2_15_6
        );

    \I__10502\ : Odrv4
    port map (
            O => \N__44363\,
            I => data_out_frame2_15_6
        );

    \I__10501\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44351\
        );

    \I__10500\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44348\
        );

    \I__10499\ : InMux
    port map (
            O => \N__44354\,
            I => \N__44342\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__44351\,
            I => \N__44339\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__44348\,
            I => \N__44336\
        );

    \I__10496\ : InMux
    port map (
            O => \N__44347\,
            I => \N__44333\
        );

    \I__10495\ : InMux
    port map (
            O => \N__44346\,
            I => \N__44328\
        );

    \I__10494\ : InMux
    port map (
            O => \N__44345\,
            I => \N__44328\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__44342\,
            I => \N__44323\
        );

    \I__10492\ : Span4Mux_v
    port map (
            O => \N__44339\,
            I => \N__44323\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__44336\,
            I => \N__44320\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__44333\,
            I => \N__44315\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__44328\,
            I => \N__44315\
        );

    \I__10488\ : Odrv4
    port map (
            O => \N__44323\,
            I => data_out_frame2_7_6
        );

    \I__10487\ : Odrv4
    port map (
            O => \N__44320\,
            I => data_out_frame2_7_6
        );

    \I__10486\ : Odrv12
    port map (
            O => \N__44315\,
            I => data_out_frame2_7_6
        );

    \I__10485\ : InMux
    port map (
            O => \N__44308\,
            I => \N__44304\
        );

    \I__10484\ : InMux
    port map (
            O => \N__44307\,
            I => \N__44301\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__44304\,
            I => \N__44298\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__44301\,
            I => \N__44295\
        );

    \I__10481\ : Sp12to4
    port map (
            O => \N__44298\,
            I => \N__44292\
        );

    \I__10480\ : Span4Mux_h
    port map (
            O => \N__44295\,
            I => \N__44289\
        );

    \I__10479\ : Odrv12
    port map (
            O => \N__44292\,
            I => \c0.n17127\
        );

    \I__10478\ : Odrv4
    port map (
            O => \N__44289\,
            I => \c0.n17127\
        );

    \I__10477\ : InMux
    port map (
            O => \N__44284\,
            I => \N__44279\
        );

    \I__10476\ : CascadeMux
    port map (
            O => \N__44283\,
            I => \N__44276\
        );

    \I__10475\ : InMux
    port map (
            O => \N__44282\,
            I => \N__44273\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__44279\,
            I => \N__44269\
        );

    \I__10473\ : InMux
    port map (
            O => \N__44276\,
            I => \N__44266\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__44273\,
            I => \N__44263\
        );

    \I__10471\ : InMux
    port map (
            O => \N__44272\,
            I => \N__44260\
        );

    \I__10470\ : Span4Mux_h
    port map (
            O => \N__44269\,
            I => \N__44257\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__44266\,
            I => \N__44254\
        );

    \I__10468\ : Span4Mux_h
    port map (
            O => \N__44263\,
            I => \N__44251\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__44260\,
            I => data_out_frame2_8_7
        );

    \I__10466\ : Odrv4
    port map (
            O => \N__44257\,
            I => data_out_frame2_8_7
        );

    \I__10465\ : Odrv4
    port map (
            O => \N__44254\,
            I => data_out_frame2_8_7
        );

    \I__10464\ : Odrv4
    port map (
            O => \N__44251\,
            I => data_out_frame2_8_7
        );

    \I__10463\ : InMux
    port map (
            O => \N__44242\,
            I => \N__44238\
        );

    \I__10462\ : InMux
    port map (
            O => \N__44241\,
            I => \N__44235\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__44238\,
            I => \N__44232\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__44235\,
            I => \N__44225\
        );

    \I__10459\ : Span4Mux_v
    port map (
            O => \N__44232\,
            I => \N__44225\
        );

    \I__10458\ : InMux
    port map (
            O => \N__44231\,
            I => \N__44222\
        );

    \I__10457\ : InMux
    port map (
            O => \N__44230\,
            I => \N__44218\
        );

    \I__10456\ : Span4Mux_v
    port map (
            O => \N__44225\,
            I => \N__44215\
        );

    \I__10455\ : LocalMux
    port map (
            O => \N__44222\,
            I => \N__44212\
        );

    \I__10454\ : InMux
    port map (
            O => \N__44221\,
            I => \N__44209\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__44218\,
            I => data_out_frame2_11_6
        );

    \I__10452\ : Odrv4
    port map (
            O => \N__44215\,
            I => data_out_frame2_11_6
        );

    \I__10451\ : Odrv12
    port map (
            O => \N__44212\,
            I => data_out_frame2_11_6
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__44209\,
            I => data_out_frame2_11_6
        );

    \I__10449\ : InMux
    port map (
            O => \N__44200\,
            I => \N__44197\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__44197\,
            I => \N__44192\
        );

    \I__10447\ : InMux
    port map (
            O => \N__44196\,
            I => \N__44189\
        );

    \I__10446\ : InMux
    port map (
            O => \N__44195\,
            I => \N__44186\
        );

    \I__10445\ : Span4Mux_v
    port map (
            O => \N__44192\,
            I => \N__44183\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__44189\,
            I => \N__44180\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__44186\,
            I => data_out_frame2_14_7
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__44183\,
            I => data_out_frame2_14_7
        );

    \I__10441\ : Odrv4
    port map (
            O => \N__44180\,
            I => data_out_frame2_14_7
        );

    \I__10440\ : CascadeMux
    port map (
            O => \N__44173\,
            I => \N__44169\
        );

    \I__10439\ : InMux
    port map (
            O => \N__44172\,
            I => \N__44166\
        );

    \I__10438\ : InMux
    port map (
            O => \N__44169\,
            I => \N__44161\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__44166\,
            I => \N__44157\
        );

    \I__10436\ : InMux
    port map (
            O => \N__44165\,
            I => \N__44154\
        );

    \I__10435\ : CascadeMux
    port map (
            O => \N__44164\,
            I => \N__44151\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__44161\,
            I => \N__44148\
        );

    \I__10433\ : InMux
    port map (
            O => \N__44160\,
            I => \N__44145\
        );

    \I__10432\ : Span4Mux_v
    port map (
            O => \N__44157\,
            I => \N__44140\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__44154\,
            I => \N__44140\
        );

    \I__10430\ : InMux
    port map (
            O => \N__44151\,
            I => \N__44136\
        );

    \I__10429\ : Span4Mux_h
    port map (
            O => \N__44148\,
            I => \N__44133\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__44145\,
            I => \N__44130\
        );

    \I__10427\ : Span4Mux_h
    port map (
            O => \N__44140\,
            I => \N__44127\
        );

    \I__10426\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44124\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__44136\,
            I => \N__44121\
        );

    \I__10424\ : Odrv4
    port map (
            O => \N__44133\,
            I => rand_data_12
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__44130\,
            I => rand_data_12
        );

    \I__10422\ : Odrv4
    port map (
            O => \N__44127\,
            I => rand_data_12
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__44124\,
            I => rand_data_12
        );

    \I__10420\ : Odrv12
    port map (
            O => \N__44121\,
            I => rand_data_12
        );

    \I__10419\ : CascadeMux
    port map (
            O => \N__44110\,
            I => \N__44107\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44107\,
            I => \N__44103\
        );

    \I__10417\ : InMux
    port map (
            O => \N__44106\,
            I => \N__44100\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__44103\,
            I => \N__44097\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__44100\,
            I => data_out_frame2_17_4
        );

    \I__10414\ : Odrv4
    port map (
            O => \N__44097\,
            I => data_out_frame2_17_4
        );

    \I__10413\ : InMux
    port map (
            O => \N__44092\,
            I => \N__44087\
        );

    \I__10412\ : InMux
    port map (
            O => \N__44091\,
            I => \N__44082\
        );

    \I__10411\ : InMux
    port map (
            O => \N__44090\,
            I => \N__44082\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__44087\,
            I => \N__44078\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__44082\,
            I => \N__44075\
        );

    \I__10408\ : InMux
    port map (
            O => \N__44081\,
            I => \N__44072\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__44078\,
            I => \N__44069\
        );

    \I__10406\ : Span4Mux_v
    port map (
            O => \N__44075\,
            I => \N__44065\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__44072\,
            I => \N__44062\
        );

    \I__10404\ : Span4Mux_v
    port map (
            O => \N__44069\,
            I => \N__44059\
        );

    \I__10403\ : InMux
    port map (
            O => \N__44068\,
            I => \N__44056\
        );

    \I__10402\ : Span4Mux_h
    port map (
            O => \N__44065\,
            I => \N__44051\
        );

    \I__10401\ : Span4Mux_s2_v
    port map (
            O => \N__44062\,
            I => \N__44051\
        );

    \I__10400\ : Odrv4
    port map (
            O => \N__44059\,
            I => rand_data_23
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__44056\,
            I => rand_data_23
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__44051\,
            I => rand_data_23
        );

    \I__10397\ : InMux
    port map (
            O => \N__44044\,
            I => \N__44041\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__44041\,
            I => \N__44035\
        );

    \I__10395\ : InMux
    port map (
            O => \N__44040\,
            I => \N__44032\
        );

    \I__10394\ : InMux
    port map (
            O => \N__44039\,
            I => \N__44029\
        );

    \I__10393\ : InMux
    port map (
            O => \N__44038\,
            I => \N__44026\
        );

    \I__10392\ : Span4Mux_h
    port map (
            O => \N__44035\,
            I => \N__44019\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__44032\,
            I => \N__44019\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__44029\,
            I => \N__44019\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__44026\,
            I => data_out_frame2_6_7
        );

    \I__10388\ : Odrv4
    port map (
            O => \N__44019\,
            I => data_out_frame2_6_7
        );

    \I__10387\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44009\
        );

    \I__10386\ : InMux
    port map (
            O => \N__44013\,
            I => \N__44006\
        );

    \I__10385\ : InMux
    port map (
            O => \N__44012\,
            I => \N__44003\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__44009\,
            I => \N__43997\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__44006\,
            I => \N__43997\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__44003\,
            I => \N__43994\
        );

    \I__10381\ : InMux
    port map (
            O => \N__44002\,
            I => \N__43991\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__43997\,
            I => \N__43987\
        );

    \I__10379\ : Span4Mux_v
    port map (
            O => \N__43994\,
            I => \N__43984\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__43991\,
            I => \N__43981\
        );

    \I__10377\ : InMux
    port map (
            O => \N__43990\,
            I => \N__43978\
        );

    \I__10376\ : Span4Mux_v
    port map (
            O => \N__43987\,
            I => \N__43973\
        );

    \I__10375\ : Span4Mux_v
    port map (
            O => \N__43984\,
            I => \N__43973\
        );

    \I__10374\ : Span4Mux_s2_v
    port map (
            O => \N__43981\,
            I => \N__43970\
        );

    \I__10373\ : LocalMux
    port map (
            O => \N__43978\,
            I => rand_data_31
        );

    \I__10372\ : Odrv4
    port map (
            O => \N__43973\,
            I => rand_data_31
        );

    \I__10371\ : Odrv4
    port map (
            O => \N__43970\,
            I => rand_data_31
        );

    \I__10370\ : InMux
    port map (
            O => \N__43963\,
            I => \N__43960\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__43960\,
            I => \N__43955\
        );

    \I__10368\ : InMux
    port map (
            O => \N__43959\,
            I => \N__43952\
        );

    \I__10367\ : CascadeMux
    port map (
            O => \N__43958\,
            I => \N__43949\
        );

    \I__10366\ : Span4Mux_v
    port map (
            O => \N__43955\,
            I => \N__43944\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__43952\,
            I => \N__43941\
        );

    \I__10364\ : InMux
    port map (
            O => \N__43949\,
            I => \N__43938\
        );

    \I__10363\ : InMux
    port map (
            O => \N__43948\,
            I => \N__43935\
        );

    \I__10362\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43932\
        );

    \I__10361\ : Span4Mux_h
    port map (
            O => \N__43944\,
            I => \N__43929\
        );

    \I__10360\ : Span4Mux_h
    port map (
            O => \N__43941\,
            I => \N__43924\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__43938\,
            I => \N__43924\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__43935\,
            I => data_out_frame2_5_7
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__43932\,
            I => data_out_frame2_5_7
        );

    \I__10356\ : Odrv4
    port map (
            O => \N__43929\,
            I => data_out_frame2_5_7
        );

    \I__10355\ : Odrv4
    port map (
            O => \N__43924\,
            I => data_out_frame2_5_7
        );

    \I__10354\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43912\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__43912\,
            I => \c0.n24_adj_2272\
        );

    \I__10352\ : CascadeMux
    port map (
            O => \N__43909\,
            I => \N__43903\
        );

    \I__10351\ : CascadeMux
    port map (
            O => \N__43908\,
            I => \N__43899\
        );

    \I__10350\ : InMux
    port map (
            O => \N__43907\,
            I => \N__43896\
        );

    \I__10349\ : InMux
    port map (
            O => \N__43906\,
            I => \N__43891\
        );

    \I__10348\ : InMux
    port map (
            O => \N__43903\,
            I => \N__43891\
        );

    \I__10347\ : InMux
    port map (
            O => \N__43902\,
            I => \N__43888\
        );

    \I__10346\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43885\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__43896\,
            I => \N__43881\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__43891\,
            I => \N__43878\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__43888\,
            I => \N__43873\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__43885\,
            I => \N__43873\
        );

    \I__10341\ : InMux
    port map (
            O => \N__43884\,
            I => \N__43870\
        );

    \I__10340\ : Span4Mux_v
    port map (
            O => \N__43881\,
            I => \N__43867\
        );

    \I__10339\ : Span4Mux_v
    port map (
            O => \N__43878\,
            I => \N__43864\
        );

    \I__10338\ : Span4Mux_v
    port map (
            O => \N__43873\,
            I => \N__43861\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__43870\,
            I => \N__43852\
        );

    \I__10336\ : Span4Mux_h
    port map (
            O => \N__43867\,
            I => \N__43852\
        );

    \I__10335\ : Span4Mux_h
    port map (
            O => \N__43864\,
            I => \N__43852\
        );

    \I__10334\ : Span4Mux_v
    port map (
            O => \N__43861\,
            I => \N__43852\
        );

    \I__10333\ : Odrv4
    port map (
            O => \N__43852\,
            I => data_out_frame2_9_2
        );

    \I__10332\ : InMux
    port map (
            O => \N__43849\,
            I => \N__43844\
        );

    \I__10331\ : InMux
    port map (
            O => \N__43848\,
            I => \N__43841\
        );

    \I__10330\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43838\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__43844\,
            I => \N__43833\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__43841\,
            I => \N__43833\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__43838\,
            I => \N__43828\
        );

    \I__10326\ : Sp12to4
    port map (
            O => \N__43833\,
            I => \N__43825\
        );

    \I__10325\ : InMux
    port map (
            O => \N__43832\,
            I => \N__43822\
        );

    \I__10324\ : InMux
    port map (
            O => \N__43831\,
            I => \N__43819\
        );

    \I__10323\ : Span4Mux_h
    port map (
            O => \N__43828\,
            I => \N__43816\
        );

    \I__10322\ : Span12Mux_v
    port map (
            O => \N__43825\,
            I => \N__43811\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__43822\,
            I => \N__43811\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__43819\,
            I => data_out_frame2_16_0
        );

    \I__10319\ : Odrv4
    port map (
            O => \N__43816\,
            I => data_out_frame2_16_0
        );

    \I__10318\ : Odrv12
    port map (
            O => \N__43811\,
            I => data_out_frame2_16_0
        );

    \I__10317\ : InMux
    port map (
            O => \N__43804\,
            I => \N__43801\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__43801\,
            I => \N__43798\
        );

    \I__10315\ : Odrv4
    port map (
            O => \N__43798\,
            I => \c0.n9892\
        );

    \I__10314\ : CascadeMux
    port map (
            O => \N__43795\,
            I => \N__43792\
        );

    \I__10313\ : InMux
    port map (
            O => \N__43792\,
            I => \N__43789\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__43789\,
            I => \N__43786\
        );

    \I__10311\ : Odrv4
    port map (
            O => \N__43786\,
            I => \c0.n20_adj_2205\
        );

    \I__10310\ : InMux
    port map (
            O => \N__43783\,
            I => \N__43780\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__43780\,
            I => \N__43777\
        );

    \I__10308\ : Odrv12
    port map (
            O => \N__43777\,
            I => \c0.n18071\
        );

    \I__10307\ : CascadeMux
    port map (
            O => \N__43774\,
            I => \c0.n18074_cascade_\
        );

    \I__10306\ : InMux
    port map (
            O => \N__43771\,
            I => \N__43768\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__43768\,
            I => \N__43763\
        );

    \I__10304\ : InMux
    port map (
            O => \N__43767\,
            I => \N__43760\
        );

    \I__10303\ : InMux
    port map (
            O => \N__43766\,
            I => \N__43757\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__43763\,
            I => \N__43753\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__43760\,
            I => \N__43750\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__43757\,
            I => \N__43747\
        );

    \I__10299\ : InMux
    port map (
            O => \N__43756\,
            I => \N__43744\
        );

    \I__10298\ : Span4Mux_h
    port map (
            O => \N__43753\,
            I => \N__43739\
        );

    \I__10297\ : Span4Mux_v
    port map (
            O => \N__43750\,
            I => \N__43739\
        );

    \I__10296\ : Odrv12
    port map (
            O => \N__43747\,
            I => data_out_frame2_12_7
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__43744\,
            I => data_out_frame2_12_7
        );

    \I__10294\ : Odrv4
    port map (
            O => \N__43739\,
            I => data_out_frame2_12_7
        );

    \I__10293\ : InMux
    port map (
            O => \N__43732\,
            I => \N__43729\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__43729\,
            I => \N__43725\
        );

    \I__10291\ : CascadeMux
    port map (
            O => \N__43728\,
            I => \N__43721\
        );

    \I__10290\ : Span4Mux_v
    port map (
            O => \N__43725\,
            I => \N__43718\
        );

    \I__10289\ : InMux
    port map (
            O => \N__43724\,
            I => \N__43715\
        );

    \I__10288\ : InMux
    port map (
            O => \N__43721\,
            I => \N__43712\
        );

    \I__10287\ : Span4Mux_h
    port map (
            O => \N__43718\,
            I => \N__43709\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__43715\,
            I => \N__43704\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__43712\,
            I => \N__43704\
        );

    \I__10284\ : Odrv4
    port map (
            O => \N__43709\,
            I => data_out_frame2_13_7
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__43704\,
            I => data_out_frame2_13_7
        );

    \I__10282\ : CascadeMux
    port map (
            O => \N__43699\,
            I => \c0.n18065_cascade_\
        );

    \I__10281\ : InMux
    port map (
            O => \N__43696\,
            I => \N__43693\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__43693\,
            I => \c0.n18068\
        );

    \I__10279\ : InMux
    port map (
            O => \N__43690\,
            I => \N__43687\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__43687\,
            I => \N__43683\
        );

    \I__10277\ : InMux
    port map (
            O => \N__43686\,
            I => \N__43679\
        );

    \I__10276\ : Span4Mux_h
    port map (
            O => \N__43683\,
            I => \N__43675\
        );

    \I__10275\ : InMux
    port map (
            O => \N__43682\,
            I => \N__43672\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__43679\,
            I => \N__43669\
        );

    \I__10273\ : InMux
    port map (
            O => \N__43678\,
            I => \N__43666\
        );

    \I__10272\ : Sp12to4
    port map (
            O => \N__43675\,
            I => \N__43663\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__43672\,
            I => \N__43658\
        );

    \I__10270\ : Span4Mux_h
    port map (
            O => \N__43669\,
            I => \N__43658\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__43666\,
            I => data_out_frame2_14_6
        );

    \I__10268\ : Odrv12
    port map (
            O => \N__43663\,
            I => data_out_frame2_14_6
        );

    \I__10267\ : Odrv4
    port map (
            O => \N__43658\,
            I => data_out_frame2_14_6
        );

    \I__10266\ : InMux
    port map (
            O => \N__43651\,
            I => \N__43648\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__43648\,
            I => \N__43643\
        );

    \I__10264\ : InMux
    port map (
            O => \N__43647\,
            I => \N__43640\
        );

    \I__10263\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43637\
        );

    \I__10262\ : Span4Mux_h
    port map (
            O => \N__43643\,
            I => \N__43633\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__43640\,
            I => \N__43630\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__43637\,
            I => \N__43627\
        );

    \I__10259\ : InMux
    port map (
            O => \N__43636\,
            I => \N__43623\
        );

    \I__10258\ : Span4Mux_v
    port map (
            O => \N__43633\,
            I => \N__43620\
        );

    \I__10257\ : Span4Mux_h
    port map (
            O => \N__43630\,
            I => \N__43617\
        );

    \I__10256\ : Span4Mux_h
    port map (
            O => \N__43627\,
            I => \N__43614\
        );

    \I__10255\ : InMux
    port map (
            O => \N__43626\,
            I => \N__43611\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__43623\,
            I => data_out_frame2_12_6
        );

    \I__10253\ : Odrv4
    port map (
            O => \N__43620\,
            I => data_out_frame2_12_6
        );

    \I__10252\ : Odrv4
    port map (
            O => \N__43617\,
            I => data_out_frame2_12_6
        );

    \I__10251\ : Odrv4
    port map (
            O => \N__43614\,
            I => data_out_frame2_12_6
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__43611\,
            I => data_out_frame2_12_6
        );

    \I__10249\ : CascadeMux
    port map (
            O => \N__43600\,
            I => \c0.n18005_cascade_\
        );

    \I__10248\ : CascadeMux
    port map (
            O => \N__43597\,
            I => \N__43594\
        );

    \I__10247\ : InMux
    port map (
            O => \N__43594\,
            I => \N__43591\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__43591\,
            I => \N__43588\
        );

    \I__10245\ : Odrv4
    port map (
            O => \N__43588\,
            I => \c0.n18008\
        );

    \I__10244\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43581\
        );

    \I__10243\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43578\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__43581\,
            I => \N__43575\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__43578\,
            I => \N__43569\
        );

    \I__10240\ : Span4Mux_v
    port map (
            O => \N__43575\,
            I => \N__43566\
        );

    \I__10239\ : InMux
    port map (
            O => \N__43574\,
            I => \N__43563\
        );

    \I__10238\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43560\
        );

    \I__10237\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43557\
        );

    \I__10236\ : Span4Mux_v
    port map (
            O => \N__43569\,
            I => \N__43554\
        );

    \I__10235\ : Span4Mux_h
    port map (
            O => \N__43566\,
            I => \N__43549\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__43563\,
            I => \N__43549\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__43560\,
            I => \N__43546\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__43557\,
            I => data_out_frame2_10_0
        );

    \I__10231\ : Odrv4
    port map (
            O => \N__43554\,
            I => data_out_frame2_10_0
        );

    \I__10230\ : Odrv4
    port map (
            O => \N__43549\,
            I => data_out_frame2_10_0
        );

    \I__10229\ : Odrv4
    port map (
            O => \N__43546\,
            I => data_out_frame2_10_0
        );

    \I__10228\ : InMux
    port map (
            O => \N__43537\,
            I => \N__43534\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__43534\,
            I => \N__43531\
        );

    \I__10226\ : Span4Mux_v
    port map (
            O => \N__43531\,
            I => \N__43528\
        );

    \I__10225\ : Odrv4
    port map (
            O => \N__43528\,
            I => \c0.n17347\
        );

    \I__10224\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43520\
        );

    \I__10223\ : InMux
    port map (
            O => \N__43524\,
            I => \N__43516\
        );

    \I__10222\ : InMux
    port map (
            O => \N__43523\,
            I => \N__43513\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__43520\,
            I => \N__43510\
        );

    \I__10220\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43507\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__43516\,
            I => \N__43504\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__43513\,
            I => \N__43501\
        );

    \I__10217\ : Span4Mux_h
    port map (
            O => \N__43510\,
            I => \N__43498\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__43507\,
            I => data_out_frame2_5_4
        );

    \I__10215\ : Odrv4
    port map (
            O => \N__43504\,
            I => data_out_frame2_5_4
        );

    \I__10214\ : Odrv12
    port map (
            O => \N__43501\,
            I => data_out_frame2_5_4
        );

    \I__10213\ : Odrv4
    port map (
            O => \N__43498\,
            I => data_out_frame2_5_4
        );

    \I__10212\ : InMux
    port map (
            O => \N__43489\,
            I => \N__43486\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__43486\,
            I => \N__43483\
        );

    \I__10210\ : Span4Mux_v
    port map (
            O => \N__43483\,
            I => \N__43480\
        );

    \I__10209\ : Odrv4
    port map (
            O => \N__43480\,
            I => \c0.n17495\
        );

    \I__10208\ : InMux
    port map (
            O => \N__43477\,
            I => \N__43474\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__43474\,
            I => \N__43469\
        );

    \I__10206\ : InMux
    port map (
            O => \N__43473\,
            I => \N__43466\
        );

    \I__10205\ : InMux
    port map (
            O => \N__43472\,
            I => \N__43460\
        );

    \I__10204\ : Span4Mux_v
    port map (
            O => \N__43469\,
            I => \N__43457\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__43466\,
            I => \N__43454\
        );

    \I__10202\ : InMux
    port map (
            O => \N__43465\,
            I => \N__43451\
        );

    \I__10201\ : InMux
    port map (
            O => \N__43464\,
            I => \N__43448\
        );

    \I__10200\ : InMux
    port map (
            O => \N__43463\,
            I => \N__43445\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__43460\,
            I => \N__43438\
        );

    \I__10198\ : Span4Mux_h
    port map (
            O => \N__43457\,
            I => \N__43438\
        );

    \I__10197\ : Span4Mux_v
    port map (
            O => \N__43454\,
            I => \N__43438\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__43451\,
            I => \N__43433\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__43448\,
            I => \N__43433\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__43445\,
            I => \N__43430\
        );

    \I__10193\ : Sp12to4
    port map (
            O => \N__43438\,
            I => \N__43427\
        );

    \I__10192\ : Span4Mux_h
    port map (
            O => \N__43433\,
            I => \N__43424\
        );

    \I__10191\ : Odrv12
    port map (
            O => \N__43430\,
            I => data_out_frame2_9_6
        );

    \I__10190\ : Odrv12
    port map (
            O => \N__43427\,
            I => data_out_frame2_9_6
        );

    \I__10189\ : Odrv4
    port map (
            O => \N__43424\,
            I => data_out_frame2_9_6
        );

    \I__10188\ : InMux
    port map (
            O => \N__43417\,
            I => \N__43414\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__43414\,
            I => \c0.n18047\
        );

    \I__10186\ : InMux
    port map (
            O => \N__43411\,
            I => \N__43407\
        );

    \I__10185\ : InMux
    port map (
            O => \N__43410\,
            I => \N__43404\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__43407\,
            I => \N__43401\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__43404\,
            I => \N__43398\
        );

    \I__10182\ : Span4Mux_h
    port map (
            O => \N__43401\,
            I => \N__43395\
        );

    \I__10181\ : Span4Mux_v
    port map (
            O => \N__43398\,
            I => \N__43392\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__43395\,
            I => \c0.n9859\
        );

    \I__10179\ : Odrv4
    port map (
            O => \N__43392\,
            I => \c0.n9859\
        );

    \I__10178\ : CascadeMux
    port map (
            O => \N__43387\,
            I => \N__43384\
        );

    \I__10177\ : InMux
    port map (
            O => \N__43384\,
            I => \N__43381\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43377\
        );

    \I__10175\ : InMux
    port map (
            O => \N__43380\,
            I => \N__43374\
        );

    \I__10174\ : Span4Mux_v
    port map (
            O => \N__43377\,
            I => \N__43369\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__43374\,
            I => \N__43366\
        );

    \I__10172\ : InMux
    port map (
            O => \N__43373\,
            I => \N__43363\
        );

    \I__10171\ : InMux
    port map (
            O => \N__43372\,
            I => \N__43360\
        );

    \I__10170\ : Span4Mux_v
    port map (
            O => \N__43369\,
            I => \N__43357\
        );

    \I__10169\ : Span4Mux_v
    port map (
            O => \N__43366\,
            I => \N__43354\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__43363\,
            I => \N__43351\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__43360\,
            I => \N__43346\
        );

    \I__10166\ : Span4Mux_h
    port map (
            O => \N__43357\,
            I => \N__43346\
        );

    \I__10165\ : Span4Mux_h
    port map (
            O => \N__43354\,
            I => \N__43341\
        );

    \I__10164\ : Span4Mux_v
    port map (
            O => \N__43351\,
            I => \N__43341\
        );

    \I__10163\ : Odrv4
    port map (
            O => \N__43346\,
            I => data_out_frame2_13_2
        );

    \I__10162\ : Odrv4
    port map (
            O => \N__43341\,
            I => data_out_frame2_13_2
        );

    \I__10161\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43332\
        );

    \I__10160\ : InMux
    port map (
            O => \N__43335\,
            I => \N__43329\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__43332\,
            I => \N__43324\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__43329\,
            I => \N__43324\
        );

    \I__10157\ : Span4Mux_h
    port map (
            O => \N__43324\,
            I => \N__43321\
        );

    \I__10156\ : Odrv4
    port map (
            O => \N__43321\,
            I => \c0.n17133\
        );

    \I__10155\ : InMux
    port map (
            O => \N__43318\,
            I => \N__43315\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__43315\,
            I => \N__43312\
        );

    \I__10153\ : Odrv4
    port map (
            O => \N__43312\,
            I => \c0.n27_adj_2277\
        );

    \I__10152\ : InMux
    port map (
            O => \N__43309\,
            I => \N__43306\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__43306\,
            I => \N__43301\
        );

    \I__10150\ : CascadeMux
    port map (
            O => \N__43305\,
            I => \N__43297\
        );

    \I__10149\ : InMux
    port map (
            O => \N__43304\,
            I => \N__43294\
        );

    \I__10148\ : Span4Mux_v
    port map (
            O => \N__43301\,
            I => \N__43291\
        );

    \I__10147\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43286\
        );

    \I__10146\ : InMux
    port map (
            O => \N__43297\,
            I => \N__43286\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__43294\,
            I => data_out_frame2_8_6
        );

    \I__10144\ : Odrv4
    port map (
            O => \N__43291\,
            I => data_out_frame2_8_6
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__43286\,
            I => data_out_frame2_8_6
        );

    \I__10142\ : InMux
    port map (
            O => \N__43279\,
            I => \N__43274\
        );

    \I__10141\ : InMux
    port map (
            O => \N__43278\,
            I => \N__43271\
        );

    \I__10140\ : InMux
    port map (
            O => \N__43277\,
            I => \N__43268\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__43274\,
            I => \N__43263\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__43271\,
            I => \N__43258\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__43268\,
            I => \N__43258\
        );

    \I__10136\ : CascadeMux
    port map (
            O => \N__43267\,
            I => \N__43255\
        );

    \I__10135\ : InMux
    port map (
            O => \N__43266\,
            I => \N__43252\
        );

    \I__10134\ : Span4Mux_h
    port map (
            O => \N__43263\,
            I => \N__43247\
        );

    \I__10133\ : Span4Mux_h
    port map (
            O => \N__43258\,
            I => \N__43247\
        );

    \I__10132\ : InMux
    port map (
            O => \N__43255\,
            I => \N__43244\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__43252\,
            I => data_out_frame2_6_6
        );

    \I__10130\ : Odrv4
    port map (
            O => \N__43247\,
            I => data_out_frame2_6_6
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__43244\,
            I => data_out_frame2_6_6
        );

    \I__10128\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43234\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__43234\,
            I => \c0.n18050\
        );

    \I__10126\ : InMux
    port map (
            O => \N__43231\,
            I => \N__43228\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__43228\,
            I => \N__43224\
        );

    \I__10124\ : InMux
    port map (
            O => \N__43227\,
            I => \N__43221\
        );

    \I__10123\ : Odrv4
    port map (
            O => \N__43224\,
            I => \c0.n9671\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__43221\,
            I => \c0.n9671\
        );

    \I__10121\ : InMux
    port map (
            O => \N__43216\,
            I => \N__43212\
        );

    \I__10120\ : InMux
    port map (
            O => \N__43215\,
            I => \N__43209\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__43212\,
            I => \c0.n17016\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__43209\,
            I => \c0.n17016\
        );

    \I__10117\ : InMux
    port map (
            O => \N__43204\,
            I => \N__43201\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__43201\,
            I => \N__43198\
        );

    \I__10115\ : Span4Mux_h
    port map (
            O => \N__43198\,
            I => \N__43195\
        );

    \I__10114\ : Span4Mux_h
    port map (
            O => \N__43195\,
            I => \N__43192\
        );

    \I__10113\ : Odrv4
    port map (
            O => \N__43192\,
            I => \c0.n6_adj_2293\
        );

    \I__10112\ : InMux
    port map (
            O => \N__43189\,
            I => \N__43186\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__43186\,
            I => \N__43183\
        );

    \I__10110\ : Span4Mux_h
    port map (
            O => \N__43183\,
            I => \N__43179\
        );

    \I__10109\ : InMux
    port map (
            O => \N__43182\,
            I => \N__43176\
        );

    \I__10108\ : Odrv4
    port map (
            O => \N__43179\,
            I => \c0.n16960\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__43176\,
            I => \c0.n16960\
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__43171\,
            I => \c0.n18017_cascade_\
        );

    \I__10105\ : InMux
    port map (
            O => \N__43168\,
            I => \N__43165\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__43165\,
            I => \c0.n17593\
        );

    \I__10103\ : InMux
    port map (
            O => \N__43162\,
            I => \N__43159\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__43159\,
            I => \c0.n10_adj_2154\
        );

    \I__10101\ : CascadeMux
    port map (
            O => \N__43156\,
            I => \c0.n18020_cascade_\
        );

    \I__10100\ : InMux
    port map (
            O => \N__43153\,
            I => \N__43143\
        );

    \I__10099\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43140\
        );

    \I__10098\ : InMux
    port map (
            O => \N__43151\,
            I => \N__43136\
        );

    \I__10097\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43133\
        );

    \I__10096\ : InMux
    port map (
            O => \N__43149\,
            I => \N__43130\
        );

    \I__10095\ : InMux
    port map (
            O => \N__43148\,
            I => \N__43127\
        );

    \I__10094\ : InMux
    port map (
            O => \N__43147\,
            I => \N__43124\
        );

    \I__10093\ : InMux
    port map (
            O => \N__43146\,
            I => \N__43121\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__43143\,
            I => \N__43116\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__43140\,
            I => \N__43113\
        );

    \I__10090\ : CascadeMux
    port map (
            O => \N__43139\,
            I => \N__43109\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__43136\,
            I => \N__43106\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__43133\,
            I => \N__43103\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__43130\,
            I => \N__43096\
        );

    \I__10086\ : LocalMux
    port map (
            O => \N__43127\,
            I => \N__43096\
        );

    \I__10085\ : LocalMux
    port map (
            O => \N__43124\,
            I => \N__43096\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__43121\,
            I => \N__43093\
        );

    \I__10083\ : InMux
    port map (
            O => \N__43120\,
            I => \N__43090\
        );

    \I__10082\ : InMux
    port map (
            O => \N__43119\,
            I => \N__43087\
        );

    \I__10081\ : Span4Mux_v
    port map (
            O => \N__43116\,
            I => \N__43082\
        );

    \I__10080\ : Span4Mux_v
    port map (
            O => \N__43113\,
            I => \N__43082\
        );

    \I__10079\ : InMux
    port map (
            O => \N__43112\,
            I => \N__43079\
        );

    \I__10078\ : InMux
    port map (
            O => \N__43109\,
            I => \N__43075\
        );

    \I__10077\ : Span4Mux_s1_v
    port map (
            O => \N__43106\,
            I => \N__43072\
        );

    \I__10076\ : Span4Mux_h
    port map (
            O => \N__43103\,
            I => \N__43069\
        );

    \I__10075\ : Span4Mux_v
    port map (
            O => \N__43096\,
            I => \N__43064\
        );

    \I__10074\ : Span4Mux_s1_v
    port map (
            O => \N__43093\,
            I => \N__43064\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__43090\,
            I => \N__43055\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__43087\,
            I => \N__43055\
        );

    \I__10071\ : Sp12to4
    port map (
            O => \N__43082\,
            I => \N__43055\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__43079\,
            I => \N__43055\
        );

    \I__10069\ : InMux
    port map (
            O => \N__43078\,
            I => \N__43052\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__43075\,
            I => byte_transmit_counter_3
        );

    \I__10067\ : Odrv4
    port map (
            O => \N__43072\,
            I => byte_transmit_counter_3
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__43069\,
            I => byte_transmit_counter_3
        );

    \I__10065\ : Odrv4
    port map (
            O => \N__43064\,
            I => byte_transmit_counter_3
        );

    \I__10064\ : Odrv12
    port map (
            O => \N__43055\,
            I => byte_transmit_counter_3
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__43052\,
            I => byte_transmit_counter_3
        );

    \I__10062\ : InMux
    port map (
            O => \N__43039\,
            I => \N__43036\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__43036\,
            I => \N__43033\
        );

    \I__10060\ : Odrv12
    port map (
            O => \N__43033\,
            I => \c0.n10_adj_2155\
        );

    \I__10059\ : InMux
    port map (
            O => \N__43030\,
            I => \N__43027\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__43027\,
            I => \N__43024\
        );

    \I__10057\ : Odrv4
    port map (
            O => \N__43024\,
            I => \c0.n10_adj_2268\
        );

    \I__10056\ : InMux
    port map (
            O => \N__43021\,
            I => \N__43017\
        );

    \I__10055\ : InMux
    port map (
            O => \N__43020\,
            I => \N__43014\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__43017\,
            I => \N__43008\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__43014\,
            I => \N__43005\
        );

    \I__10052\ : InMux
    port map (
            O => \N__43013\,
            I => \N__43002\
        );

    \I__10051\ : InMux
    port map (
            O => \N__43012\,
            I => \N__42999\
        );

    \I__10050\ : InMux
    port map (
            O => \N__43011\,
            I => \N__42996\
        );

    \I__10049\ : Span4Mux_s3_v
    port map (
            O => \N__43008\,
            I => \N__42989\
        );

    \I__10048\ : Span4Mux_v
    port map (
            O => \N__43005\,
            I => \N__42989\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__43002\,
            I => \N__42989\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__42999\,
            I => \c0.data_out_8_3\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__42996\,
            I => \c0.data_out_8_3\
        );

    \I__10044\ : Odrv4
    port map (
            O => \N__42989\,
            I => \c0.data_out_8_3\
        );

    \I__10043\ : CascadeMux
    port map (
            O => \N__42982\,
            I => \N__42978\
        );

    \I__10042\ : InMux
    port map (
            O => \N__42981\,
            I => \N__42975\
        );

    \I__10041\ : InMux
    port map (
            O => \N__42978\,
            I => \N__42972\
        );

    \I__10040\ : LocalMux
    port map (
            O => \N__42975\,
            I => \N__42969\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__42972\,
            I => \N__42965\
        );

    \I__10038\ : Span4Mux_s3_v
    port map (
            O => \N__42969\,
            I => \N__42962\
        );

    \I__10037\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42959\
        );

    \I__10036\ : Span4Mux_h
    port map (
            O => \N__42965\,
            I => \N__42954\
        );

    \I__10035\ : Span4Mux_h
    port map (
            O => \N__42962\,
            I => \N__42949\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__42959\,
            I => \N__42949\
        );

    \I__10033\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42944\
        );

    \I__10032\ : InMux
    port map (
            O => \N__42957\,
            I => \N__42944\
        );

    \I__10031\ : Odrv4
    port map (
            O => \N__42954\,
            I => data_out_8_4
        );

    \I__10030\ : Odrv4
    port map (
            O => \N__42949\,
            I => data_out_8_4
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__42944\,
            I => data_out_8_4
        );

    \I__10028\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42933\
        );

    \I__10027\ : InMux
    port map (
            O => \N__42936\,
            I => \N__42930\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__42933\,
            I => \N__42927\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__42930\,
            I => \N__42922\
        );

    \I__10024\ : Span4Mux_s2_v
    port map (
            O => \N__42927\,
            I => \N__42922\
        );

    \I__10023\ : Span4Mux_h
    port map (
            O => \N__42922\,
            I => \N__42918\
        );

    \I__10022\ : InMux
    port map (
            O => \N__42921\,
            I => \N__42915\
        );

    \I__10021\ : Odrv4
    port map (
            O => \N__42918\,
            I => \c0.data_out_9_1\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__42915\,
            I => \c0.data_out_9_1\
        );

    \I__10019\ : InMux
    port map (
            O => \N__42910\,
            I => \N__42906\
        );

    \I__10018\ : InMux
    port map (
            O => \N__42909\,
            I => \N__42903\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__42906\,
            I => data_out_3_4
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__42903\,
            I => data_out_3_4
        );

    \I__10015\ : InMux
    port map (
            O => \N__42898\,
            I => \N__42895\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__42895\,
            I => \N__42892\
        );

    \I__10013\ : Span4Mux_s2_v
    port map (
            O => \N__42892\,
            I => \N__42889\
        );

    \I__10012\ : Span4Mux_h
    port map (
            O => \N__42889\,
            I => \N__42886\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__42886\,
            I => \c0.n17591\
        );

    \I__10010\ : InMux
    port map (
            O => \N__42883\,
            I => \N__42879\
        );

    \I__10009\ : CascadeMux
    port map (
            O => \N__42882\,
            I => \N__42876\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__42879\,
            I => \N__42873\
        );

    \I__10007\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42870\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__42873\,
            I => rand_setpoint_16
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__42870\,
            I => rand_setpoint_16
        );

    \I__10004\ : InMux
    port map (
            O => \N__42865\,
            I => \N__42855\
        );

    \I__10003\ : InMux
    port map (
            O => \N__42864\,
            I => \N__42855\
        );

    \I__10002\ : InMux
    port map (
            O => \N__42863\,
            I => \N__42852\
        );

    \I__10001\ : CascadeMux
    port map (
            O => \N__42862\,
            I => \N__42848\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__42861\,
            I => \N__42844\
        );

    \I__9999\ : CascadeMux
    port map (
            O => \N__42860\,
            I => \N__42839\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__42855\,
            I => \N__42835\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__42852\,
            I => \N__42832\
        );

    \I__9996\ : InMux
    port map (
            O => \N__42851\,
            I => \N__42829\
        );

    \I__9995\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42826\
        );

    \I__9994\ : InMux
    port map (
            O => \N__42847\,
            I => \N__42823\
        );

    \I__9993\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42817\
        );

    \I__9992\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42817\
        );

    \I__9991\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42812\
        );

    \I__9990\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42812\
        );

    \I__9989\ : InMux
    port map (
            O => \N__42838\,
            I => \N__42809\
        );

    \I__9988\ : Span4Mux_s3_v
    port map (
            O => \N__42835\,
            I => \N__42804\
        );

    \I__9987\ : Span4Mux_s3_v
    port map (
            O => \N__42832\,
            I => \N__42804\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__42829\,
            I => \N__42799\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__42826\,
            I => \N__42799\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__42823\,
            I => \N__42795\
        );

    \I__9983\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42792\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__42817\,
            I => \N__42781\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__42812\,
            I => \N__42781\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__42809\,
            I => \N__42781\
        );

    \I__9979\ : Span4Mux_v
    port map (
            O => \N__42804\,
            I => \N__42781\
        );

    \I__9978\ : Span4Mux_s3_v
    port map (
            O => \N__42799\,
            I => \N__42781\
        );

    \I__9977\ : InMux
    port map (
            O => \N__42798\,
            I => \N__42778\
        );

    \I__9976\ : Span4Mux_v
    port map (
            O => \N__42795\,
            I => \N__42775\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__42792\,
            I => \N__42770\
        );

    \I__9974\ : Span4Mux_h
    port map (
            O => \N__42781\,
            I => \N__42770\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__42778\,
            I => n2547
        );

    \I__9972\ : Odrv4
    port map (
            O => \N__42775\,
            I => n2547
        );

    \I__9971\ : Odrv4
    port map (
            O => \N__42770\,
            I => n2547
        );

    \I__9970\ : CascadeMux
    port map (
            O => \N__42763\,
            I => \N__42755\
        );

    \I__9969\ : CascadeMux
    port map (
            O => \N__42762\,
            I => \N__42746\
        );

    \I__9968\ : CascadeMux
    port map (
            O => \N__42761\,
            I => \N__42742\
        );

    \I__9967\ : InMux
    port map (
            O => \N__42760\,
            I => \N__42739\
        );

    \I__9966\ : InMux
    port map (
            O => \N__42759\,
            I => \N__42736\
        );

    \I__9965\ : InMux
    port map (
            O => \N__42758\,
            I => \N__42733\
        );

    \I__9964\ : InMux
    port map (
            O => \N__42755\,
            I => \N__42728\
        );

    \I__9963\ : InMux
    port map (
            O => \N__42754\,
            I => \N__42728\
        );

    \I__9962\ : InMux
    port map (
            O => \N__42753\,
            I => \N__42722\
        );

    \I__9961\ : InMux
    port map (
            O => \N__42752\,
            I => \N__42719\
        );

    \I__9960\ : CascadeMux
    port map (
            O => \N__42751\,
            I => \N__42716\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__42750\,
            I => \N__42713\
        );

    \I__9958\ : CascadeMux
    port map (
            O => \N__42749\,
            I => \N__42705\
        );

    \I__9957\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42702\
        );

    \I__9956\ : InMux
    port map (
            O => \N__42745\,
            I => \N__42698\
        );

    \I__9955\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42695\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__42739\,
            I => \N__42692\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__42736\,
            I => \N__42687\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__42733\,
            I => \N__42687\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__42728\,
            I => \N__42684\
        );

    \I__9950\ : InMux
    port map (
            O => \N__42727\,
            I => \N__42681\
        );

    \I__9949\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42675\
        );

    \I__9948\ : InMux
    port map (
            O => \N__42725\,
            I => \N__42675\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__42722\,
            I => \N__42670\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__42719\,
            I => \N__42670\
        );

    \I__9945\ : InMux
    port map (
            O => \N__42716\,
            I => \N__42661\
        );

    \I__9944\ : InMux
    port map (
            O => \N__42713\,
            I => \N__42661\
        );

    \I__9943\ : InMux
    port map (
            O => \N__42712\,
            I => \N__42661\
        );

    \I__9942\ : InMux
    port map (
            O => \N__42711\,
            I => \N__42661\
        );

    \I__9941\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42657\
        );

    \I__9940\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42654\
        );

    \I__9939\ : CascadeMux
    port map (
            O => \N__42708\,
            I => \N__42649\
        );

    \I__9938\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42641\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__42702\,
            I => \N__42638\
        );

    \I__9936\ : InMux
    port map (
            O => \N__42701\,
            I => \N__42635\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__42698\,
            I => \N__42624\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__42695\,
            I => \N__42624\
        );

    \I__9933\ : Span4Mux_s3_v
    port map (
            O => \N__42692\,
            I => \N__42624\
        );

    \I__9932\ : Span4Mux_s3_v
    port map (
            O => \N__42687\,
            I => \N__42624\
        );

    \I__9931\ : Span4Mux_v
    port map (
            O => \N__42684\,
            I => \N__42624\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__42681\,
            I => \N__42619\
        );

    \I__9929\ : InMux
    port map (
            O => \N__42680\,
            I => \N__42616\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__42675\,
            I => \N__42611\
        );

    \I__9927\ : Span4Mux_v
    port map (
            O => \N__42670\,
            I => \N__42611\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__42661\,
            I => \N__42608\
        );

    \I__9925\ : CascadeMux
    port map (
            O => \N__42660\,
            I => \N__42604\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__42657\,
            I => \N__42598\
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__42654\,
            I => \N__42598\
        );

    \I__9922\ : InMux
    port map (
            O => \N__42653\,
            I => \N__42593\
        );

    \I__9921\ : InMux
    port map (
            O => \N__42652\,
            I => \N__42593\
        );

    \I__9920\ : InMux
    port map (
            O => \N__42649\,
            I => \N__42589\
        );

    \I__9919\ : InMux
    port map (
            O => \N__42648\,
            I => \N__42584\
        );

    \I__9918\ : InMux
    port map (
            O => \N__42647\,
            I => \N__42584\
        );

    \I__9917\ : InMux
    port map (
            O => \N__42646\,
            I => \N__42581\
        );

    \I__9916\ : CascadeMux
    port map (
            O => \N__42645\,
            I => \N__42577\
        );

    \I__9915\ : InMux
    port map (
            O => \N__42644\,
            I => \N__42571\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__42641\,
            I => \N__42568\
        );

    \I__9913\ : Span4Mux_h
    port map (
            O => \N__42638\,
            I => \N__42561\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__42635\,
            I => \N__42561\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__42624\,
            I => \N__42561\
        );

    \I__9910\ : CascadeMux
    port map (
            O => \N__42623\,
            I => \N__42558\
        );

    \I__9909\ : CascadeMux
    port map (
            O => \N__42622\,
            I => \N__42555\
        );

    \I__9908\ : Span4Mux_h
    port map (
            O => \N__42619\,
            I => \N__42546\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__42616\,
            I => \N__42546\
        );

    \I__9906\ : Span4Mux_s2_v
    port map (
            O => \N__42611\,
            I => \N__42546\
        );

    \I__9905\ : Span4Mux_s2_v
    port map (
            O => \N__42608\,
            I => \N__42546\
        );

    \I__9904\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42543\
        );

    \I__9903\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42538\
        );

    \I__9902\ : InMux
    port map (
            O => \N__42603\,
            I => \N__42538\
        );

    \I__9901\ : Span4Mux_v
    port map (
            O => \N__42598\,
            I => \N__42533\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__42593\,
            I => \N__42533\
        );

    \I__9899\ : InMux
    port map (
            O => \N__42592\,
            I => \N__42530\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__42589\,
            I => \N__42525\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__42584\,
            I => \N__42525\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__42581\,
            I => \N__42522\
        );

    \I__9895\ : InMux
    port map (
            O => \N__42580\,
            I => \N__42515\
        );

    \I__9894\ : InMux
    port map (
            O => \N__42577\,
            I => \N__42515\
        );

    \I__9893\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42515\
        );

    \I__9892\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42510\
        );

    \I__9891\ : InMux
    port map (
            O => \N__42574\,
            I => \N__42510\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__42571\,
            I => \N__42503\
        );

    \I__9889\ : Span4Mux_h
    port map (
            O => \N__42568\,
            I => \N__42503\
        );

    \I__9888\ : Span4Mux_h
    port map (
            O => \N__42561\,
            I => \N__42503\
        );

    \I__9887\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42498\
        );

    \I__9886\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42498\
        );

    \I__9885\ : Span4Mux_h
    port map (
            O => \N__42546\,
            I => \N__42495\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__42543\,
            I => \N__42484\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__42538\,
            I => \N__42484\
        );

    \I__9882\ : Sp12to4
    port map (
            O => \N__42533\,
            I => \N__42484\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__42530\,
            I => \N__42484\
        );

    \I__9880\ : Span12Mux_v
    port map (
            O => \N__42525\,
            I => \N__42484\
        );

    \I__9879\ : Odrv4
    port map (
            O => \N__42522\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__42515\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__42510\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__9876\ : Odrv4
    port map (
            O => \N__42503\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__42498\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__9874\ : Odrv4
    port map (
            O => \N__42495\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__9873\ : Odrv12
    port map (
            O => \N__42484\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__9872\ : InMux
    port map (
            O => \N__42469\,
            I => \N__42461\
        );

    \I__9871\ : InMux
    port map (
            O => \N__42468\,
            I => \N__42458\
        );

    \I__9870\ : InMux
    port map (
            O => \N__42467\,
            I => \N__42455\
        );

    \I__9869\ : InMux
    port map (
            O => \N__42466\,
            I => \N__42452\
        );

    \I__9868\ : InMux
    port map (
            O => \N__42465\,
            I => \N__42449\
        );

    \I__9867\ : InMux
    port map (
            O => \N__42464\,
            I => \N__42446\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__42461\,
            I => \N__42443\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__42458\,
            I => \N__42440\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__42455\,
            I => \N__42436\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__42452\,
            I => \N__42431\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__42449\,
            I => \N__42431\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__42446\,
            I => \N__42428\
        );

    \I__9860\ : Span4Mux_v
    port map (
            O => \N__42443\,
            I => \N__42425\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__42440\,
            I => \N__42422\
        );

    \I__9858\ : InMux
    port map (
            O => \N__42439\,
            I => \N__42419\
        );

    \I__9857\ : Span4Mux_h
    port map (
            O => \N__42436\,
            I => \N__42414\
        );

    \I__9856\ : Span4Mux_h
    port map (
            O => \N__42431\,
            I => \N__42414\
        );

    \I__9855\ : Odrv12
    port map (
            O => \N__42428\,
            I => \c0.data_out_5_3\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__42425\,
            I => \c0.data_out_5_3\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__42422\,
            I => \c0.data_out_5_3\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__42419\,
            I => \c0.data_out_5_3\
        );

    \I__9851\ : Odrv4
    port map (
            O => \N__42414\,
            I => \c0.data_out_5_3\
        );

    \I__9850\ : InMux
    port map (
            O => \N__42403\,
            I => \N__42397\
        );

    \I__9849\ : InMux
    port map (
            O => \N__42402\,
            I => \N__42393\
        );

    \I__9848\ : InMux
    port map (
            O => \N__42401\,
            I => \N__42390\
        );

    \I__9847\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42387\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__42397\,
            I => \N__42384\
        );

    \I__9845\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42380\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__42393\,
            I => \N__42375\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__42390\,
            I => \N__42375\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__42387\,
            I => \N__42372\
        );

    \I__9841\ : Span4Mux_v
    port map (
            O => \N__42384\,
            I => \N__42368\
        );

    \I__9840\ : InMux
    port map (
            O => \N__42383\,
            I => \N__42365\
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__42380\,
            I => \N__42362\
        );

    \I__9838\ : Span4Mux_v
    port map (
            O => \N__42375\,
            I => \N__42357\
        );

    \I__9837\ : Span4Mux_v
    port map (
            O => \N__42372\,
            I => \N__42357\
        );

    \I__9836\ : InMux
    port map (
            O => \N__42371\,
            I => \N__42354\
        );

    \I__9835\ : Sp12to4
    port map (
            O => \N__42368\,
            I => \N__42349\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__42365\,
            I => \N__42349\
        );

    \I__9833\ : Odrv12
    port map (
            O => \N__42362\,
            I => \c0.data_out_5_4\
        );

    \I__9832\ : Odrv4
    port map (
            O => \N__42357\,
            I => \c0.data_out_5_4\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__42354\,
            I => \c0.data_out_5_4\
        );

    \I__9830\ : Odrv12
    port map (
            O => \N__42349\,
            I => \c0.data_out_5_4\
        );

    \I__9829\ : InMux
    port map (
            O => \N__42340\,
            I => \N__42337\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__42337\,
            I => \N__42334\
        );

    \I__9827\ : Odrv12
    port map (
            O => \N__42334\,
            I => \c0.n9783\
        );

    \I__9826\ : InMux
    port map (
            O => \N__42331\,
            I => \N__42328\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__42328\,
            I => \N__42323\
        );

    \I__9824\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42320\
        );

    \I__9823\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42317\
        );

    \I__9822\ : Span4Mux_h
    port map (
            O => \N__42323\,
            I => \N__42310\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__42320\,
            I => \N__42310\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__42317\,
            I => \N__42307\
        );

    \I__9819\ : InMux
    port map (
            O => \N__42316\,
            I => \N__42302\
        );

    \I__9818\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42302\
        );

    \I__9817\ : Span4Mux_v
    port map (
            O => \N__42310\,
            I => \N__42299\
        );

    \I__9816\ : Span4Mux_h
    port map (
            O => \N__42307\,
            I => \N__42296\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__42302\,
            I => data_out_frame2_10_6
        );

    \I__9814\ : Odrv4
    port map (
            O => \N__42299\,
            I => data_out_frame2_10_6
        );

    \I__9813\ : Odrv4
    port map (
            O => \N__42296\,
            I => data_out_frame2_10_6
        );

    \I__9812\ : InMux
    port map (
            O => \N__42289\,
            I => \N__42285\
        );

    \I__9811\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42281\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__42285\,
            I => \N__42278\
        );

    \I__9809\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42275\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__42281\,
            I => \N__42270\
        );

    \I__9807\ : Span4Mux_h
    port map (
            O => \N__42278\,
            I => \N__42270\
        );

    \I__9806\ : LocalMux
    port map (
            O => \N__42275\,
            I => \N__42267\
        );

    \I__9805\ : Span4Mux_h
    port map (
            O => \N__42270\,
            I => \N__42264\
        );

    \I__9804\ : Odrv4
    port map (
            O => \N__42267\,
            I => \c0.data_out_7_3\
        );

    \I__9803\ : Odrv4
    port map (
            O => \N__42264\,
            I => \c0.data_out_7_3\
        );

    \I__9802\ : InMux
    port map (
            O => \N__42259\,
            I => \N__42256\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__42256\,
            I => \c0.n8_adj_2153\
        );

    \I__9800\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42250\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__42250\,
            I => \N__42246\
        );

    \I__9798\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42243\
        );

    \I__9797\ : Odrv4
    port map (
            O => \N__42246\,
            I => \c0.n17070\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__42243\,
            I => \c0.n17070\
        );

    \I__9795\ : CascadeMux
    port map (
            O => \N__42238\,
            I => \N__42235\
        );

    \I__9794\ : InMux
    port map (
            O => \N__42235\,
            I => \N__42232\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__42232\,
            I => \N__42229\
        );

    \I__9792\ : Span4Mux_h
    port map (
            O => \N__42229\,
            I => \N__42225\
        );

    \I__9791\ : InMux
    port map (
            O => \N__42228\,
            I => \N__42222\
        );

    \I__9790\ : Odrv4
    port map (
            O => \N__42225\,
            I => \c0.n9737\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__42222\,
            I => \c0.n9737\
        );

    \I__9788\ : CascadeMux
    port map (
            O => \N__42217\,
            I => \N__42214\
        );

    \I__9787\ : InMux
    port map (
            O => \N__42214\,
            I => \N__42211\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__42211\,
            I => \N__42208\
        );

    \I__9785\ : Odrv4
    port map (
            O => \N__42208\,
            I => \c0.n12_adj_2285\
        );

    \I__9784\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42199\
        );

    \I__9783\ : InMux
    port map (
            O => \N__42204\,
            I => \N__42194\
        );

    \I__9782\ : InMux
    port map (
            O => \N__42203\,
            I => \N__42194\
        );

    \I__9781\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42191\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__42199\,
            I => \N__42188\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__42194\,
            I => \N__42185\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__42191\,
            I => \N__42180\
        );

    \I__9777\ : Span4Mux_v
    port map (
            O => \N__42188\,
            I => \N__42180\
        );

    \I__9776\ : Span4Mux_h
    port map (
            O => \N__42185\,
            I => \N__42177\
        );

    \I__9775\ : Odrv4
    port map (
            O => \N__42180\,
            I => \c0.data_out_6_3\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__42177\,
            I => \c0.data_out_6_3\
        );

    \I__9773\ : InMux
    port map (
            O => \N__42172\,
            I => \N__42166\
        );

    \I__9772\ : InMux
    port map (
            O => \N__42171\,
            I => \N__42166\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__42166\,
            I => \c0.data_out_2_3\
        );

    \I__9770\ : CascadeMux
    port map (
            O => \N__42163\,
            I => \N__42160\
        );

    \I__9769\ : InMux
    port map (
            O => \N__42160\,
            I => \N__42157\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__42157\,
            I => \N__42152\
        );

    \I__9767\ : InMux
    port map (
            O => \N__42156\,
            I => \N__42149\
        );

    \I__9766\ : CascadeMux
    port map (
            O => \N__42155\,
            I => \N__42146\
        );

    \I__9765\ : Span4Mux_v
    port map (
            O => \N__42152\,
            I => \N__42141\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__42149\,
            I => \N__42141\
        );

    \I__9763\ : InMux
    port map (
            O => \N__42146\,
            I => \N__42138\
        );

    \I__9762\ : Span4Mux_h
    port map (
            O => \N__42141\,
            I => \N__42135\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__42138\,
            I => \N__42132\
        );

    \I__9760\ : Span4Mux_v
    port map (
            O => \N__42135\,
            I => \N__42126\
        );

    \I__9759\ : Span4Mux_v
    port map (
            O => \N__42132\,
            I => \N__42126\
        );

    \I__9758\ : InMux
    port map (
            O => \N__42131\,
            I => \N__42123\
        );

    \I__9757\ : Odrv4
    port map (
            O => \N__42126\,
            I => n2652
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__42123\,
            I => n2652
        );

    \I__9755\ : InMux
    port map (
            O => \N__42118\,
            I => \N__42115\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__42115\,
            I => \c0.n5_adj_2350\
        );

    \I__9753\ : CascadeMux
    port map (
            O => \N__42112\,
            I => \c0.n17546_cascade_\
        );

    \I__9752\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42106\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__42106\,
            I => \N__42103\
        );

    \I__9750\ : Span4Mux_v
    port map (
            O => \N__42103\,
            I => \N__42100\
        );

    \I__9749\ : Span4Mux_h
    port map (
            O => \N__42100\,
            I => \N__42097\
        );

    \I__9748\ : Odrv4
    port map (
            O => \N__42097\,
            I => \c0.n17592\
        );

    \I__9747\ : CascadeMux
    port map (
            O => \N__42094\,
            I => \c0.n18059_cascade_\
        );

    \I__9746\ : InMux
    port map (
            O => \N__42091\,
            I => \N__42088\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__42088\,
            I => \N__42085\
        );

    \I__9744\ : Span4Mux_v
    port map (
            O => \N__42085\,
            I => \N__42082\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__42082\,
            I => \N__42079\
        );

    \I__9742\ : Odrv4
    port map (
            O => \N__42079\,
            I => \c0.data_out_frame2_20_7\
        );

    \I__9741\ : CascadeMux
    port map (
            O => \N__42076\,
            I => \c0.n18062_cascade_\
        );

    \I__9740\ : InMux
    port map (
            O => \N__42073\,
            I => \N__42069\
        );

    \I__9739\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42063\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__42069\,
            I => \N__42060\
        );

    \I__9737\ : InMux
    port map (
            O => \N__42068\,
            I => \N__42057\
        );

    \I__9736\ : InMux
    port map (
            O => \N__42067\,
            I => \N__42054\
        );

    \I__9735\ : InMux
    port map (
            O => \N__42066\,
            I => \N__42051\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__42063\,
            I => \N__42048\
        );

    \I__9733\ : Span4Mux_h
    port map (
            O => \N__42060\,
            I => \N__42043\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__42057\,
            I => \N__42043\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__42054\,
            I => data_out_frame2_11_4
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__42051\,
            I => data_out_frame2_11_4
        );

    \I__9729\ : Odrv12
    port map (
            O => \N__42048\,
            I => data_out_frame2_11_4
        );

    \I__9728\ : Odrv4
    port map (
            O => \N__42043\,
            I => data_out_frame2_11_4
        );

    \I__9727\ : InMux
    port map (
            O => \N__42034\,
            I => \N__42028\
        );

    \I__9726\ : InMux
    port map (
            O => \N__42033\,
            I => \N__42028\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__42028\,
            I => data_out_frame2_17_7
        );

    \I__9724\ : InMux
    port map (
            O => \N__42025\,
            I => \N__42020\
        );

    \I__9723\ : InMux
    port map (
            O => \N__42024\,
            I => \N__42015\
        );

    \I__9722\ : InMux
    port map (
            O => \N__42023\,
            I => \N__42015\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__42020\,
            I => data_out_frame2_14_0
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__42015\,
            I => data_out_frame2_14_0
        );

    \I__9719\ : CascadeMux
    port map (
            O => \N__42010\,
            I => \N__42007\
        );

    \I__9718\ : InMux
    port map (
            O => \N__42007\,
            I => \N__42004\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__42004\,
            I => \N__42001\
        );

    \I__9716\ : Span12Mux_v
    port map (
            O => \N__42001\,
            I => \N__41998\
        );

    \I__9715\ : Odrv12
    port map (
            O => \N__41998\,
            I => \c0.n9853\
        );

    \I__9714\ : CascadeMux
    port map (
            O => \N__41995\,
            I => \N__41991\
        );

    \I__9713\ : InMux
    port map (
            O => \N__41994\,
            I => \N__41988\
        );

    \I__9712\ : InMux
    port map (
            O => \N__41991\,
            I => \N__41985\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__41988\,
            I => \N__41982\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__41985\,
            I => \N__41979\
        );

    \I__9709\ : Span4Mux_v
    port map (
            O => \N__41982\,
            I => \N__41974\
        );

    \I__9708\ : Span4Mux_v
    port map (
            O => \N__41979\,
            I => \N__41974\
        );

    \I__9707\ : Odrv4
    port map (
            O => \N__41974\,
            I => \c0.n9589\
        );

    \I__9706\ : CascadeMux
    port map (
            O => \N__41971\,
            I => \c0.n9853_cascade_\
        );

    \I__9705\ : CascadeMux
    port map (
            O => \N__41968\,
            I => \N__41965\
        );

    \I__9704\ : InMux
    port map (
            O => \N__41965\,
            I => \N__41962\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__41962\,
            I => \N__41959\
        );

    \I__9702\ : Span12Mux_v
    port map (
            O => \N__41959\,
            I => \N__41953\
        );

    \I__9701\ : InMux
    port map (
            O => \N__41958\,
            I => \N__41950\
        );

    \I__9700\ : InMux
    port map (
            O => \N__41957\,
            I => \N__41945\
        );

    \I__9699\ : InMux
    port map (
            O => \N__41956\,
            I => \N__41945\
        );

    \I__9698\ : Odrv12
    port map (
            O => \N__41953\,
            I => data_out_frame2_13_0
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__41950\,
            I => data_out_frame2_13_0
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__41945\,
            I => data_out_frame2_13_0
        );

    \I__9695\ : InMux
    port map (
            O => \N__41938\,
            I => \N__41935\
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__41935\,
            I => \N__41931\
        );

    \I__9693\ : InMux
    port map (
            O => \N__41934\,
            I => \N__41928\
        );

    \I__9692\ : Span4Mux_v
    port map (
            O => \N__41931\,
            I => \N__41923\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__41928\,
            I => \N__41923\
        );

    \I__9690\ : Span4Mux_h
    port map (
            O => \N__41923\,
            I => \N__41920\
        );

    \I__9689\ : Span4Mux_v
    port map (
            O => \N__41920\,
            I => \N__41917\
        );

    \I__9688\ : Span4Mux_h
    port map (
            O => \N__41917\,
            I => \N__41914\
        );

    \I__9687\ : Odrv4
    port map (
            O => \N__41914\,
            I => \c0.n17046\
        );

    \I__9686\ : InMux
    port map (
            O => \N__41911\,
            I => \N__41908\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__41908\,
            I => \N__41905\
        );

    \I__9684\ : Span4Mux_h
    port map (
            O => \N__41905\,
            I => \N__41902\
        );

    \I__9683\ : Span4Mux_h
    port map (
            O => \N__41902\,
            I => \N__41899\
        );

    \I__9682\ : Odrv4
    port map (
            O => \N__41899\,
            I => \c0.n17581\
        );

    \I__9681\ : SRMux
    port map (
            O => \N__41896\,
            I => \N__41893\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__41893\,
            I => \N__41890\
        );

    \I__9679\ : Span4Mux_h
    port map (
            O => \N__41890\,
            I => \N__41886\
        );

    \I__9678\ : SRMux
    port map (
            O => \N__41889\,
            I => \N__41883\
        );

    \I__9677\ : Span4Mux_s0_v
    port map (
            O => \N__41886\,
            I => \N__41878\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41878\
        );

    \I__9675\ : Span4Mux_v
    port map (
            O => \N__41878\,
            I => \N__41875\
        );

    \I__9674\ : Odrv4
    port map (
            O => \N__41875\,
            I => \c0.n10259\
        );

    \I__9673\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41869\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__41869\,
            I => \N__41863\
        );

    \I__9671\ : InMux
    port map (
            O => \N__41868\,
            I => \N__41860\
        );

    \I__9670\ : InMux
    port map (
            O => \N__41867\,
            I => \N__41856\
        );

    \I__9669\ : InMux
    port map (
            O => \N__41866\,
            I => \N__41853\
        );

    \I__9668\ : Span4Mux_h
    port map (
            O => \N__41863\,
            I => \N__41850\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__41860\,
            I => \N__41847\
        );

    \I__9666\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41844\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__41856\,
            I => data_out_frame2_8_5
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__41853\,
            I => data_out_frame2_8_5
        );

    \I__9663\ : Odrv4
    port map (
            O => \N__41850\,
            I => data_out_frame2_8_5
        );

    \I__9662\ : Odrv12
    port map (
            O => \N__41847\,
            I => data_out_frame2_8_5
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__41844\,
            I => data_out_frame2_8_5
        );

    \I__9660\ : InMux
    port map (
            O => \N__41833\,
            I => \N__41828\
        );

    \I__9659\ : InMux
    port map (
            O => \N__41832\,
            I => \N__41825\
        );

    \I__9658\ : InMux
    port map (
            O => \N__41831\,
            I => \N__41822\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__41828\,
            I => \N__41819\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__41825\,
            I => \N__41816\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__41822\,
            I => \N__41812\
        );

    \I__9654\ : Span4Mux_v
    port map (
            O => \N__41819\,
            I => \N__41809\
        );

    \I__9653\ : Span4Mux_h
    port map (
            O => \N__41816\,
            I => \N__41806\
        );

    \I__9652\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41803\
        );

    \I__9651\ : Span4Mux_h
    port map (
            O => \N__41812\,
            I => \N__41800\
        );

    \I__9650\ : Span4Mux_h
    port map (
            O => \N__41809\,
            I => \N__41795\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__41806\,
            I => \N__41795\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__41803\,
            I => data_out_frame2_10_3
        );

    \I__9647\ : Odrv4
    port map (
            O => \N__41800\,
            I => data_out_frame2_10_3
        );

    \I__9646\ : Odrv4
    port map (
            O => \N__41795\,
            I => data_out_frame2_10_3
        );

    \I__9645\ : InMux
    port map (
            O => \N__41788\,
            I => \N__41785\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__41785\,
            I => \N__41782\
        );

    \I__9643\ : Span4Mux_h
    port map (
            O => \N__41782\,
            I => \N__41779\
        );

    \I__9642\ : Span4Mux_v
    port map (
            O => \N__41779\,
            I => \N__41776\
        );

    \I__9641\ : Odrv4
    port map (
            O => \N__41776\,
            I => \c0.n20_adj_2252\
        );

    \I__9640\ : InMux
    port map (
            O => \N__41773\,
            I => \N__41770\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__41770\,
            I => \c0.n17322\
        );

    \I__9638\ : CascadeMux
    port map (
            O => \N__41767\,
            I => \c0.n17323_cascade_\
        );

    \I__9637\ : CascadeMux
    port map (
            O => \N__41764\,
            I => \N__41761\
        );

    \I__9636\ : InMux
    port map (
            O => \N__41761\,
            I => \N__41758\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__41758\,
            I => \c0.n18053\
        );

    \I__9634\ : InMux
    port map (
            O => \N__41755\,
            I => \N__41749\
        );

    \I__9633\ : InMux
    port map (
            O => \N__41754\,
            I => \N__41746\
        );

    \I__9632\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41743\
        );

    \I__9631\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41740\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__41749\,
            I => \N__41737\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__41746\,
            I => \N__41734\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__41743\,
            I => \N__41730\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__41740\,
            I => \N__41727\
        );

    \I__9626\ : Span4Mux_v
    port map (
            O => \N__41737\,
            I => \N__41724\
        );

    \I__9625\ : Span4Mux_v
    port map (
            O => \N__41734\,
            I => \N__41721\
        );

    \I__9624\ : InMux
    port map (
            O => \N__41733\,
            I => \N__41718\
        );

    \I__9623\ : Span4Mux_v
    port map (
            O => \N__41730\,
            I => \N__41713\
        );

    \I__9622\ : Span4Mux_s3_v
    port map (
            O => \N__41727\,
            I => \N__41713\
        );

    \I__9621\ : Odrv4
    port map (
            O => \N__41724\,
            I => rand_data_16
        );

    \I__9620\ : Odrv4
    port map (
            O => \N__41721\,
            I => rand_data_16
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__41718\,
            I => rand_data_16
        );

    \I__9618\ : Odrv4
    port map (
            O => \N__41713\,
            I => rand_data_16
        );

    \I__9617\ : InMux
    port map (
            O => \N__41704\,
            I => \N__41700\
        );

    \I__9616\ : InMux
    port map (
            O => \N__41703\,
            I => \N__41697\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__41700\,
            I => \N__41691\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__41697\,
            I => \N__41691\
        );

    \I__9613\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41686\
        );

    \I__9612\ : Span12Mux_h
    port map (
            O => \N__41691\,
            I => \N__41683\
        );

    \I__9611\ : InMux
    port map (
            O => \N__41690\,
            I => \N__41680\
        );

    \I__9610\ : InMux
    port map (
            O => \N__41689\,
            I => \N__41677\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__41686\,
            I => data_out_frame2_9_1
        );

    \I__9608\ : Odrv12
    port map (
            O => \N__41683\,
            I => data_out_frame2_9_1
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__41680\,
            I => data_out_frame2_9_1
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__41677\,
            I => data_out_frame2_9_1
        );

    \I__9605\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41665\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__41665\,
            I => \c0.n17921\
        );

    \I__9603\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41659\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__41659\,
            I => \N__41656\
        );

    \I__9601\ : Span4Mux_h
    port map (
            O => \N__41656\,
            I => \N__41653\
        );

    \I__9600\ : Span4Mux_h
    port map (
            O => \N__41653\,
            I => \N__41650\
        );

    \I__9599\ : Odrv4
    port map (
            O => \N__41650\,
            I => \c0.n17924\
        );

    \I__9598\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41641\
        );

    \I__9597\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41641\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__41641\,
            I => data_out_frame2_18_7
        );

    \I__9595\ : CascadeMux
    port map (
            O => \N__41638\,
            I => \N__41635\
        );

    \I__9594\ : InMux
    port map (
            O => \N__41635\,
            I => \N__41632\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__41632\,
            I => \N__41629\
        );

    \I__9592\ : Span4Mux_v
    port map (
            O => \N__41629\,
            I => \N__41626\
        );

    \I__9591\ : Odrv4
    port map (
            O => \N__41626\,
            I => \c0.data_out_frame2_19_7\
        );

    \I__9590\ : CascadeMux
    port map (
            O => \N__41623\,
            I => \N__41620\
        );

    \I__9589\ : InMux
    port map (
            O => \N__41620\,
            I => \N__41617\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__41617\,
            I => \N__41614\
        );

    \I__9587\ : Odrv4
    port map (
            O => \N__41614\,
            I => \c0.n17034\
        );

    \I__9586\ : CascadeMux
    port map (
            O => \N__41611\,
            I => \c0.n17034_cascade_\
        );

    \I__9585\ : InMux
    port map (
            O => \N__41608\,
            I => \N__41605\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__41605\,
            I => \N__41602\
        );

    \I__9583\ : Span4Mux_h
    port map (
            O => \N__41602\,
            I => \N__41599\
        );

    \I__9582\ : Odrv4
    port map (
            O => \N__41599\,
            I => \c0.n9688\
        );

    \I__9581\ : InMux
    port map (
            O => \N__41596\,
            I => \N__41591\
        );

    \I__9580\ : InMux
    port map (
            O => \N__41595\,
            I => \N__41588\
        );

    \I__9579\ : InMux
    port map (
            O => \N__41594\,
            I => \N__41585\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__41591\,
            I => \N__41582\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__41588\,
            I => \N__41579\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__41585\,
            I => \N__41576\
        );

    \I__9575\ : Span4Mux_v
    port map (
            O => \N__41582\,
            I => \N__41571\
        );

    \I__9574\ : Span4Mux_v
    port map (
            O => \N__41579\,
            I => \N__41571\
        );

    \I__9573\ : Span4Mux_v
    port map (
            O => \N__41576\,
            I => \N__41566\
        );

    \I__9572\ : Span4Mux_h
    port map (
            O => \N__41571\,
            I => \N__41563\
        );

    \I__9571\ : InMux
    port map (
            O => \N__41570\,
            I => \N__41558\
        );

    \I__9570\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41558\
        );

    \I__9569\ : Odrv4
    port map (
            O => \N__41566\,
            I => data_out_frame2_12_1
        );

    \I__9568\ : Odrv4
    port map (
            O => \N__41563\,
            I => data_out_frame2_12_1
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__41558\,
            I => data_out_frame2_12_1
        );

    \I__9566\ : CascadeMux
    port map (
            O => \N__41551\,
            I => \c0.n9688_cascade_\
        );

    \I__9565\ : InMux
    port map (
            O => \N__41548\,
            I => \N__41545\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__41545\,
            I => \c0.n6_adj_2325\
        );

    \I__9563\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41539\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__41539\,
            I => \N__41536\
        );

    \I__9561\ : Span4Mux_h
    port map (
            O => \N__41536\,
            I => \N__41531\
        );

    \I__9560\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41526\
        );

    \I__9559\ : InMux
    port map (
            O => \N__41534\,
            I => \N__41526\
        );

    \I__9558\ : Odrv4
    port map (
            O => \N__41531\,
            I => data_out_frame2_11_1
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__41526\,
            I => data_out_frame2_11_1
        );

    \I__9556\ : InMux
    port map (
            O => \N__41521\,
            I => \N__41518\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__41518\,
            I => \N__41515\
        );

    \I__9554\ : Span4Mux_h
    port map (
            O => \N__41515\,
            I => \N__41510\
        );

    \I__9553\ : InMux
    port map (
            O => \N__41514\,
            I => \N__41506\
        );

    \I__9552\ : InMux
    port map (
            O => \N__41513\,
            I => \N__41503\
        );

    \I__9551\ : Span4Mux_h
    port map (
            O => \N__41510\,
            I => \N__41500\
        );

    \I__9550\ : InMux
    port map (
            O => \N__41509\,
            I => \N__41497\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__41506\,
            I => data_out_frame2_6_1
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__41503\,
            I => data_out_frame2_6_1
        );

    \I__9547\ : Odrv4
    port map (
            O => \N__41500\,
            I => data_out_frame2_6_1
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__41497\,
            I => data_out_frame2_6_1
        );

    \I__9545\ : InMux
    port map (
            O => \N__41488\,
            I => \N__41484\
        );

    \I__9544\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41481\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__41484\,
            I => \N__41476\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__41481\,
            I => \N__41476\
        );

    \I__9541\ : Sp12to4
    port map (
            O => \N__41476\,
            I => \N__41473\
        );

    \I__9540\ : Odrv12
    port map (
            O => \N__41473\,
            I => \c0.n17115\
        );

    \I__9539\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41466\
        );

    \I__9538\ : InMux
    port map (
            O => \N__41469\,
            I => \N__41461\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__41466\,
            I => \N__41458\
        );

    \I__9536\ : InMux
    port map (
            O => \N__41465\,
            I => \N__41455\
        );

    \I__9535\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41451\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__41461\,
            I => \N__41448\
        );

    \I__9533\ : Span4Mux_h
    port map (
            O => \N__41458\,
            I => \N__41445\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__41455\,
            I => \N__41441\
        );

    \I__9531\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41438\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__41451\,
            I => \N__41433\
        );

    \I__9529\ : Span12Mux_v
    port map (
            O => \N__41448\,
            I => \N__41433\
        );

    \I__9528\ : Span4Mux_v
    port map (
            O => \N__41445\,
            I => \N__41430\
        );

    \I__9527\ : InMux
    port map (
            O => \N__41444\,
            I => \N__41427\
        );

    \I__9526\ : Span4Mux_v
    port map (
            O => \N__41441\,
            I => \N__41424\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__41438\,
            I => rand_data_5
        );

    \I__9524\ : Odrv12
    port map (
            O => \N__41433\,
            I => rand_data_5
        );

    \I__9523\ : Odrv4
    port map (
            O => \N__41430\,
            I => rand_data_5
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__41427\,
            I => rand_data_5
        );

    \I__9521\ : Odrv4
    port map (
            O => \N__41424\,
            I => rand_data_5
        );

    \I__9520\ : CascadeMux
    port map (
            O => \N__41413\,
            I => \N__41410\
        );

    \I__9519\ : InMux
    port map (
            O => \N__41410\,
            I => \N__41407\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__41407\,
            I => \N__41403\
        );

    \I__9517\ : InMux
    port map (
            O => \N__41406\,
            I => \N__41400\
        );

    \I__9516\ : Span4Mux_h
    port map (
            O => \N__41403\,
            I => \N__41395\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__41400\,
            I => \N__41392\
        );

    \I__9514\ : InMux
    port map (
            O => \N__41399\,
            I => \N__41387\
        );

    \I__9513\ : InMux
    port map (
            O => \N__41398\,
            I => \N__41387\
        );

    \I__9512\ : Odrv4
    port map (
            O => \N__41395\,
            I => data_out_frame2_16_5
        );

    \I__9511\ : Odrv12
    port map (
            O => \N__41392\,
            I => data_out_frame2_16_5
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__41387\,
            I => data_out_frame2_16_5
        );

    \I__9509\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41376\
        );

    \I__9508\ : InMux
    port map (
            O => \N__41379\,
            I => \N__41373\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__41376\,
            I => \N__41370\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__41373\,
            I => \N__41367\
        );

    \I__9505\ : Span4Mux_v
    port map (
            O => \N__41370\,
            I => \N__41364\
        );

    \I__9504\ : Odrv12
    port map (
            O => \N__41367\,
            I => \c0.n17040\
        );

    \I__9503\ : Odrv4
    port map (
            O => \N__41364\,
            I => \c0.n17040\
        );

    \I__9502\ : InMux
    port map (
            O => \N__41359\,
            I => \N__41356\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__41356\,
            I => \c0.n16972\
        );

    \I__9500\ : InMux
    port map (
            O => \N__41353\,
            I => \N__41350\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__41350\,
            I => \c0.n30_adj_2295\
        );

    \I__9498\ : InMux
    port map (
            O => \N__41347\,
            I => \N__41340\
        );

    \I__9497\ : InMux
    port map (
            O => \N__41346\,
            I => \N__41337\
        );

    \I__9496\ : InMux
    port map (
            O => \N__41345\,
            I => \N__41334\
        );

    \I__9495\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41331\
        );

    \I__9494\ : InMux
    port map (
            O => \N__41343\,
            I => \N__41328\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__41340\,
            I => \N__41325\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__41337\,
            I => \N__41322\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__41334\,
            I => \N__41319\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__41331\,
            I => \N__41313\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__41328\,
            I => \N__41313\
        );

    \I__9488\ : Span4Mux_v
    port map (
            O => \N__41325\,
            I => \N__41308\
        );

    \I__9487\ : Span4Mux_v
    port map (
            O => \N__41322\,
            I => \N__41308\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__41319\,
            I => \N__41305\
        );

    \I__9485\ : InMux
    port map (
            O => \N__41318\,
            I => \N__41302\
        );

    \I__9484\ : Span4Mux_v
    port map (
            O => \N__41313\,
            I => \N__41297\
        );

    \I__9483\ : Span4Mux_h
    port map (
            O => \N__41308\,
            I => \N__41297\
        );

    \I__9482\ : Span4Mux_h
    port map (
            O => \N__41305\,
            I => \N__41294\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__41302\,
            I => data_out_frame2_7_7
        );

    \I__9480\ : Odrv4
    port map (
            O => \N__41297\,
            I => data_out_frame2_7_7
        );

    \I__9479\ : Odrv4
    port map (
            O => \N__41294\,
            I => data_out_frame2_7_7
        );

    \I__9478\ : CascadeMux
    port map (
            O => \N__41287\,
            I => \N__41284\
        );

    \I__9477\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41281\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41278\
        );

    \I__9475\ : Span4Mux_h
    port map (
            O => \N__41278\,
            I => \N__41275\
        );

    \I__9474\ : Span4Mux_h
    port map (
            O => \N__41275\,
            I => \N__41272\
        );

    \I__9473\ : Odrv4
    port map (
            O => \N__41272\,
            I => \c0.n5_adj_2351\
        );

    \I__9472\ : CascadeMux
    port map (
            O => \N__41269\,
            I => \N__41265\
        );

    \I__9471\ : InMux
    port map (
            O => \N__41268\,
            I => \N__41260\
        );

    \I__9470\ : InMux
    port map (
            O => \N__41265\,
            I => \N__41255\
        );

    \I__9469\ : InMux
    port map (
            O => \N__41264\,
            I => \N__41255\
        );

    \I__9468\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41252\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__41260\,
            I => \N__41249\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__41255\,
            I => data_out_frame2_11_3
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__41252\,
            I => data_out_frame2_11_3
        );

    \I__9464\ : Odrv4
    port map (
            O => \N__41249\,
            I => data_out_frame2_11_3
        );

    \I__9463\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41239\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__41239\,
            I => \N__41235\
        );

    \I__9461\ : InMux
    port map (
            O => \N__41238\,
            I => \N__41232\
        );

    \I__9460\ : Span4Mux_h
    port map (
            O => \N__41235\,
            I => \N__41229\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__41232\,
            I => \N__41226\
        );

    \I__9458\ : Odrv4
    port map (
            O => \N__41229\,
            I => \c0.n9695\
        );

    \I__9457\ : Odrv12
    port map (
            O => \N__41226\,
            I => \c0.n9695\
        );

    \I__9456\ : CascadeMux
    port map (
            O => \N__41221\,
            I => \c0.n9695_cascade_\
        );

    \I__9455\ : InMux
    port map (
            O => \N__41218\,
            I => \N__41214\
        );

    \I__9454\ : CascadeMux
    port map (
            O => \N__41217\,
            I => \N__41211\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__41214\,
            I => \N__41208\
        );

    \I__9452\ : InMux
    port map (
            O => \N__41211\,
            I => \N__41205\
        );

    \I__9451\ : Span4Mux_h
    port map (
            O => \N__41208\,
            I => \N__41198\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__41205\,
            I => \N__41198\
        );

    \I__9449\ : InMux
    port map (
            O => \N__41204\,
            I => \N__41195\
        );

    \I__9448\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41192\
        );

    \I__9447\ : Span4Mux_h
    port map (
            O => \N__41198\,
            I => \N__41189\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__41195\,
            I => \N__41186\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__41192\,
            I => \N__41182\
        );

    \I__9444\ : Span4Mux_v
    port map (
            O => \N__41189\,
            I => \N__41179\
        );

    \I__9443\ : Span4Mux_v
    port map (
            O => \N__41186\,
            I => \N__41176\
        );

    \I__9442\ : InMux
    port map (
            O => \N__41185\,
            I => \N__41173\
        );

    \I__9441\ : Span4Mux_s2_v
    port map (
            O => \N__41182\,
            I => \N__41170\
        );

    \I__9440\ : Odrv4
    port map (
            O => \N__41179\,
            I => rand_data_22
        );

    \I__9439\ : Odrv4
    port map (
            O => \N__41176\,
            I => rand_data_22
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__41173\,
            I => rand_data_22
        );

    \I__9437\ : Odrv4
    port map (
            O => \N__41170\,
            I => rand_data_22
        );

    \I__9436\ : InMux
    port map (
            O => \N__41161\,
            I => \N__41155\
        );

    \I__9435\ : InMux
    port map (
            O => \N__41160\,
            I => \N__41150\
        );

    \I__9434\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41150\
        );

    \I__9433\ : InMux
    port map (
            O => \N__41158\,
            I => \N__41147\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__41155\,
            I => data_out_frame2_11_7
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__41150\,
            I => data_out_frame2_11_7
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__41147\,
            I => data_out_frame2_11_7
        );

    \I__9429\ : InMux
    port map (
            O => \N__41140\,
            I => \N__41137\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__41137\,
            I => \N__41132\
        );

    \I__9427\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41128\
        );

    \I__9426\ : InMux
    port map (
            O => \N__41135\,
            I => \N__41125\
        );

    \I__9425\ : Span4Mux_h
    port map (
            O => \N__41132\,
            I => \N__41122\
        );

    \I__9424\ : InMux
    port map (
            O => \N__41131\,
            I => \N__41119\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__41128\,
            I => data_out_frame2_11_5
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__41125\,
            I => data_out_frame2_11_5
        );

    \I__9421\ : Odrv4
    port map (
            O => \N__41122\,
            I => data_out_frame2_11_5
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__41119\,
            I => data_out_frame2_11_5
        );

    \I__9419\ : InMux
    port map (
            O => \N__41110\,
            I => \N__41106\
        );

    \I__9418\ : InMux
    port map (
            O => \N__41109\,
            I => \N__41103\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__41106\,
            I => \N__41100\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__41103\,
            I => \N__41097\
        );

    \I__9415\ : Span4Mux_v
    port map (
            O => \N__41100\,
            I => \N__41094\
        );

    \I__9414\ : Span12Mux_s11_v
    port map (
            O => \N__41097\,
            I => \N__41091\
        );

    \I__9413\ : Odrv4
    port map (
            O => \N__41094\,
            I => \c0.n9919\
        );

    \I__9412\ : Odrv12
    port map (
            O => \N__41091\,
            I => \c0.n9919\
        );

    \I__9411\ : InMux
    port map (
            O => \N__41086\,
            I => \N__41083\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__41083\,
            I => \N__41080\
        );

    \I__9409\ : Span4Mux_h
    port map (
            O => \N__41080\,
            I => \N__41077\
        );

    \I__9408\ : Odrv4
    port map (
            O => \N__41077\,
            I => \c0.n9901\
        );

    \I__9407\ : InMux
    port map (
            O => \N__41074\,
            I => \N__41071\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__41071\,
            I => \c0.n10_adj_2292\
        );

    \I__9405\ : InMux
    port map (
            O => \N__41068\,
            I => \N__41064\
        );

    \I__9404\ : CascadeMux
    port map (
            O => \N__41067\,
            I => \N__41061\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__41064\,
            I => \N__41058\
        );

    \I__9402\ : InMux
    port map (
            O => \N__41061\,
            I => \N__41055\
        );

    \I__9401\ : Span4Mux_v
    port map (
            O => \N__41058\,
            I => \N__41050\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__41055\,
            I => \N__41050\
        );

    \I__9399\ : Span4Mux_v
    port map (
            O => \N__41050\,
            I => \N__41046\
        );

    \I__9398\ : InMux
    port map (
            O => \N__41049\,
            I => \N__41043\
        );

    \I__9397\ : Span4Mux_h
    port map (
            O => \N__41046\,
            I => \N__41037\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__41043\,
            I => \N__41034\
        );

    \I__9395\ : InMux
    port map (
            O => \N__41042\,
            I => \N__41031\
        );

    \I__9394\ : InMux
    port map (
            O => \N__41041\,
            I => \N__41026\
        );

    \I__9393\ : InMux
    port map (
            O => \N__41040\,
            I => \N__41026\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__41037\,
            I => data_out_frame2_7_4
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__41034\,
            I => data_out_frame2_7_4
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__41031\,
            I => data_out_frame2_7_4
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__41026\,
            I => data_out_frame2_7_4
        );

    \I__9388\ : InMux
    port map (
            O => \N__41017\,
            I => \N__41014\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__41014\,
            I => \N__41011\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__41011\,
            I => \N__41008\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__41008\,
            I => \c0.n9913\
        );

    \I__9384\ : InMux
    port map (
            O => \N__41005\,
            I => \N__41002\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__41002\,
            I => \c0.n29_adj_2296\
        );

    \I__9382\ : InMux
    port map (
            O => \N__40999\,
            I => \N__40996\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__40996\,
            I => \N__40993\
        );

    \I__9380\ : Span4Mux_v
    port map (
            O => \N__40993\,
            I => \N__40990\
        );

    \I__9379\ : Odrv4
    port map (
            O => \N__40990\,
            I => \c0.n16933\
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__40987\,
            I => \c0.n16915_cascade_\
        );

    \I__9377\ : InMux
    port map (
            O => \N__40984\,
            I => \N__40980\
        );

    \I__9376\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40974\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__40980\,
            I => \N__40971\
        );

    \I__9374\ : InMux
    port map (
            O => \N__40979\,
            I => \N__40968\
        );

    \I__9373\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40965\
        );

    \I__9372\ : InMux
    port map (
            O => \N__40977\,
            I => \N__40962\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__40974\,
            I => \N__40957\
        );

    \I__9370\ : Span4Mux_h
    port map (
            O => \N__40971\,
            I => \N__40957\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__40968\,
            I => \N__40954\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__40965\,
            I => \N__40949\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__40962\,
            I => \N__40949\
        );

    \I__9366\ : Odrv4
    port map (
            O => \N__40957\,
            I => data_out_frame2_7_2
        );

    \I__9365\ : Odrv4
    port map (
            O => \N__40954\,
            I => data_out_frame2_7_2
        );

    \I__9364\ : Odrv12
    port map (
            O => \N__40949\,
            I => data_out_frame2_7_2
        );

    \I__9363\ : InMux
    port map (
            O => \N__40942\,
            I => \N__40939\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__40939\,
            I => \c0.n19_adj_2303\
        );

    \I__9361\ : CascadeMux
    port map (
            O => \N__40936\,
            I => \c0.n20_adj_2302_cascade_\
        );

    \I__9360\ : InMux
    port map (
            O => \N__40933\,
            I => \N__40930\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__40930\,
            I => \N__40927\
        );

    \I__9358\ : Odrv4
    port map (
            O => \N__40927\,
            I => \c0.n21_adj_2304\
        );

    \I__9357\ : CascadeMux
    port map (
            O => \N__40924\,
            I => \N__40921\
        );

    \I__9356\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40918\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__40918\,
            I => \N__40915\
        );

    \I__9354\ : Odrv4
    port map (
            O => \N__40915\,
            I => \c0.data_out_frame2_19_6\
        );

    \I__9353\ : InMux
    port map (
            O => \N__40912\,
            I => \N__40909\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__40909\,
            I => \N__40906\
        );

    \I__9351\ : Span4Mux_v
    port map (
            O => \N__40906\,
            I => \N__40901\
        );

    \I__9350\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40895\
        );

    \I__9349\ : InMux
    port map (
            O => \N__40904\,
            I => \N__40895\
        );

    \I__9348\ : Span4Mux_h
    port map (
            O => \N__40901\,
            I => \N__40892\
        );

    \I__9347\ : InMux
    port map (
            O => \N__40900\,
            I => \N__40889\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__40895\,
            I => \N__40886\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__40892\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__40889\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9343\ : Odrv12
    port map (
            O => \N__40886\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9342\ : CascadeMux
    port map (
            O => \N__40879\,
            I => \c0.n16972_cascade_\
        );

    \I__9341\ : InMux
    port map (
            O => \N__40876\,
            I => \N__40872\
        );

    \I__9340\ : InMux
    port map (
            O => \N__40875\,
            I => \N__40868\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__40872\,
            I => \N__40865\
        );

    \I__9338\ : InMux
    port map (
            O => \N__40871\,
            I => \N__40862\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__40868\,
            I => \N__40857\
        );

    \I__9336\ : Span4Mux_h
    port map (
            O => \N__40865\,
            I => \N__40852\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__40862\,
            I => \N__40852\
        );

    \I__9334\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40849\
        );

    \I__9333\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40846\
        );

    \I__9332\ : Span12Mux_v
    port map (
            O => \N__40857\,
            I => \N__40843\
        );

    \I__9331\ : Span4Mux_h
    port map (
            O => \N__40852\,
            I => \N__40840\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__40849\,
            I => \N__40835\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__40846\,
            I => \N__40835\
        );

    \I__9328\ : Odrv12
    port map (
            O => \N__40843\,
            I => data_out_frame2_11_2
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__40840\,
            I => data_out_frame2_11_2
        );

    \I__9326\ : Odrv12
    port map (
            O => \N__40835\,
            I => data_out_frame2_11_2
        );

    \I__9325\ : InMux
    port map (
            O => \N__40828\,
            I => \N__40825\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__40825\,
            I => \N__40822\
        );

    \I__9323\ : Span4Mux_v
    port map (
            O => \N__40822\,
            I => \N__40819\
        );

    \I__9322\ : Span4Mux_h
    port map (
            O => \N__40819\,
            I => \N__40816\
        );

    \I__9321\ : Odrv4
    port map (
            O => \N__40816\,
            I => \c0.n10_adj_2281\
        );

    \I__9320\ : InMux
    port map (
            O => \N__40813\,
            I => \N__40810\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__40810\,
            I => \N__40807\
        );

    \I__9318\ : Odrv12
    port map (
            O => \N__40807\,
            I => \c0.n17969\
        );

    \I__9317\ : InMux
    port map (
            O => \N__40804\,
            I => \N__40800\
        );

    \I__9316\ : InMux
    port map (
            O => \N__40803\,
            I => \N__40796\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__40800\,
            I => \N__40793\
        );

    \I__9314\ : InMux
    port map (
            O => \N__40799\,
            I => \N__40790\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__40796\,
            I => \N__40783\
        );

    \I__9312\ : Span4Mux_v
    port map (
            O => \N__40793\,
            I => \N__40783\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__40790\,
            I => \N__40783\
        );

    \I__9310\ : Span4Mux_h
    port map (
            O => \N__40783\,
            I => \N__40778\
        );

    \I__9309\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40775\
        );

    \I__9308\ : InMux
    port map (
            O => \N__40781\,
            I => \N__40771\
        );

    \I__9307\ : Span4Mux_v
    port map (
            O => \N__40778\,
            I => \N__40768\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__40775\,
            I => \N__40765\
        );

    \I__9305\ : InMux
    port map (
            O => \N__40774\,
            I => \N__40762\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__40771\,
            I => data_out_frame2_16_4
        );

    \I__9303\ : Odrv4
    port map (
            O => \N__40768\,
            I => data_out_frame2_16_4
        );

    \I__9302\ : Odrv4
    port map (
            O => \N__40765\,
            I => data_out_frame2_16_4
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__40762\,
            I => data_out_frame2_16_4
        );

    \I__9300\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40750\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__40750\,
            I => \c0.data_out_frame2_20_4\
        );

    \I__9298\ : CascadeMux
    port map (
            O => \N__40747\,
            I => \c0.n17972_cascade_\
        );

    \I__9297\ : CascadeMux
    port map (
            O => \N__40744\,
            I => \N__40741\
        );

    \I__9296\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40738\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__40738\,
            I => \N__40735\
        );

    \I__9294\ : Span4Mux_h
    port map (
            O => \N__40735\,
            I => \N__40732\
        );

    \I__9293\ : Odrv4
    port map (
            O => \N__40732\,
            I => \c0.n17576\
        );

    \I__9292\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40726\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__40726\,
            I => \N__40721\
        );

    \I__9290\ : InMux
    port map (
            O => \N__40725\,
            I => \N__40718\
        );

    \I__9289\ : InMux
    port map (
            O => \N__40724\,
            I => \N__40714\
        );

    \I__9288\ : Span4Mux_h
    port map (
            O => \N__40721\,
            I => \N__40711\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__40718\,
            I => \N__40708\
        );

    \I__9286\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40705\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__40714\,
            I => data_out_frame2_8_3
        );

    \I__9284\ : Odrv4
    port map (
            O => \N__40711\,
            I => data_out_frame2_8_3
        );

    \I__9283\ : Odrv4
    port map (
            O => \N__40708\,
            I => data_out_frame2_8_3
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__40705\,
            I => data_out_frame2_8_3
        );

    \I__9281\ : CascadeMux
    port map (
            O => \N__40696\,
            I => \N__40693\
        );

    \I__9280\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40689\
        );

    \I__9279\ : CascadeMux
    port map (
            O => \N__40692\,
            I => \N__40686\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__40689\,
            I => \N__40683\
        );

    \I__9277\ : InMux
    port map (
            O => \N__40686\,
            I => \N__40680\
        );

    \I__9276\ : Span4Mux_h
    port map (
            O => \N__40683\,
            I => \N__40677\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__40680\,
            I => \N__40674\
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__40677\,
            I => \c0.n9839\
        );

    \I__9273\ : Odrv4
    port map (
            O => \N__40674\,
            I => \c0.n9839\
        );

    \I__9272\ : InMux
    port map (
            O => \N__40669\,
            I => \N__40665\
        );

    \I__9271\ : InMux
    port map (
            O => \N__40668\,
            I => \N__40662\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__40665\,
            I => \N__40659\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__40662\,
            I => data_out_frame2_18_6
        );

    \I__9268\ : Odrv4
    port map (
            O => \N__40659\,
            I => data_out_frame2_18_6
        );

    \I__9267\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40651\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__40651\,
            I => \N__40648\
        );

    \I__9265\ : Odrv4
    port map (
            O => \N__40648\,
            I => \c0.n16994\
        );

    \I__9264\ : InMux
    port map (
            O => \N__40645\,
            I => \N__40642\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__40642\,
            I => \N__40638\
        );

    \I__9262\ : InMux
    port map (
            O => \N__40641\,
            I => \N__40635\
        );

    \I__9261\ : Span4Mux_v
    port map (
            O => \N__40638\,
            I => \N__40631\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__40635\,
            I => \N__40628\
        );

    \I__9259\ : InMux
    port map (
            O => \N__40634\,
            I => \N__40625\
        );

    \I__9258\ : Span4Mux_h
    port map (
            O => \N__40631\,
            I => \N__40620\
        );

    \I__9257\ : Span4Mux_h
    port map (
            O => \N__40628\,
            I => \N__40620\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__40625\,
            I => \N__40615\
        );

    \I__9255\ : Span4Mux_v
    port map (
            O => \N__40620\,
            I => \N__40612\
        );

    \I__9254\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40609\
        );

    \I__9253\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40606\
        );

    \I__9252\ : Span4Mux_s2_v
    port map (
            O => \N__40615\,
            I => \N__40603\
        );

    \I__9251\ : Odrv4
    port map (
            O => \N__40612\,
            I => rand_data_21
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__40609\,
            I => rand_data_21
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__40606\,
            I => rand_data_21
        );

    \I__9248\ : Odrv4
    port map (
            O => \N__40603\,
            I => rand_data_21
        );

    \I__9247\ : InMux
    port map (
            O => \N__40594\,
            I => \N__40591\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__40591\,
            I => \N__40588\
        );

    \I__9245\ : Span4Mux_v
    port map (
            O => \N__40588\,
            I => \N__40585\
        );

    \I__9244\ : Odrv4
    port map (
            O => \N__40585\,
            I => \c0.n28_adj_2294\
        );

    \I__9243\ : CascadeMux
    port map (
            O => \N__40582\,
            I => \c0.n32_cascade_\
        );

    \I__9242\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40576\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__40576\,
            I => \c0.n31\
        );

    \I__9240\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40570\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__40570\,
            I => \N__40566\
        );

    \I__9238\ : CascadeMux
    port map (
            O => \N__40569\,
            I => \N__40563\
        );

    \I__9237\ : Span4Mux_h
    port map (
            O => \N__40566\,
            I => \N__40560\
        );

    \I__9236\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40557\
        );

    \I__9235\ : Odrv4
    port map (
            O => \N__40560\,
            I => rand_setpoint_1
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__40557\,
            I => rand_setpoint_1
        );

    \I__9233\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40547\
        );

    \I__9232\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40544\
        );

    \I__9231\ : InMux
    port map (
            O => \N__40550\,
            I => \N__40541\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__40547\,
            I => \N__40536\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__40544\,
            I => \N__40536\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__40541\,
            I => \N__40533\
        );

    \I__9227\ : Span4Mux_v
    port map (
            O => \N__40536\,
            I => \N__40530\
        );

    \I__9226\ : Odrv4
    port map (
            O => \N__40533\,
            I => \c0.data_out_7_1\
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__40530\,
            I => \c0.data_out_7_1\
        );

    \I__9224\ : CascadeMux
    port map (
            O => \N__40525\,
            I => \N__40521\
        );

    \I__9223\ : CascadeMux
    port map (
            O => \N__40524\,
            I => \N__40518\
        );

    \I__9222\ : InMux
    port map (
            O => \N__40521\,
            I => \N__40515\
        );

    \I__9221\ : InMux
    port map (
            O => \N__40518\,
            I => \N__40512\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__40515\,
            I => \N__40509\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__40512\,
            I => \N__40505\
        );

    \I__9218\ : Span4Mux_v
    port map (
            O => \N__40509\,
            I => \N__40501\
        );

    \I__9217\ : InMux
    port map (
            O => \N__40508\,
            I => \N__40498\
        );

    \I__9216\ : Span4Mux_s3_v
    port map (
            O => \N__40505\,
            I => \N__40495\
        );

    \I__9215\ : InMux
    port map (
            O => \N__40504\,
            I => \N__40492\
        );

    \I__9214\ : Span4Mux_h
    port map (
            O => \N__40501\,
            I => \N__40487\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__40498\,
            I => \N__40487\
        );

    \I__9212\ : Odrv4
    port map (
            O => \N__40495\,
            I => \c0.data_out_9_0\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__40492\,
            I => \c0.data_out_9_0\
        );

    \I__9210\ : Odrv4
    port map (
            O => \N__40487\,
            I => \c0.data_out_9_0\
        );

    \I__9209\ : InMux
    port map (
            O => \N__40480\,
            I => \N__40475\
        );

    \I__9208\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40471\
        );

    \I__9207\ : InMux
    port map (
            O => \N__40478\,
            I => \N__40468\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__40475\,
            I => \N__40465\
        );

    \I__9205\ : InMux
    port map (
            O => \N__40474\,
            I => \N__40462\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__40471\,
            I => \N__40459\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__40468\,
            I => \N__40456\
        );

    \I__9202\ : Span4Mux_v
    port map (
            O => \N__40465\,
            I => \N__40449\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__40462\,
            I => \N__40449\
        );

    \I__9200\ : Span4Mux_v
    port map (
            O => \N__40459\,
            I => \N__40444\
        );

    \I__9199\ : Span4Mux_h
    port map (
            O => \N__40456\,
            I => \N__40444\
        );

    \I__9198\ : InMux
    port map (
            O => \N__40455\,
            I => \N__40439\
        );

    \I__9197\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40439\
        );

    \I__9196\ : Span4Mux_v
    port map (
            O => \N__40449\,
            I => \N__40436\
        );

    \I__9195\ : Odrv4
    port map (
            O => \N__40444\,
            I => \c0.data_out_5_2\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__40439\,
            I => \c0.data_out_5_2\
        );

    \I__9193\ : Odrv4
    port map (
            O => \N__40436\,
            I => \c0.data_out_5_2\
        );

    \I__9192\ : CascadeMux
    port map (
            O => \N__40429\,
            I => \N__40426\
        );

    \I__9191\ : InMux
    port map (
            O => \N__40426\,
            I => \N__40420\
        );

    \I__9190\ : InMux
    port map (
            O => \N__40425\,
            I => \N__40420\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__40420\,
            I => \N__40417\
        );

    \I__9188\ : Odrv4
    port map (
            O => \N__40417\,
            I => \c0.n9522\
        );

    \I__9187\ : InMux
    port map (
            O => \N__40414\,
            I => \N__40409\
        );

    \I__9186\ : CascadeMux
    port map (
            O => \N__40413\,
            I => \N__40405\
        );

    \I__9185\ : InMux
    port map (
            O => \N__40412\,
            I => \N__40402\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__40409\,
            I => \N__40399\
        );

    \I__9183\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40396\
        );

    \I__9182\ : InMux
    port map (
            O => \N__40405\,
            I => \N__40393\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__40402\,
            I => \N__40386\
        );

    \I__9180\ : Span4Mux_v
    port map (
            O => \N__40399\,
            I => \N__40386\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__40396\,
            I => \N__40386\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__40393\,
            I => \N__40381\
        );

    \I__9177\ : Span4Mux_h
    port map (
            O => \N__40386\,
            I => \N__40378\
        );

    \I__9176\ : InMux
    port map (
            O => \N__40385\,
            I => \N__40373\
        );

    \I__9175\ : InMux
    port map (
            O => \N__40384\,
            I => \N__40373\
        );

    \I__9174\ : Odrv4
    port map (
            O => \N__40381\,
            I => data_out_8_1
        );

    \I__9173\ : Odrv4
    port map (
            O => \N__40378\,
            I => data_out_8_1
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__40373\,
            I => data_out_8_1
        );

    \I__9171\ : InMux
    port map (
            O => \N__40366\,
            I => \N__40363\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__40363\,
            I => \N__40360\
        );

    \I__9169\ : Span4Mux_s1_v
    port map (
            O => \N__40360\,
            I => \N__40357\
        );

    \I__9168\ : Span4Mux_h
    port map (
            O => \N__40357\,
            I => \N__40354\
        );

    \I__9167\ : Odrv4
    port map (
            O => \N__40354\,
            I => \c0.n18077\
        );

    \I__9166\ : InMux
    port map (
            O => \N__40351\,
            I => \N__40348\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__40348\,
            I => \N__40345\
        );

    \I__9164\ : Span4Mux_h
    port map (
            O => \N__40345\,
            I => \N__40342\
        );

    \I__9163\ : Span4Mux_v
    port map (
            O => \N__40342\,
            I => \N__40337\
        );

    \I__9162\ : InMux
    port map (
            O => \N__40341\,
            I => \N__40332\
        );

    \I__9161\ : InMux
    port map (
            O => \N__40340\,
            I => \N__40329\
        );

    \I__9160\ : Span4Mux_v
    port map (
            O => \N__40337\,
            I => \N__40326\
        );

    \I__9159\ : InMux
    port map (
            O => \N__40336\,
            I => \N__40323\
        );

    \I__9158\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40319\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__40332\,
            I => \N__40316\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__40329\,
            I => \N__40313\
        );

    \I__9155\ : Span4Mux_v
    port map (
            O => \N__40326\,
            I => \N__40308\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__40323\,
            I => \N__40308\
        );

    \I__9153\ : InMux
    port map (
            O => \N__40322\,
            I => \N__40305\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__40319\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__9151\ : Odrv4
    port map (
            O => \N__40316\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__9150\ : Odrv4
    port map (
            O => \N__40313\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__9149\ : Odrv4
    port map (
            O => \N__40308\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__40305\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__9147\ : InMux
    port map (
            O => \N__40294\,
            I => \N__40291\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__40291\,
            I => \N__40287\
        );

    \I__9145\ : CascadeMux
    port map (
            O => \N__40290\,
            I => \N__40284\
        );

    \I__9144\ : Span4Mux_h
    port map (
            O => \N__40287\,
            I => \N__40281\
        );

    \I__9143\ : InMux
    port map (
            O => \N__40284\,
            I => \N__40278\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__40281\,
            I => rand_setpoint_23
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__40278\,
            I => rand_setpoint_23
        );

    \I__9140\ : CascadeMux
    port map (
            O => \N__40273\,
            I => \c0.n17532_cascade_\
        );

    \I__9139\ : InMux
    port map (
            O => \N__40270\,
            I => \N__40266\
        );

    \I__9138\ : InMux
    port map (
            O => \N__40269\,
            I => \N__40263\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__40266\,
            I => \N__40260\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__40263\,
            I => \N__40254\
        );

    \I__9135\ : Span4Mux_s2_v
    port map (
            O => \N__40260\,
            I => \N__40254\
        );

    \I__9134\ : InMux
    port map (
            O => \N__40259\,
            I => \N__40251\
        );

    \I__9133\ : Span4Mux_h
    port map (
            O => \N__40254\,
            I => \N__40248\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__40251\,
            I => \c0.data_out_6_7\
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__40248\,
            I => \c0.data_out_6_7\
        );

    \I__9130\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40238\
        );

    \I__9129\ : InMux
    port map (
            O => \N__40242\,
            I => \N__40235\
        );

    \I__9128\ : InMux
    port map (
            O => \N__40241\,
            I => \N__40232\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__40238\,
            I => \N__40229\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__40235\,
            I => \N__40223\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__40232\,
            I => \N__40223\
        );

    \I__9124\ : Span4Mux_v
    port map (
            O => \N__40229\,
            I => \N__40220\
        );

    \I__9123\ : InMux
    port map (
            O => \N__40228\,
            I => \N__40216\
        );

    \I__9122\ : Span4Mux_s2_v
    port map (
            O => \N__40223\,
            I => \N__40211\
        );

    \I__9121\ : Span4Mux_h
    port map (
            O => \N__40220\,
            I => \N__40211\
        );

    \I__9120\ : InMux
    port map (
            O => \N__40219\,
            I => \N__40208\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__40216\,
            I => \N__40205\
        );

    \I__9118\ : Span4Mux_h
    port map (
            O => \N__40211\,
            I => \N__40202\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__40208\,
            I => \c0.data_out_5_5\
        );

    \I__9116\ : Odrv12
    port map (
            O => \N__40205\,
            I => \c0.data_out_5_5\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__40202\,
            I => \c0.data_out_5_5\
        );

    \I__9114\ : CascadeMux
    port map (
            O => \N__40195\,
            I => \N__40192\
        );

    \I__9113\ : InMux
    port map (
            O => \N__40192\,
            I => \N__40189\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__40189\,
            I => \N__40184\
        );

    \I__9111\ : CascadeMux
    port map (
            O => \N__40188\,
            I => \N__40181\
        );

    \I__9110\ : CascadeMux
    port map (
            O => \N__40187\,
            I => \N__40178\
        );

    \I__9109\ : Span4Mux_s1_v
    port map (
            O => \N__40184\,
            I => \N__40175\
        );

    \I__9108\ : InMux
    port map (
            O => \N__40181\,
            I => \N__40170\
        );

    \I__9107\ : InMux
    port map (
            O => \N__40178\,
            I => \N__40170\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__40175\,
            I => \N__40167\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__40170\,
            I => \c0.n17025\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__40167\,
            I => \c0.n17025\
        );

    \I__9103\ : InMux
    port map (
            O => \N__40162\,
            I => \N__40159\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__40159\,
            I => \N__40156\
        );

    \I__9101\ : Odrv12
    port map (
            O => \N__40156\,
            I => \c0.n17534\
        );

    \I__9100\ : InMux
    port map (
            O => \N__40153\,
            I => \N__40149\
        );

    \I__9099\ : InMux
    port map (
            O => \N__40152\,
            I => \N__40143\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__40149\,
            I => \N__40140\
        );

    \I__9097\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40137\
        );

    \I__9096\ : InMux
    port map (
            O => \N__40147\,
            I => \N__40132\
        );

    \I__9095\ : InMux
    port map (
            O => \N__40146\,
            I => \N__40132\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__40143\,
            I => \N__40129\
        );

    \I__9093\ : Span4Mux_h
    port map (
            O => \N__40140\,
            I => \N__40126\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__40137\,
            I => \N__40121\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__40132\,
            I => \N__40121\
        );

    \I__9090\ : Span4Mux_h
    port map (
            O => \N__40129\,
            I => \N__40118\
        );

    \I__9089\ : Span4Mux_v
    port map (
            O => \N__40126\,
            I => \N__40115\
        );

    \I__9088\ : Span4Mux_h
    port map (
            O => \N__40121\,
            I => \N__40112\
        );

    \I__9087\ : Odrv4
    port map (
            O => \N__40118\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__9086\ : Odrv4
    port map (
            O => \N__40115\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__9085\ : Odrv4
    port map (
            O => \N__40112\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__9084\ : InMux
    port map (
            O => \N__40105\,
            I => \N__40101\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__40104\,
            I => \N__40098\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__40101\,
            I => \N__40095\
        );

    \I__9081\ : InMux
    port map (
            O => \N__40098\,
            I => \N__40092\
        );

    \I__9080\ : Odrv4
    port map (
            O => \N__40095\,
            I => rand_setpoint_5
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__40092\,
            I => rand_setpoint_5
        );

    \I__9078\ : InMux
    port map (
            O => \N__40087\,
            I => \N__40084\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__40084\,
            I => \N__40081\
        );

    \I__9076\ : Span4Mux_v
    port map (
            O => \N__40081\,
            I => \N__40074\
        );

    \I__9075\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40067\
        );

    \I__9074\ : InMux
    port map (
            O => \N__40079\,
            I => \N__40067\
        );

    \I__9073\ : InMux
    port map (
            O => \N__40078\,
            I => \N__40067\
        );

    \I__9072\ : InMux
    port map (
            O => \N__40077\,
            I => \N__40064\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__40074\,
            I => data_out_8_5
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__40067\,
            I => data_out_8_5
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__40064\,
            I => data_out_8_5
        );

    \I__9068\ : InMux
    port map (
            O => \N__40057\,
            I => \N__40053\
        );

    \I__9067\ : InMux
    port map (
            O => \N__40056\,
            I => \N__40050\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__40053\,
            I => \c0.n28_adj_2287\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__40050\,
            I => \c0.n28_adj_2287\
        );

    \I__9064\ : InMux
    port map (
            O => \N__40045\,
            I => \N__40041\
        );

    \I__9063\ : CascadeMux
    port map (
            O => \N__40044\,
            I => \N__40038\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__40041\,
            I => \N__40035\
        );

    \I__9061\ : InMux
    port map (
            O => \N__40038\,
            I => \N__40032\
        );

    \I__9060\ : Odrv12
    port map (
            O => \N__40035\,
            I => rand_setpoint_6
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__40032\,
            I => rand_setpoint_6
        );

    \I__9058\ : InMux
    port map (
            O => \N__40027\,
            I => \N__40018\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40026\,
            I => \N__40018\
        );

    \I__9056\ : InMux
    port map (
            O => \N__40025\,
            I => \N__40013\
        );

    \I__9055\ : InMux
    port map (
            O => \N__40024\,
            I => \N__40013\
        );

    \I__9054\ : InMux
    port map (
            O => \N__40023\,
            I => \N__40010\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__40018\,
            I => \N__40005\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__40013\,
            I => \N__40005\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__40010\,
            I => data_out_8_6
        );

    \I__9050\ : Odrv4
    port map (
            O => \N__40005\,
            I => data_out_8_6
        );

    \I__9049\ : InMux
    port map (
            O => \N__40000\,
            I => \N__39997\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__39997\,
            I => \N__39994\
        );

    \I__9047\ : Span4Mux_h
    port map (
            O => \N__39994\,
            I => \N__39990\
        );

    \I__9046\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39987\
        );

    \I__9045\ : Span4Mux_h
    port map (
            O => \N__39990\,
            I => \N__39984\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__39987\,
            I => \N__39981\
        );

    \I__9043\ : Odrv4
    port map (
            O => \N__39984\,
            I => \c0.data_out_10_7\
        );

    \I__9042\ : Odrv4
    port map (
            O => \N__39981\,
            I => \c0.data_out_10_7\
        );

    \I__9041\ : InMux
    port map (
            O => \N__39976\,
            I => \N__39973\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__39973\,
            I => \c0.n8_adj_2166\
        );

    \I__9039\ : CascadeMux
    port map (
            O => \N__39970\,
            I => \N__39967\
        );

    \I__9038\ : InMux
    port map (
            O => \N__39967\,
            I => \N__39964\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__39964\,
            I => \N__39961\
        );

    \I__9036\ : Odrv12
    port map (
            O => \N__39961\,
            I => n10_adj_2425
        );

    \I__9035\ : InMux
    port map (
            O => \N__39958\,
            I => \N__39954\
        );

    \I__9034\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39951\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__39954\,
            I => \N__39948\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__39951\,
            I => \N__39945\
        );

    \I__9031\ : Span4Mux_s3_v
    port map (
            O => \N__39948\,
            I => \N__39942\
        );

    \I__9030\ : Span4Mux_v
    port map (
            O => \N__39945\,
            I => \N__39939\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__39942\,
            I => \c0.n17055\
        );

    \I__9028\ : Odrv4
    port map (
            O => \N__39939\,
            I => \c0.n17055\
        );

    \I__9027\ : InMux
    port map (
            O => \N__39934\,
            I => \N__39929\
        );

    \I__9026\ : InMux
    port map (
            O => \N__39933\,
            I => \N__39924\
        );

    \I__9025\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39924\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__39929\,
            I => \N__39919\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__39924\,
            I => \N__39919\
        );

    \I__9022\ : Odrv4
    port map (
            O => \N__39919\,
            I => \c0.data_out_9_5\
        );

    \I__9021\ : CascadeMux
    port map (
            O => \N__39916\,
            I => \N__39912\
        );

    \I__9020\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39909\
        );

    \I__9019\ : InMux
    port map (
            O => \N__39912\,
            I => \N__39906\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__39909\,
            I => \N__39903\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__39906\,
            I => \N__39900\
        );

    \I__9016\ : Span4Mux_v
    port map (
            O => \N__39903\,
            I => \N__39895\
        );

    \I__9015\ : Span4Mux_v
    port map (
            O => \N__39900\,
            I => \N__39892\
        );

    \I__9014\ : InMux
    port map (
            O => \N__39899\,
            I => \N__39887\
        );

    \I__9013\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39887\
        );

    \I__9012\ : Span4Mux_h
    port map (
            O => \N__39895\,
            I => \N__39884\
        );

    \I__9011\ : Odrv4
    port map (
            O => \N__39892\,
            I => \c0.data_out_10_1\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__39887\,
            I => \c0.data_out_10_1\
        );

    \I__9009\ : Odrv4
    port map (
            O => \N__39884\,
            I => \c0.data_out_10_1\
        );

    \I__9008\ : InMux
    port map (
            O => \N__39877\,
            I => \N__39872\
        );

    \I__9007\ : InMux
    port map (
            O => \N__39876\,
            I => \N__39868\
        );

    \I__9006\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39865\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__39872\,
            I => \N__39862\
        );

    \I__9004\ : InMux
    port map (
            O => \N__39871\,
            I => \N__39859\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__39868\,
            I => \N__39851\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__39865\,
            I => \N__39851\
        );

    \I__9001\ : Span4Mux_v
    port map (
            O => \N__39862\,
            I => \N__39851\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__39859\,
            I => \N__39848\
        );

    \I__8999\ : InMux
    port map (
            O => \N__39858\,
            I => \N__39845\
        );

    \I__8998\ : Odrv4
    port map (
            O => \N__39851\,
            I => \c0.data_out_8_2\
        );

    \I__8997\ : Odrv4
    port map (
            O => \N__39848\,
            I => \c0.data_out_8_2\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__39845\,
            I => \c0.data_out_8_2\
        );

    \I__8995\ : CascadeMux
    port map (
            O => \N__39838\,
            I => \N__39834\
        );

    \I__8994\ : InMux
    port map (
            O => \N__39837\,
            I => \N__39827\
        );

    \I__8993\ : InMux
    port map (
            O => \N__39834\,
            I => \N__39827\
        );

    \I__8992\ : InMux
    port map (
            O => \N__39833\,
            I => \N__39822\
        );

    \I__8991\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39822\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__39827\,
            I => \c0.data_out_10_5\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__39822\,
            I => \c0.data_out_10_5\
        );

    \I__8988\ : InMux
    port map (
            O => \N__39817\,
            I => \N__39814\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__39814\,
            I => \N__39809\
        );

    \I__8986\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39806\
        );

    \I__8985\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39803\
        );

    \I__8984\ : Span4Mux_s3_v
    port map (
            O => \N__39809\,
            I => \N__39800\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__39806\,
            I => \N__39795\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__39803\,
            I => \N__39795\
        );

    \I__8981\ : Span4Mux_h
    port map (
            O => \N__39800\,
            I => \N__39792\
        );

    \I__8980\ : Odrv4
    port map (
            O => \N__39795\,
            I => \c0.data_out_6_4\
        );

    \I__8979\ : Odrv4
    port map (
            O => \N__39792\,
            I => \c0.data_out_6_4\
        );

    \I__8978\ : CascadeMux
    port map (
            O => \N__39787\,
            I => \N__39783\
        );

    \I__8977\ : InMux
    port map (
            O => \N__39786\,
            I => \N__39779\
        );

    \I__8976\ : InMux
    port map (
            O => \N__39783\,
            I => \N__39776\
        );

    \I__8975\ : CascadeMux
    port map (
            O => \N__39782\,
            I => \N__39773\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__39779\,
            I => \N__39768\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__39776\,
            I => \N__39768\
        );

    \I__8972\ : InMux
    port map (
            O => \N__39773\,
            I => \N__39765\
        );

    \I__8971\ : Odrv12
    port map (
            O => \N__39768\,
            I => \c0.data_out_10_0\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__39765\,
            I => \c0.data_out_10_0\
        );

    \I__8969\ : InMux
    port map (
            O => \N__39760\,
            I => \N__39757\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__39757\,
            I => \N__39754\
        );

    \I__8967\ : Span4Mux_v
    port map (
            O => \N__39754\,
            I => \N__39751\
        );

    \I__8966\ : Span4Mux_h
    port map (
            O => \N__39751\,
            I => \N__39748\
        );

    \I__8965\ : Odrv4
    port map (
            O => \N__39748\,
            I => \c0.n16966\
        );

    \I__8964\ : CascadeMux
    port map (
            O => \N__39745\,
            I => \c0.n16966_cascade_\
        );

    \I__8963\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39739\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__39739\,
            I => \N__39736\
        );

    \I__8961\ : Odrv4
    port map (
            O => \N__39736\,
            I => \c0.n16918\
        );

    \I__8960\ : CascadeMux
    port map (
            O => \N__39733\,
            I => \c0.n10_adj_2288_cascade_\
        );

    \I__8959\ : InMux
    port map (
            O => \N__39730\,
            I => \N__39724\
        );

    \I__8958\ : InMux
    port map (
            O => \N__39729\,
            I => \N__39724\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__39724\,
            I => \c0.n17109\
        );

    \I__8956\ : InMux
    port map (
            O => \N__39721\,
            I => \N__39717\
        );

    \I__8955\ : InMux
    port map (
            O => \N__39720\,
            I => \N__39714\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__39717\,
            I => \N__39709\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__39714\,
            I => \N__39709\
        );

    \I__8952\ : Odrv12
    port map (
            O => \N__39709\,
            I => \c0.n16990\
        );

    \I__8951\ : CascadeMux
    port map (
            O => \N__39706\,
            I => \N__39701\
        );

    \I__8950\ : InMux
    port map (
            O => \N__39705\,
            I => \N__39698\
        );

    \I__8949\ : InMux
    port map (
            O => \N__39704\,
            I => \N__39695\
        );

    \I__8948\ : InMux
    port map (
            O => \N__39701\,
            I => \N__39692\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__39698\,
            I => \N__39689\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__39695\,
            I => \N__39686\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__39692\,
            I => \N__39683\
        );

    \I__8944\ : Span4Mux_h
    port map (
            O => \N__39689\,
            I => \N__39680\
        );

    \I__8943\ : Span4Mux_h
    port map (
            O => \N__39686\,
            I => \N__39675\
        );

    \I__8942\ : Span4Mux_h
    port map (
            O => \N__39683\,
            I => \N__39675\
        );

    \I__8941\ : Odrv4
    port map (
            O => \N__39680\,
            I => \c0.data_out_6_1\
        );

    \I__8940\ : Odrv4
    port map (
            O => \N__39675\,
            I => \c0.data_out_6_1\
        );

    \I__8939\ : InMux
    port map (
            O => \N__39670\,
            I => \N__39661\
        );

    \I__8938\ : InMux
    port map (
            O => \N__39669\,
            I => \N__39661\
        );

    \I__8937\ : InMux
    port map (
            O => \N__39668\,
            I => \N__39661\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__39661\,
            I => \N__39657\
        );

    \I__8935\ : InMux
    port map (
            O => \N__39660\,
            I => \N__39654\
        );

    \I__8934\ : Sp12to4
    port map (
            O => \N__39657\,
            I => \N__39651\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__39654\,
            I => data_out_frame2_7_0
        );

    \I__8932\ : Odrv12
    port map (
            O => \N__39651\,
            I => data_out_frame2_7_0
        );

    \I__8931\ : InMux
    port map (
            O => \N__39646\,
            I => \N__39643\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__39643\,
            I => \N__39640\
        );

    \I__8929\ : Odrv4
    port map (
            O => \N__39640\,
            I => \c0.n17346\
        );

    \I__8928\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39631\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__39636\,
            I => \N__39628\
        );

    \I__8926\ : InMux
    port map (
            O => \N__39635\,
            I => \N__39623\
        );

    \I__8925\ : InMux
    port map (
            O => \N__39634\,
            I => \N__39623\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__39631\,
            I => \N__39619\
        );

    \I__8923\ : InMux
    port map (
            O => \N__39628\,
            I => \N__39616\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__39623\,
            I => \N__39613\
        );

    \I__8921\ : InMux
    port map (
            O => \N__39622\,
            I => \N__39610\
        );

    \I__8920\ : Span12Mux_h
    port map (
            O => \N__39619\,
            I => \N__39605\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__39616\,
            I => \N__39605\
        );

    \I__8918\ : Odrv4
    port map (
            O => \N__39613\,
            I => rand_data_26
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__39610\,
            I => rand_data_26
        );

    \I__8916\ : Odrv12
    port map (
            O => \N__39605\,
            I => rand_data_26
        );

    \I__8915\ : InMux
    port map (
            O => \N__39598\,
            I => \N__39594\
        );

    \I__8914\ : InMux
    port map (
            O => \N__39597\,
            I => \N__39590\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__39594\,
            I => \N__39586\
        );

    \I__8912\ : InMux
    port map (
            O => \N__39593\,
            I => \N__39583\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__39590\,
            I => \N__39580\
        );

    \I__8910\ : InMux
    port map (
            O => \N__39589\,
            I => \N__39577\
        );

    \I__8909\ : Span4Mux_h
    port map (
            O => \N__39586\,
            I => \N__39573\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__39583\,
            I => \N__39568\
        );

    \I__8907\ : Span4Mux_h
    port map (
            O => \N__39580\,
            I => \N__39568\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__39577\,
            I => \N__39565\
        );

    \I__8905\ : InMux
    port map (
            O => \N__39576\,
            I => \N__39562\
        );

    \I__8904\ : Span4Mux_v
    port map (
            O => \N__39573\,
            I => \N__39559\
        );

    \I__8903\ : Span4Mux_v
    port map (
            O => \N__39568\,
            I => \N__39554\
        );

    \I__8902\ : Span4Mux_h
    port map (
            O => \N__39565\,
            I => \N__39554\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__39562\,
            I => data_out_frame2_14_2
        );

    \I__8900\ : Odrv4
    port map (
            O => \N__39559\,
            I => data_out_frame2_14_2
        );

    \I__8899\ : Odrv4
    port map (
            O => \N__39554\,
            I => data_out_frame2_14_2
        );

    \I__8898\ : CascadeMux
    port map (
            O => \N__39547\,
            I => \N__39542\
        );

    \I__8897\ : InMux
    port map (
            O => \N__39546\,
            I => \N__39539\
        );

    \I__8896\ : InMux
    port map (
            O => \N__39545\,
            I => \N__39534\
        );

    \I__8895\ : InMux
    port map (
            O => \N__39542\,
            I => \N__39534\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__39539\,
            I => \N__39529\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__39534\,
            I => \N__39526\
        );

    \I__8892\ : CascadeMux
    port map (
            O => \N__39533\,
            I => \N__39523\
        );

    \I__8891\ : InMux
    port map (
            O => \N__39532\,
            I => \N__39519\
        );

    \I__8890\ : Span4Mux_v
    port map (
            O => \N__39529\,
            I => \N__39514\
        );

    \I__8889\ : Span4Mux_v
    port map (
            O => \N__39526\,
            I => \N__39514\
        );

    \I__8888\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39511\
        );

    \I__8887\ : InMux
    port map (
            O => \N__39522\,
            I => \N__39508\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__39519\,
            I => \N__39505\
        );

    \I__8885\ : Odrv4
    port map (
            O => \N__39514\,
            I => rand_data_0
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__39511\,
            I => rand_data_0
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__39508\,
            I => rand_data_0
        );

    \I__8882\ : Odrv12
    port map (
            O => \N__39505\,
            I => rand_data_0
        );

    \I__8881\ : InMux
    port map (
            O => \N__39496\,
            I => \N__39491\
        );

    \I__8880\ : CascadeMux
    port map (
            O => \N__39495\,
            I => \N__39488\
        );

    \I__8879\ : InMux
    port map (
            O => \N__39494\,
            I => \N__39485\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__39491\,
            I => \N__39482\
        );

    \I__8877\ : InMux
    port map (
            O => \N__39488\,
            I => \N__39479\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__39485\,
            I => \N__39474\
        );

    \I__8875\ : Span4Mux_v
    port map (
            O => \N__39482\,
            I => \N__39469\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__39479\,
            I => \N__39469\
        );

    \I__8873\ : InMux
    port map (
            O => \N__39478\,
            I => \N__39464\
        );

    \I__8872\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39464\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__39474\,
            I => \N__39459\
        );

    \I__8870\ : Span4Mux_v
    port map (
            O => \N__39469\,
            I => \N__39459\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__39464\,
            I => data_out_frame2_9_0
        );

    \I__8868\ : Odrv4
    port map (
            O => \N__39459\,
            I => data_out_frame2_9_0
        );

    \I__8867\ : InMux
    port map (
            O => \N__39454\,
            I => \N__39451\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__39451\,
            I => \N__39448\
        );

    \I__8865\ : Span4Mux_h
    port map (
            O => \N__39448\,
            I => \N__39445\
        );

    \I__8864\ : Odrv4
    port map (
            O => \N__39445\,
            I => \c0.n32_adj_2297\
        );

    \I__8863\ : InMux
    port map (
            O => \N__39442\,
            I => \N__39439\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__39439\,
            I => \N__39436\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__39436\,
            I => \N__39431\
        );

    \I__8860\ : InMux
    port map (
            O => \N__39435\,
            I => \N__39428\
        );

    \I__8859\ : InMux
    port map (
            O => \N__39434\,
            I => \N__39425\
        );

    \I__8858\ : Span4Mux_v
    port map (
            O => \N__39431\,
            I => \N__39422\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__39428\,
            I => \N__39419\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__39425\,
            I => \N__39416\
        );

    \I__8855\ : Sp12to4
    port map (
            O => \N__39422\,
            I => \N__39413\
        );

    \I__8854\ : Span4Mux_h
    port map (
            O => \N__39419\,
            I => \N__39408\
        );

    \I__8853\ : Span4Mux_h
    port map (
            O => \N__39416\,
            I => \N__39408\
        );

    \I__8852\ : Odrv12
    port map (
            O => \N__39413\,
            I => \c0.n9814\
        );

    \I__8851\ : Odrv4
    port map (
            O => \N__39408\,
            I => \c0.n9814\
        );

    \I__8850\ : InMux
    port map (
            O => \N__39403\,
            I => \N__39400\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__39400\,
            I => \N__39397\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__39397\,
            I => \N__39393\
        );

    \I__8847\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39390\
        );

    \I__8846\ : Odrv4
    port map (
            O => \N__39393\,
            I => \c0.n16987\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__39390\,
            I => \c0.n16987\
        );

    \I__8844\ : InMux
    port map (
            O => \N__39385\,
            I => \N__39382\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__39382\,
            I => \N__39379\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__39379\,
            I => \c0.n25_adj_2275\
        );

    \I__8841\ : InMux
    port map (
            O => \N__39376\,
            I => \N__39369\
        );

    \I__8840\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39369\
        );

    \I__8839\ : InMux
    port map (
            O => \N__39374\,
            I => \N__39365\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__39369\,
            I => \N__39362\
        );

    \I__8837\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39359\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__39365\,
            I => \N__39355\
        );

    \I__8835\ : Span4Mux_v
    port map (
            O => \N__39362\,
            I => \N__39352\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__39359\,
            I => \N__39349\
        );

    \I__8833\ : InMux
    port map (
            O => \N__39358\,
            I => \N__39346\
        );

    \I__8832\ : Span4Mux_s3_v
    port map (
            O => \N__39355\,
            I => \N__39343\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__39352\,
            I => rand_data_17
        );

    \I__8830\ : Odrv4
    port map (
            O => \N__39349\,
            I => rand_data_17
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__39346\,
            I => rand_data_17
        );

    \I__8828\ : Odrv4
    port map (
            O => \N__39343\,
            I => rand_data_17
        );

    \I__8827\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39330\
        );

    \I__8826\ : InMux
    port map (
            O => \N__39333\,
            I => \N__39327\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__39330\,
            I => \N__39322\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__39327\,
            I => \N__39319\
        );

    \I__8823\ : InMux
    port map (
            O => \N__39326\,
            I => \N__39314\
        );

    \I__8822\ : InMux
    port map (
            O => \N__39325\,
            I => \N__39314\
        );

    \I__8821\ : Span4Mux_v
    port map (
            O => \N__39322\,
            I => \N__39311\
        );

    \I__8820\ : Odrv12
    port map (
            O => \N__39319\,
            I => data_out_frame2_6_4
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__39314\,
            I => data_out_frame2_6_4
        );

    \I__8818\ : Odrv4
    port map (
            O => \N__39311\,
            I => data_out_frame2_6_4
        );

    \I__8817\ : CascadeMux
    port map (
            O => \N__39304\,
            I => \c0.n5_adj_2141_cascade_\
        );

    \I__8816\ : InMux
    port map (
            O => \N__39301\,
            I => \N__39298\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__39298\,
            I => \N__39295\
        );

    \I__8814\ : Span4Mux_h
    port map (
            O => \N__39295\,
            I => \N__39292\
        );

    \I__8813\ : Odrv4
    port map (
            O => \N__39292\,
            I => \c0.n17987\
        );

    \I__8812\ : InMux
    port map (
            O => \N__39289\,
            I => \N__39286\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__39286\,
            I => \N__39283\
        );

    \I__8810\ : Span4Mux_h
    port map (
            O => \N__39283\,
            I => \N__39280\
        );

    \I__8809\ : Odrv4
    port map (
            O => \N__39280\,
            I => \c0.n17951\
        );

    \I__8808\ : InMux
    port map (
            O => \N__39277\,
            I => \N__39271\
        );

    \I__8807\ : InMux
    port map (
            O => \N__39276\,
            I => \N__39268\
        );

    \I__8806\ : InMux
    port map (
            O => \N__39275\,
            I => \N__39265\
        );

    \I__8805\ : InMux
    port map (
            O => \N__39274\,
            I => \N__39262\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__39271\,
            I => \N__39259\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__39268\,
            I => \N__39256\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__39265\,
            I => \N__39253\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__39262\,
            I => data_out_frame2_13_3
        );

    \I__8800\ : Odrv4
    port map (
            O => \N__39259\,
            I => data_out_frame2_13_3
        );

    \I__8799\ : Odrv4
    port map (
            O => \N__39256\,
            I => data_out_frame2_13_3
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__39253\,
            I => data_out_frame2_13_3
        );

    \I__8797\ : CascadeMux
    port map (
            O => \N__39244\,
            I => \N__39241\
        );

    \I__8796\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39238\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__39238\,
            I => \N__39235\
        );

    \I__8794\ : Span4Mux_v
    port map (
            O => \N__39235\,
            I => \N__39232\
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__39232\,
            I => \c0.n17954\
        );

    \I__8792\ : InMux
    port map (
            O => \N__39229\,
            I => \N__39226\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__39226\,
            I => \N__39223\
        );

    \I__8790\ : Span4Mux_h
    port map (
            O => \N__39223\,
            I => \N__39220\
        );

    \I__8789\ : Span4Mux_v
    port map (
            O => \N__39220\,
            I => \N__39217\
        );

    \I__8788\ : Odrv4
    port map (
            O => \N__39217\,
            I => \c0.n18056\
        );

    \I__8787\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39211\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__39211\,
            I => \N__39207\
        );

    \I__8785\ : InMux
    port map (
            O => \N__39210\,
            I => \N__39204\
        );

    \I__8784\ : Span4Mux_h
    port map (
            O => \N__39207\,
            I => \N__39199\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__39204\,
            I => \N__39195\
        );

    \I__8782\ : InMux
    port map (
            O => \N__39203\,
            I => \N__39192\
        );

    \I__8781\ : InMux
    port map (
            O => \N__39202\,
            I => \N__39189\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__39199\,
            I => \N__39186\
        );

    \I__8779\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39183\
        );

    \I__8778\ : Span4Mux_v
    port map (
            O => \N__39195\,
            I => \N__39180\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__39192\,
            I => \N__39175\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__39189\,
            I => \N__39175\
        );

    \I__8775\ : Span4Mux_h
    port map (
            O => \N__39186\,
            I => \N__39172\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__39183\,
            I => rand_data_28
        );

    \I__8773\ : Odrv4
    port map (
            O => \N__39180\,
            I => rand_data_28
        );

    \I__8772\ : Odrv12
    port map (
            O => \N__39175\,
            I => rand_data_28
        );

    \I__8771\ : Odrv4
    port map (
            O => \N__39172\,
            I => rand_data_28
        );

    \I__8770\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39160\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__39160\,
            I => \N__39156\
        );

    \I__8768\ : CascadeMux
    port map (
            O => \N__39159\,
            I => \N__39153\
        );

    \I__8767\ : Span4Mux_h
    port map (
            O => \N__39156\,
            I => \N__39148\
        );

    \I__8766\ : InMux
    port map (
            O => \N__39153\,
            I => \N__39145\
        );

    \I__8765\ : InMux
    port map (
            O => \N__39152\,
            I => \N__39140\
        );

    \I__8764\ : InMux
    port map (
            O => \N__39151\,
            I => \N__39140\
        );

    \I__8763\ : Odrv4
    port map (
            O => \N__39148\,
            I => data_out_frame2_15_2
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__39145\,
            I => data_out_frame2_15_2
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__39140\,
            I => data_out_frame2_15_2
        );

    \I__8760\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39129\
        );

    \I__8759\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39123\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__39129\,
            I => \N__39120\
        );

    \I__8757\ : InMux
    port map (
            O => \N__39128\,
            I => \N__39117\
        );

    \I__8756\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39114\
        );

    \I__8755\ : InMux
    port map (
            O => \N__39126\,
            I => \N__39111\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__39123\,
            I => \N__39108\
        );

    \I__8753\ : Span4Mux_v
    port map (
            O => \N__39120\,
            I => \N__39103\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__39117\,
            I => \N__39103\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__39114\,
            I => data_out_frame2_16_1
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__39111\,
            I => data_out_frame2_16_1
        );

    \I__8749\ : Odrv12
    port map (
            O => \N__39108\,
            I => data_out_frame2_16_1
        );

    \I__8748\ : Odrv4
    port map (
            O => \N__39103\,
            I => data_out_frame2_16_1
        );

    \I__8747\ : CascadeMux
    port map (
            O => \N__39094\,
            I => \N__39091\
        );

    \I__8746\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39087\
        );

    \I__8745\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39084\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__39087\,
            I => \N__39077\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__39084\,
            I => \N__39077\
        );

    \I__8742\ : CascadeMux
    port map (
            O => \N__39083\,
            I => \N__39074\
        );

    \I__8741\ : InMux
    port map (
            O => \N__39082\,
            I => \N__39070\
        );

    \I__8740\ : Span4Mux_v
    port map (
            O => \N__39077\,
            I => \N__39067\
        );

    \I__8739\ : InMux
    port map (
            O => \N__39074\,
            I => \N__39064\
        );

    \I__8738\ : InMux
    port map (
            O => \N__39073\,
            I => \N__39061\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__39070\,
            I => \N__39058\
        );

    \I__8736\ : Odrv4
    port map (
            O => \N__39067\,
            I => rand_data_20
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__39064\,
            I => rand_data_20
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39061\,
            I => rand_data_20
        );

    \I__8733\ : Odrv12
    port map (
            O => \N__39058\,
            I => rand_data_20
        );

    \I__8732\ : InMux
    port map (
            O => \N__39049\,
            I => \N__39045\
        );

    \I__8731\ : InMux
    port map (
            O => \N__39048\,
            I => \N__39042\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__39045\,
            I => \N__39039\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__39042\,
            I => \N__39035\
        );

    \I__8728\ : Span4Mux_h
    port map (
            O => \N__39039\,
            I => \N__39032\
        );

    \I__8727\ : InMux
    port map (
            O => \N__39038\,
            I => \N__39029\
        );

    \I__8726\ : Odrv4
    port map (
            O => \N__39035\,
            I => \c0.n9749\
        );

    \I__8725\ : Odrv4
    port map (
            O => \N__39032\,
            I => \c0.n9749\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__39029\,
            I => \c0.n9749\
        );

    \I__8723\ : InMux
    port map (
            O => \N__39022\,
            I => \N__39018\
        );

    \I__8722\ : InMux
    port map (
            O => \N__39021\,
            I => \N__39015\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__39018\,
            I => \N__39010\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__39015\,
            I => \N__39007\
        );

    \I__8719\ : InMux
    port map (
            O => \N__39014\,
            I => \N__39004\
        );

    \I__8718\ : InMux
    port map (
            O => \N__39013\,
            I => \N__39001\
        );

    \I__8717\ : Span4Mux_v
    port map (
            O => \N__39010\,
            I => \N__38998\
        );

    \I__8716\ : Span4Mux_h
    port map (
            O => \N__39007\,
            I => \N__38993\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__39004\,
            I => \N__38993\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__39001\,
            I => data_out_frame2_5_1
        );

    \I__8713\ : Odrv4
    port map (
            O => \N__38998\,
            I => data_out_frame2_5_1
        );

    \I__8712\ : Odrv4
    port map (
            O => \N__38993\,
            I => data_out_frame2_5_1
        );

    \I__8711\ : CascadeMux
    port map (
            O => \N__38986\,
            I => \N__38983\
        );

    \I__8710\ : InMux
    port map (
            O => \N__38983\,
            I => \N__38980\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__38980\,
            I => \c0.n9776\
        );

    \I__8708\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38973\
        );

    \I__8707\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38970\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__38973\,
            I => \c0.n9555\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__38970\,
            I => \c0.n9555\
        );

    \I__8704\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38962\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__38962\,
            I => \N__38959\
        );

    \I__8702\ : Span4Mux_h
    port map (
            O => \N__38959\,
            I => \N__38956\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__38956\,
            I => \c0.n16946\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__38953\,
            I => \c0.n22_adj_2207_cascade_\
        );

    \I__8699\ : InMux
    port map (
            O => \N__38950\,
            I => \N__38947\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__38947\,
            I => \N__38944\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__38944\,
            I => \N__38941\
        );

    \I__8696\ : Odrv4
    port map (
            O => \N__38941\,
            I => \c0.n18_adj_2251\
        );

    \I__8695\ : CascadeMux
    port map (
            O => \N__38938\,
            I => \c0.n9892_cascade_\
        );

    \I__8694\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38932\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__38932\,
            I => \N__38929\
        );

    \I__8692\ : Odrv4
    port map (
            O => \N__38929\,
            I => \c0.n17079\
        );

    \I__8691\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38923\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__38923\,
            I => \N__38920\
        );

    \I__8689\ : Odrv4
    port map (
            O => \N__38920\,
            I => \c0.n20_adj_2202\
        );

    \I__8688\ : CascadeMux
    port map (
            O => \N__38917\,
            I => \c0.n17079_cascade_\
        );

    \I__8687\ : InMux
    port map (
            O => \N__38914\,
            I => \N__38911\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__38911\,
            I => \N__38908\
        );

    \I__8685\ : Odrv12
    port map (
            O => \N__38908\,
            I => \c0.n24\
        );

    \I__8684\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38902\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__38902\,
            I => \N__38899\
        );

    \I__8682\ : Span4Mux_h
    port map (
            O => \N__38899\,
            I => \N__38896\
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__38896\,
            I => \c0.data_out_frame2_20_5\
        );

    \I__8680\ : InMux
    port map (
            O => \N__38893\,
            I => \N__38887\
        );

    \I__8679\ : InMux
    port map (
            O => \N__38892\,
            I => \N__38884\
        );

    \I__8678\ : InMux
    port map (
            O => \N__38891\,
            I => \N__38881\
        );

    \I__8677\ : InMux
    port map (
            O => \N__38890\,
            I => \N__38878\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__38887\,
            I => \N__38873\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__38884\,
            I => \N__38873\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__38881\,
            I => data_out_frame2_10_7
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__38878\,
            I => data_out_frame2_10_7
        );

    \I__8672\ : Odrv4
    port map (
            O => \N__38873\,
            I => data_out_frame2_10_7
        );

    \I__8671\ : CascadeMux
    port map (
            O => \N__38866\,
            I => \c0.n15_adj_2320_cascade_\
        );

    \I__8670\ : InMux
    port map (
            O => \N__38863\,
            I => \N__38859\
        );

    \I__8669\ : InMux
    port map (
            O => \N__38862\,
            I => \N__38856\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__38859\,
            I => \N__38851\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__38856\,
            I => \N__38851\
        );

    \I__8666\ : Odrv4
    port map (
            O => \N__38851\,
            I => \c0.n17088\
        );

    \I__8665\ : InMux
    port map (
            O => \N__38848\,
            I => \N__38845\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__38845\,
            I => \N__38842\
        );

    \I__8663\ : Odrv12
    port map (
            O => \N__38842\,
            I => \c0.data_out_frame2_19_2\
        );

    \I__8662\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38836\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__38836\,
            I => \c0.n14_adj_2323\
        );

    \I__8660\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38829\
        );

    \I__8659\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38826\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__38829\,
            I => \c0.n17052\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__38826\,
            I => \c0.n17052\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__38821\,
            I => \N__38818\
        );

    \I__8655\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38815\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__38815\,
            I => \N__38812\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__38812\,
            I => \N__38809\
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__38809\,
            I => \c0.n17121\
        );

    \I__8651\ : InMux
    port map (
            O => \N__38806\,
            I => \N__38803\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__38803\,
            I => \N__38800\
        );

    \I__8649\ : Span4Mux_h
    port map (
            O => \N__38800\,
            I => \N__38797\
        );

    \I__8648\ : Odrv4
    port map (
            O => \N__38797\,
            I => \c0.n19_adj_2254\
        );

    \I__8647\ : CascadeMux
    port map (
            O => \N__38794\,
            I => \c0.n21_adj_2255_cascade_\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__38791\,
            I => \N__38788\
        );

    \I__8645\ : InMux
    port map (
            O => \N__38788\,
            I => \N__38785\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__38785\,
            I => \N__38782\
        );

    \I__8643\ : Odrv4
    port map (
            O => \N__38782\,
            I => \c0.data_out_frame2_20_3\
        );

    \I__8642\ : InMux
    port map (
            O => \N__38779\,
            I => \N__38776\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__38776\,
            I => \N__38770\
        );

    \I__8640\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38767\
        );

    \I__8639\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38762\
        );

    \I__8638\ : InMux
    port map (
            O => \N__38773\,
            I => \N__38762\
        );

    \I__8637\ : Span4Mux_h
    port map (
            O => \N__38770\,
            I => \N__38759\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__38767\,
            I => data_out_frame2_14_5
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__38762\,
            I => data_out_frame2_14_5
        );

    \I__8634\ : Odrv4
    port map (
            O => \N__38759\,
            I => data_out_frame2_14_5
        );

    \I__8633\ : InMux
    port map (
            O => \N__38752\,
            I => \N__38748\
        );

    \I__8632\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38745\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__38748\,
            I => \N__38742\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__38745\,
            I => \N__38739\
        );

    \I__8629\ : Odrv4
    port map (
            O => \N__38742\,
            I => \c0.n17022\
        );

    \I__8628\ : Odrv4
    port map (
            O => \N__38739\,
            I => \c0.n17022\
        );

    \I__8627\ : InMux
    port map (
            O => \N__38734\,
            I => \N__38731\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__38731\,
            I => \c0.n26_adj_2273\
        );

    \I__8625\ : CascadeMux
    port map (
            O => \N__38728\,
            I => \N__38725\
        );

    \I__8624\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38721\
        );

    \I__8623\ : CascadeMux
    port map (
            O => \N__38724\,
            I => \N__38718\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__38721\,
            I => \N__38714\
        );

    \I__8621\ : InMux
    port map (
            O => \N__38718\,
            I => \N__38711\
        );

    \I__8620\ : CascadeMux
    port map (
            O => \N__38717\,
            I => \N__38708\
        );

    \I__8619\ : Span4Mux_h
    port map (
            O => \N__38714\,
            I => \N__38704\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__38711\,
            I => \N__38701\
        );

    \I__8617\ : InMux
    port map (
            O => \N__38708\,
            I => \N__38696\
        );

    \I__8616\ : InMux
    port map (
            O => \N__38707\,
            I => \N__38696\
        );

    \I__8615\ : Span4Mux_h
    port map (
            O => \N__38704\,
            I => \N__38693\
        );

    \I__8614\ : Span4Mux_h
    port map (
            O => \N__38701\,
            I => \N__38690\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__38696\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__8612\ : Odrv4
    port map (
            O => \N__38693\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__38690\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__8610\ : InMux
    port map (
            O => \N__38683\,
            I => \N__38680\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__38680\,
            I => \N__38676\
        );

    \I__8608\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38673\
        );

    \I__8607\ : Odrv4
    port map (
            O => \N__38676\,
            I => \c0.n17103\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__38673\,
            I => \c0.n17103\
        );

    \I__8605\ : InMux
    port map (
            O => \N__38668\,
            I => \N__38665\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__38665\,
            I => \N__38661\
        );

    \I__8603\ : InMux
    port map (
            O => \N__38664\,
            I => \N__38658\
        );

    \I__8602\ : Span4Mux_v
    port map (
            O => \N__38661\,
            I => \N__38655\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__38658\,
            I => \c0.n17067\
        );

    \I__8600\ : Odrv4
    port map (
            O => \N__38655\,
            I => \c0.n17067\
        );

    \I__8599\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38647\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__38647\,
            I => \N__38644\
        );

    \I__8597\ : Odrv4
    port map (
            O => \N__38644\,
            I => \c0.n17100\
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__38641\,
            I => \N__38637\
        );

    \I__8595\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38634\
        );

    \I__8594\ : InMux
    port map (
            O => \N__38637\,
            I => \N__38631\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__38634\,
            I => rand_setpoint_27
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__38631\,
            I => rand_setpoint_27
        );

    \I__8591\ : CascadeMux
    port map (
            O => \N__38626\,
            I => \N__38622\
        );

    \I__8590\ : InMux
    port map (
            O => \N__38625\,
            I => \N__38619\
        );

    \I__8589\ : InMux
    port map (
            O => \N__38622\,
            I => \N__38616\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__38619\,
            I => rand_setpoint_28
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__38616\,
            I => rand_setpoint_28
        );

    \I__8586\ : InMux
    port map (
            O => \N__38611\,
            I => \N__38608\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__38608\,
            I => \N__38604\
        );

    \I__8584\ : InMux
    port map (
            O => \N__38607\,
            I => \N__38601\
        );

    \I__8583\ : Span4Mux_h
    port map (
            O => \N__38604\,
            I => \N__38597\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__38601\,
            I => \N__38594\
        );

    \I__8581\ : InMux
    port map (
            O => \N__38600\,
            I => \N__38591\
        );

    \I__8580\ : Span4Mux_v
    port map (
            O => \N__38597\,
            I => \N__38586\
        );

    \I__8579\ : Span4Mux_h
    port map (
            O => \N__38594\,
            I => \N__38586\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__38591\,
            I => data_out_frame2_7_1
        );

    \I__8577\ : Odrv4
    port map (
            O => \N__38586\,
            I => data_out_frame2_7_1
        );

    \I__8576\ : InMux
    port map (
            O => \N__38581\,
            I => \N__38577\
        );

    \I__8575\ : InMux
    port map (
            O => \N__38580\,
            I => \N__38574\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__38577\,
            I => \N__38571\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__38574\,
            I => \N__38564\
        );

    \I__8572\ : Span4Mux_h
    port map (
            O => \N__38571\,
            I => \N__38564\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__38570\,
            I => \N__38561\
        );

    \I__8570\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38558\
        );

    \I__8569\ : Span4Mux_v
    port map (
            O => \N__38564\,
            I => \N__38555\
        );

    \I__8568\ : InMux
    port map (
            O => \N__38561\,
            I => \N__38552\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__38558\,
            I => data_out_frame2_10_5
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__38555\,
            I => data_out_frame2_10_5
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__38552\,
            I => data_out_frame2_10_5
        );

    \I__8564\ : InMux
    port map (
            O => \N__38545\,
            I => \N__38542\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__38542\,
            I => \N__38538\
        );

    \I__8562\ : InMux
    port map (
            O => \N__38541\,
            I => \N__38535\
        );

    \I__8561\ : Span4Mux_v
    port map (
            O => \N__38538\,
            I => \N__38532\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__38535\,
            I => \N__38529\
        );

    \I__8559\ : Odrv4
    port map (
            O => \N__38532\,
            I => \c0.n9763\
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__38529\,
            I => \c0.n9763\
        );

    \I__8557\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38519\
        );

    \I__8556\ : InMux
    port map (
            O => \N__38523\,
            I => \N__38515\
        );

    \I__8555\ : InMux
    port map (
            O => \N__38522\,
            I => \N__38511\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__38519\,
            I => \N__38508\
        );

    \I__8553\ : InMux
    port map (
            O => \N__38518\,
            I => \N__38505\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__38515\,
            I => \N__38502\
        );

    \I__8551\ : InMux
    port map (
            O => \N__38514\,
            I => \N__38499\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__38511\,
            I => \N__38494\
        );

    \I__8549\ : Span4Mux_h
    port map (
            O => \N__38508\,
            I => \N__38494\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__38505\,
            I => data_out_frame2_8_2
        );

    \I__8547\ : Odrv12
    port map (
            O => \N__38502\,
            I => data_out_frame2_8_2
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__38499\,
            I => data_out_frame2_8_2
        );

    \I__8545\ : Odrv4
    port map (
            O => \N__38494\,
            I => data_out_frame2_8_2
        );

    \I__8544\ : InMux
    port map (
            O => \N__38485\,
            I => \N__38482\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__38482\,
            I => \N__38479\
        );

    \I__8542\ : Span4Mux_h
    port map (
            O => \N__38479\,
            I => \N__38476\
        );

    \I__8541\ : Span4Mux_h
    port map (
            O => \N__38476\,
            I => \N__38473\
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__38473\,
            I => \c0.n9916\
        );

    \I__8539\ : CascadeMux
    port map (
            O => \N__38470\,
            I => \N__38466\
        );

    \I__8538\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38463\
        );

    \I__8537\ : InMux
    port map (
            O => \N__38466\,
            I => \N__38459\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__38463\,
            I => \N__38456\
        );

    \I__8535\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38452\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__38459\,
            I => \N__38447\
        );

    \I__8533\ : Span4Mux_h
    port map (
            O => \N__38456\,
            I => \N__38447\
        );

    \I__8532\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38444\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__38452\,
            I => \N__38441\
        );

    \I__8530\ : Span4Mux_v
    port map (
            O => \N__38447\,
            I => \N__38436\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__38444\,
            I => \N__38431\
        );

    \I__8528\ : Span4Mux_h
    port map (
            O => \N__38441\,
            I => \N__38431\
        );

    \I__8527\ : InMux
    port map (
            O => \N__38440\,
            I => \N__38426\
        );

    \I__8526\ : InMux
    port map (
            O => \N__38439\,
            I => \N__38426\
        );

    \I__8525\ : Odrv4
    port map (
            O => \N__38436\,
            I => data_out_frame2_12_4
        );

    \I__8524\ : Odrv4
    port map (
            O => \N__38431\,
            I => data_out_frame2_12_4
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__38426\,
            I => data_out_frame2_12_4
        );

    \I__8522\ : InMux
    port map (
            O => \N__38419\,
            I => \N__38416\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__38416\,
            I => \N__38412\
        );

    \I__8520\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38409\
        );

    \I__8519\ : Odrv12
    port map (
            O => \N__38412\,
            I => \c0.n17037\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__38409\,
            I => \c0.n17037\
        );

    \I__8517\ : CascadeMux
    port map (
            O => \N__38404\,
            I => \c0.n16933_cascade_\
        );

    \I__8516\ : InMux
    port map (
            O => \N__38401\,
            I => \N__38398\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__38398\,
            I => \c0.n17_adj_2313\
        );

    \I__8514\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38392\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__38392\,
            I => \N__38389\
        );

    \I__8512\ : Odrv4
    port map (
            O => \N__38389\,
            I => \c0.n17960\
        );

    \I__8511\ : InMux
    port map (
            O => \N__38386\,
            I => \N__38383\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__38383\,
            I => \c0.n18125\
        );

    \I__8509\ : InMux
    port map (
            O => \N__38380\,
            I => \N__38376\
        );

    \I__8508\ : InMux
    port map (
            O => \N__38379\,
            I => \N__38373\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__38376\,
            I => \N__38370\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__38373\,
            I => \N__38365\
        );

    \I__8505\ : Span4Mux_s2_v
    port map (
            O => \N__38370\,
            I => \N__38365\
        );

    \I__8504\ : Odrv4
    port map (
            O => \N__38365\,
            I => data_out_2_7
        );

    \I__8503\ : CascadeMux
    port map (
            O => \N__38362\,
            I => \N__38358\
        );

    \I__8502\ : InMux
    port map (
            O => \N__38361\,
            I => \N__38355\
        );

    \I__8501\ : InMux
    port map (
            O => \N__38358\,
            I => \N__38352\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__38355\,
            I => rand_setpoint_20
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__38352\,
            I => rand_setpoint_20
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__38347\,
            I => \N__38344\
        );

    \I__8497\ : InMux
    port map (
            O => \N__38344\,
            I => \N__38341\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__38341\,
            I => \N__38338\
        );

    \I__8495\ : Span4Mux_h
    port map (
            O => \N__38338\,
            I => \N__38335\
        );

    \I__8494\ : Odrv4
    port map (
            O => \N__38335\,
            I => \c0.n17518\
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__38332\,
            I => \N__38328\
        );

    \I__8492\ : InMux
    port map (
            O => \N__38331\,
            I => \N__38325\
        );

    \I__8491\ : InMux
    port map (
            O => \N__38328\,
            I => \N__38322\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__38325\,
            I => rand_setpoint_19
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__38322\,
            I => rand_setpoint_19
        );

    \I__8488\ : CascadeMux
    port map (
            O => \N__38317\,
            I => \N__38314\
        );

    \I__8487\ : InMux
    port map (
            O => \N__38314\,
            I => \N__38311\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__38311\,
            I => \N__38308\
        );

    \I__8485\ : Span4Mux_h
    port map (
            O => \N__38308\,
            I => \N__38305\
        );

    \I__8484\ : Span4Mux_v
    port map (
            O => \N__38305\,
            I => \N__38302\
        );

    \I__8483\ : Odrv4
    port map (
            O => \N__38302\,
            I => \c0.n17514\
        );

    \I__8482\ : CascadeMux
    port map (
            O => \N__38299\,
            I => \N__38295\
        );

    \I__8481\ : InMux
    port map (
            O => \N__38298\,
            I => \N__38292\
        );

    \I__8480\ : InMux
    port map (
            O => \N__38295\,
            I => \N__38289\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__38292\,
            I => rand_setpoint_18
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__38289\,
            I => rand_setpoint_18
        );

    \I__8477\ : CascadeMux
    port map (
            O => \N__38284\,
            I => \N__38281\
        );

    \I__8476\ : InMux
    port map (
            O => \N__38281\,
            I => \N__38278\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__38278\,
            I => \N__38275\
        );

    \I__8474\ : Odrv12
    port map (
            O => \N__38275\,
            I => \c0.n17507\
        );

    \I__8473\ : CascadeMux
    port map (
            O => \N__38272\,
            I => \N__38268\
        );

    \I__8472\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38265\
        );

    \I__8471\ : InMux
    port map (
            O => \N__38268\,
            I => \N__38262\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__38265\,
            I => rand_setpoint_17
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__38262\,
            I => rand_setpoint_17
        );

    \I__8468\ : CascadeMux
    port map (
            O => \N__38257\,
            I => \c0.n17506_cascade_\
        );

    \I__8467\ : InMux
    port map (
            O => \N__38254\,
            I => \N__38250\
        );

    \I__8466\ : InMux
    port map (
            O => \N__38253\,
            I => \N__38247\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__38250\,
            I => rand_setpoint_26
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__38247\,
            I => rand_setpoint_26
        );

    \I__8463\ : CascadeMux
    port map (
            O => \N__38242\,
            I => \N__38238\
        );

    \I__8462\ : CascadeMux
    port map (
            O => \N__38241\,
            I => \N__38235\
        );

    \I__8461\ : InMux
    port map (
            O => \N__38238\,
            I => \N__38232\
        );

    \I__8460\ : InMux
    port map (
            O => \N__38235\,
            I => \N__38229\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__38232\,
            I => rand_setpoint_29
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__38229\,
            I => rand_setpoint_29
        );

    \I__8457\ : CascadeMux
    port map (
            O => \N__38224\,
            I => \N__38220\
        );

    \I__8456\ : InMux
    port map (
            O => \N__38223\,
            I => \N__38217\
        );

    \I__8455\ : InMux
    port map (
            O => \N__38220\,
            I => \N__38214\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__38217\,
            I => rand_setpoint_24
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__38214\,
            I => rand_setpoint_24
        );

    \I__8452\ : CascadeMux
    port map (
            O => \N__38209\,
            I => \N__38206\
        );

    \I__8451\ : InMux
    port map (
            O => \N__38206\,
            I => \N__38202\
        );

    \I__8450\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38199\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__38202\,
            I => rand_setpoint_7
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__38199\,
            I => rand_setpoint_7
        );

    \I__8447\ : CascadeMux
    port map (
            O => \N__38194\,
            I => \c0.n8_adj_2169_cascade_\
        );

    \I__8446\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38188\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__38188\,
            I => \N__38185\
        );

    \I__8444\ : Span4Mux_h
    port map (
            O => \N__38185\,
            I => \N__38182\
        );

    \I__8443\ : Odrv4
    port map (
            O => \N__38182\,
            I => n10_adj_2427
        );

    \I__8442\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38176\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__38176\,
            I => \c0.n9496\
        );

    \I__8440\ : CascadeMux
    port map (
            O => \N__38173\,
            I => \N__38170\
        );

    \I__8439\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38167\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__38167\,
            I => \c0.n9716\
        );

    \I__8437\ : CascadeMux
    port map (
            O => \N__38164\,
            I => \N__38160\
        );

    \I__8436\ : CascadeMux
    port map (
            O => \N__38163\,
            I => \N__38157\
        );

    \I__8435\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38154\
        );

    \I__8434\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38151\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__38154\,
            I => rand_setpoint_2
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__38151\,
            I => rand_setpoint_2
        );

    \I__8431\ : CascadeMux
    port map (
            O => \N__38146\,
            I => \N__38143\
        );

    \I__8430\ : InMux
    port map (
            O => \N__38143\,
            I => \N__38140\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__38137\
        );

    \I__8428\ : Span4Mux_v
    port map (
            O => \N__38137\,
            I => \N__38134\
        );

    \I__8427\ : Span4Mux_h
    port map (
            O => \N__38134\,
            I => \N__38131\
        );

    \I__8426\ : Odrv4
    port map (
            O => \N__38131\,
            I => \c0.n17594\
        );

    \I__8425\ : CascadeMux
    port map (
            O => \N__38128\,
            I => \N__38125\
        );

    \I__8424\ : InMux
    port map (
            O => \N__38125\,
            I => \N__38122\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__38122\,
            I => \N__38119\
        );

    \I__8422\ : Odrv12
    port map (
            O => \N__38119\,
            I => \c0.n8_adj_2176\
        );

    \I__8421\ : InMux
    port map (
            O => \N__38116\,
            I => \N__38110\
        );

    \I__8420\ : InMux
    port map (
            O => \N__38115\,
            I => \N__38110\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__38110\,
            I => \c0.data_out_1_2\
        );

    \I__8418\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38103\
        );

    \I__8417\ : InMux
    port map (
            O => \N__38106\,
            I => \N__38098\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__38103\,
            I => \N__38093\
        );

    \I__8415\ : InMux
    port map (
            O => \N__38102\,
            I => \N__38088\
        );

    \I__8414\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38088\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__38098\,
            I => \N__38085\
        );

    \I__8412\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38082\
        );

    \I__8411\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38079\
        );

    \I__8410\ : Span4Mux_v
    port map (
            O => \N__38093\,
            I => \N__38072\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__38088\,
            I => \N__38072\
        );

    \I__8408\ : Span4Mux_h
    port map (
            O => \N__38085\,
            I => \N__38072\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__38082\,
            I => data_out_9_2
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__38079\,
            I => data_out_9_2
        );

    \I__8405\ : Odrv4
    port map (
            O => \N__38072\,
            I => data_out_9_2
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__38065\,
            I => \N__38061\
        );

    \I__8403\ : CascadeMux
    port map (
            O => \N__38064\,
            I => \N__38058\
        );

    \I__8402\ : InMux
    port map (
            O => \N__38061\,
            I => \N__38053\
        );

    \I__8401\ : InMux
    port map (
            O => \N__38058\,
            I => \N__38053\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__38053\,
            I => \N__38050\
        );

    \I__8399\ : Sp12to4
    port map (
            O => \N__38050\,
            I => \N__38047\
        );

    \I__8398\ : Span12Mux_s7_v
    port map (
            O => \N__38047\,
            I => \N__38044\
        );

    \I__8397\ : Odrv12
    port map (
            O => \N__38044\,
            I => \c0.n17064\
        );

    \I__8396\ : CascadeMux
    port map (
            O => \N__38041\,
            I => \c0.n12_adj_2289_cascade_\
        );

    \I__8395\ : InMux
    port map (
            O => \N__38038\,
            I => \N__38035\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__38035\,
            I => \N__38030\
        );

    \I__8393\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38026\
        );

    \I__8392\ : InMux
    port map (
            O => \N__38033\,
            I => \N__38022\
        );

    \I__8391\ : Span4Mux_h
    port map (
            O => \N__38030\,
            I => \N__38019\
        );

    \I__8390\ : InMux
    port map (
            O => \N__38029\,
            I => \N__38016\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__38013\
        );

    \I__8388\ : InMux
    port map (
            O => \N__38025\,
            I => \N__38010\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__38022\,
            I => \N__38007\
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__38019\,
            I => \c0.data_out_7_6\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__38016\,
            I => \c0.data_out_7_6\
        );

    \I__8384\ : Odrv12
    port map (
            O => \N__38013\,
            I => \c0.data_out_7_6\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__38010\,
            I => \c0.data_out_7_6\
        );

    \I__8382\ : Odrv4
    port map (
            O => \N__38007\,
            I => \c0.data_out_7_6\
        );

    \I__8381\ : CascadeMux
    port map (
            O => \N__37996\,
            I => \c0.n9716_cascade_\
        );

    \I__8380\ : InMux
    port map (
            O => \N__37993\,
            I => \N__37990\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__37990\,
            I => \N__37986\
        );

    \I__8378\ : InMux
    port map (
            O => \N__37989\,
            I => \N__37983\
        );

    \I__8377\ : Span4Mux_v
    port map (
            O => \N__37986\,
            I => \N__37978\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37978\
        );

    \I__8375\ : Odrv4
    port map (
            O => \N__37978\,
            I => \c0.n9728\
        );

    \I__8374\ : CascadeMux
    port map (
            O => \N__37975\,
            I => \c0.n10_adj_2162_cascade_\
        );

    \I__8373\ : InMux
    port map (
            O => \N__37972\,
            I => \N__37969\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37966\
        );

    \I__8371\ : Odrv12
    port map (
            O => \N__37966\,
            I => \data_out_9__2__N_367\
        );

    \I__8370\ : CascadeMux
    port map (
            O => \N__37963\,
            I => \data_out_9__2__N_367_cascade_\
        );

    \I__8369\ : CascadeMux
    port map (
            O => \N__37960\,
            I => \c0.n6_adj_2306_cascade_\
        );

    \I__8368\ : InMux
    port map (
            O => \N__37957\,
            I => \N__37954\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__37954\,
            I => \N__37950\
        );

    \I__8366\ : InMux
    port map (
            O => \N__37953\,
            I => \N__37947\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__37950\,
            I => \N__37940\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__37947\,
            I => \N__37940\
        );

    \I__8363\ : InMux
    port map (
            O => \N__37946\,
            I => \N__37937\
        );

    \I__8362\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37933\
        );

    \I__8361\ : Span4Mux_v
    port map (
            O => \N__37940\,
            I => \N__37930\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__37937\,
            I => \N__37927\
        );

    \I__8359\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37924\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__37933\,
            I => \N__37921\
        );

    \I__8357\ : Odrv4
    port map (
            O => \N__37930\,
            I => rand_data_27
        );

    \I__8356\ : Odrv4
    port map (
            O => \N__37927\,
            I => rand_data_27
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__37924\,
            I => rand_data_27
        );

    \I__8354\ : Odrv12
    port map (
            O => \N__37921\,
            I => rand_data_27
        );

    \I__8353\ : InMux
    port map (
            O => \N__37912\,
            I => \N__37905\
        );

    \I__8352\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37905\
        );

    \I__8351\ : InMux
    port map (
            O => \N__37910\,
            I => \N__37902\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__37905\,
            I => \N__37898\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__37902\,
            I => \N__37893\
        );

    \I__8348\ : InMux
    port map (
            O => \N__37901\,
            I => \N__37890\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__37898\,
            I => \N__37887\
        );

    \I__8346\ : InMux
    port map (
            O => \N__37897\,
            I => \N__37884\
        );

    \I__8345\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37881\
        );

    \I__8344\ : Span12Mux_h
    port map (
            O => \N__37893\,
            I => \N__37876\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__37890\,
            I => \N__37876\
        );

    \I__8342\ : Odrv4
    port map (
            O => \N__37887\,
            I => rand_data_9
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__37884\,
            I => rand_data_9
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__37881\,
            I => rand_data_9
        );

    \I__8339\ : Odrv12
    port map (
            O => \N__37876\,
            I => rand_data_9
        );

    \I__8338\ : InMux
    port map (
            O => \N__37867\,
            I => \N__37864\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__37864\,
            I => \N__37860\
        );

    \I__8336\ : InMux
    port map (
            O => \N__37863\,
            I => \N__37857\
        );

    \I__8335\ : Span4Mux_v
    port map (
            O => \N__37860\,
            I => \N__37854\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__37857\,
            I => data_out_frame2_17_1
        );

    \I__8333\ : Odrv4
    port map (
            O => \N__37854\,
            I => data_out_frame2_17_1
        );

    \I__8332\ : InMux
    port map (
            O => \N__37849\,
            I => \N__37844\
        );

    \I__8331\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37839\
        );

    \I__8330\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37839\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__37844\,
            I => \N__37834\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__37839\,
            I => \N__37831\
        );

    \I__8327\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37828\
        );

    \I__8326\ : InMux
    port map (
            O => \N__37837\,
            I => \N__37825\
        );

    \I__8325\ : Span4Mux_v
    port map (
            O => \N__37834\,
            I => \N__37822\
        );

    \I__8324\ : Span12Mux_v
    port map (
            O => \N__37831\,
            I => \N__37819\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__37828\,
            I => \N__37816\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__37825\,
            I => data_out_frame2_10_4
        );

    \I__8321\ : Odrv4
    port map (
            O => \N__37822\,
            I => data_out_frame2_10_4
        );

    \I__8320\ : Odrv12
    port map (
            O => \N__37819\,
            I => data_out_frame2_10_4
        );

    \I__8319\ : Odrv4
    port map (
            O => \N__37816\,
            I => data_out_frame2_10_4
        );

    \I__8318\ : CascadeMux
    port map (
            O => \N__37807\,
            I => \N__37804\
        );

    \I__8317\ : InMux
    port map (
            O => \N__37804\,
            I => \N__37801\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__37801\,
            I => \c0.n10_adj_2191\
        );

    \I__8315\ : InMux
    port map (
            O => \N__37798\,
            I => \N__37795\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__37795\,
            I => \N__37792\
        );

    \I__8313\ : Odrv12
    port map (
            O => \N__37792\,
            I => \c0.n14\
        );

    \I__8312\ : CascadeMux
    port map (
            O => \N__37789\,
            I => \N__37786\
        );

    \I__8311\ : InMux
    port map (
            O => \N__37786\,
            I => \N__37783\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__37783\,
            I => \N__37780\
        );

    \I__8309\ : Span4Mux_h
    port map (
            O => \N__37780\,
            I => \N__37777\
        );

    \I__8308\ : Span4Mux_v
    port map (
            O => \N__37777\,
            I => \N__37774\
        );

    \I__8307\ : Odrv4
    port map (
            O => \N__37774\,
            I => \c0.n17528\
        );

    \I__8306\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37768\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__37768\,
            I => \N__37763\
        );

    \I__8304\ : InMux
    port map (
            O => \N__37767\,
            I => \N__37760\
        );

    \I__8303\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37757\
        );

    \I__8302\ : Span4Mux_h
    port map (
            O => \N__37763\,
            I => \N__37753\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__37760\,
            I => \N__37748\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__37757\,
            I => \N__37748\
        );

    \I__8299\ : InMux
    port map (
            O => \N__37756\,
            I => \N__37745\
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__37753\,
            I => data_out_frame2_15_4
        );

    \I__8297\ : Odrv4
    port map (
            O => \N__37748\,
            I => data_out_frame2_15_4
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__37745\,
            I => data_out_frame2_15_4
        );

    \I__8295\ : CascadeMux
    port map (
            O => \N__37738\,
            I => \N__37733\
        );

    \I__8294\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37728\
        );

    \I__8293\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37725\
        );

    \I__8292\ : InMux
    port map (
            O => \N__37733\,
            I => \N__37722\
        );

    \I__8291\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37719\
        );

    \I__8290\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37716\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__37728\,
            I => \N__37713\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__37725\,
            I => \N__37708\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__37722\,
            I => \N__37708\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__37719\,
            I => \N__37703\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37703\
        );

    \I__8284\ : Span4Mux_v
    port map (
            O => \N__37713\,
            I => \N__37698\
        );

    \I__8283\ : Span4Mux_h
    port map (
            O => \N__37708\,
            I => \N__37698\
        );

    \I__8282\ : Odrv12
    port map (
            O => \N__37703\,
            I => data_out_frame2_12_5
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__37698\,
            I => data_out_frame2_12_5
        );

    \I__8280\ : InMux
    port map (
            O => \N__37693\,
            I => \N__37689\
        );

    \I__8279\ : InMux
    port map (
            O => \N__37692\,
            I => \N__37686\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__37689\,
            I => \N__37683\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__37686\,
            I => \N__37680\
        );

    \I__8276\ : Span4Mux_h
    port map (
            O => \N__37683\,
            I => \N__37675\
        );

    \I__8275\ : Span4Mux_h
    port map (
            O => \N__37680\,
            I => \N__37675\
        );

    \I__8274\ : Odrv4
    port map (
            O => \N__37675\,
            I => \c0.n17049\
        );

    \I__8273\ : CascadeMux
    port map (
            O => \N__37672\,
            I => \N__37669\
        );

    \I__8272\ : InMux
    port map (
            O => \N__37669\,
            I => \N__37665\
        );

    \I__8271\ : CascadeMux
    port map (
            O => \N__37668\,
            I => \N__37661\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__37665\,
            I => \N__37658\
        );

    \I__8269\ : InMux
    port map (
            O => \N__37664\,
            I => \N__37653\
        );

    \I__8268\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37653\
        );

    \I__8267\ : Span4Mux_h
    port map (
            O => \N__37658\,
            I => \N__37648\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__37653\,
            I => \N__37645\
        );

    \I__8265\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37642\
        );

    \I__8264\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37639\
        );

    \I__8263\ : Span4Mux_v
    port map (
            O => \N__37648\,
            I => \N__37636\
        );

    \I__8262\ : Span4Mux_h
    port map (
            O => \N__37645\,
            I => \N__37631\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__37642\,
            I => \N__37631\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__37639\,
            I => data_out_frame2_5_2
        );

    \I__8259\ : Odrv4
    port map (
            O => \N__37636\,
            I => data_out_frame2_5_2
        );

    \I__8258\ : Odrv4
    port map (
            O => \N__37631\,
            I => data_out_frame2_5_2
        );

    \I__8257\ : InMux
    port map (
            O => \N__37624\,
            I => \N__37620\
        );

    \I__8256\ : InMux
    port map (
            O => \N__37623\,
            I => \N__37617\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__37620\,
            I => \N__37614\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__37617\,
            I => \N__37611\
        );

    \I__8253\ : Odrv4
    port map (
            O => \N__37614\,
            I => \c0.n9865\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__37611\,
            I => \c0.n9865\
        );

    \I__8251\ : InMux
    port map (
            O => \N__37606\,
            I => \N__37603\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__37603\,
            I => \N__37600\
        );

    \I__8249\ : Odrv4
    port map (
            O => \N__37600\,
            I => \c0.n16908\
        );

    \I__8248\ : CascadeMux
    port map (
            O => \N__37597\,
            I => \c0.n16908_cascade_\
        );

    \I__8247\ : InMux
    port map (
            O => \N__37594\,
            I => \N__37591\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__37591\,
            I => \c0.n6_adj_2286\
        );

    \I__8245\ : InMux
    port map (
            O => \N__37588\,
            I => \N__37584\
        );

    \I__8244\ : InMux
    port map (
            O => \N__37587\,
            I => \N__37581\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__37584\,
            I => \N__37574\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__37581\,
            I => \N__37574\
        );

    \I__8241\ : InMux
    port map (
            O => \N__37580\,
            I => \N__37571\
        );

    \I__8240\ : InMux
    port map (
            O => \N__37579\,
            I => \N__37568\
        );

    \I__8239\ : Span4Mux_v
    port map (
            O => \N__37574\,
            I => \N__37565\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__37571\,
            I => \N__37562\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__37568\,
            I => data_out_frame2_14_4
        );

    \I__8236\ : Odrv4
    port map (
            O => \N__37565\,
            I => data_out_frame2_14_4
        );

    \I__8235\ : Odrv12
    port map (
            O => \N__37562\,
            I => data_out_frame2_14_4
        );

    \I__8234\ : InMux
    port map (
            O => \N__37555\,
            I => \N__37549\
        );

    \I__8233\ : InMux
    port map (
            O => \N__37554\,
            I => \N__37545\
        );

    \I__8232\ : InMux
    port map (
            O => \N__37553\,
            I => \N__37542\
        );

    \I__8231\ : InMux
    port map (
            O => \N__37552\,
            I => \N__37535\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__37549\,
            I => \N__37532\
        );

    \I__8229\ : InMux
    port map (
            O => \N__37548\,
            I => \N__37529\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__37545\,
            I => \N__37524\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__37542\,
            I => \N__37524\
        );

    \I__8226\ : InMux
    port map (
            O => \N__37541\,
            I => \N__37519\
        );

    \I__8225\ : InMux
    port map (
            O => \N__37540\,
            I => \N__37519\
        );

    \I__8224\ : InMux
    port map (
            O => \N__37539\,
            I => \N__37516\
        );

    \I__8223\ : InMux
    port map (
            O => \N__37538\,
            I => \N__37513\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__37535\,
            I => \N__37508\
        );

    \I__8221\ : Span4Mux_h
    port map (
            O => \N__37532\,
            I => \N__37508\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__37529\,
            I => \N__37505\
        );

    \I__8219\ : Span4Mux_v
    port map (
            O => \N__37524\,
            I => \N__37498\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__37519\,
            I => \N__37498\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__37516\,
            I => \N__37498\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__37513\,
            I => \N__37495\
        );

    \I__8215\ : Span4Mux_h
    port map (
            O => \N__37508\,
            I => \N__37492\
        );

    \I__8214\ : Odrv12
    port map (
            O => \N__37505\,
            I => \c0.n5543\
        );

    \I__8213\ : Odrv4
    port map (
            O => \N__37498\,
            I => \c0.n5543\
        );

    \I__8212\ : Odrv4
    port map (
            O => \N__37495\,
            I => \c0.n5543\
        );

    \I__8211\ : Odrv4
    port map (
            O => \N__37492\,
            I => \c0.n5543\
        );

    \I__8210\ : CascadeMux
    port map (
            O => \N__37483\,
            I => \N__37480\
        );

    \I__8209\ : InMux
    port map (
            O => \N__37480\,
            I => \N__37473\
        );

    \I__8208\ : InMux
    port map (
            O => \N__37479\,
            I => \N__37467\
        );

    \I__8207\ : InMux
    port map (
            O => \N__37478\,
            I => \N__37467\
        );

    \I__8206\ : InMux
    port map (
            O => \N__37477\,
            I => \N__37462\
        );

    \I__8205\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37462\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__37473\,
            I => \N__37459\
        );

    \I__8203\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37456\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__37467\,
            I => \N__37444\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__37462\,
            I => \N__37444\
        );

    \I__8200\ : Span4Mux_v
    port map (
            O => \N__37459\,
            I => \N__37444\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__37456\,
            I => \N__37444\
        );

    \I__8198\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37439\
        );

    \I__8197\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37439\
        );

    \I__8196\ : InMux
    port map (
            O => \N__37453\,
            I => \N__37436\
        );

    \I__8195\ : Span4Mux_v
    port map (
            O => \N__37444\,
            I => \N__37427\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__37439\,
            I => \N__37422\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__37436\,
            I => \N__37422\
        );

    \I__8192\ : InMux
    port map (
            O => \N__37435\,
            I => \N__37417\
        );

    \I__8191\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37417\
        );

    \I__8190\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37414\
        );

    \I__8189\ : InMux
    port map (
            O => \N__37432\,
            I => \N__37409\
        );

    \I__8188\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37409\
        );

    \I__8187\ : InMux
    port map (
            O => \N__37430\,
            I => \N__37406\
        );

    \I__8186\ : Sp12to4
    port map (
            O => \N__37427\,
            I => \N__37403\
        );

    \I__8185\ : Span4Mux_h
    port map (
            O => \N__37422\,
            I => \N__37400\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__37417\,
            I => \c0.n5545\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__37414\,
            I => \c0.n5545\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__37409\,
            I => \c0.n5545\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__37406\,
            I => \c0.n5545\
        );

    \I__8180\ : Odrv12
    port map (
            O => \N__37403\,
            I => \c0.n5545\
        );

    \I__8179\ : Odrv4
    port map (
            O => \N__37400\,
            I => \c0.n5545\
        );

    \I__8178\ : InMux
    port map (
            O => \N__37387\,
            I => \N__37384\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__37384\,
            I => \N__37379\
        );

    \I__8176\ : InMux
    port map (
            O => \N__37383\,
            I => \N__37376\
        );

    \I__8175\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37373\
        );

    \I__8174\ : Span4Mux_h
    port map (
            O => \N__37379\,
            I => \N__37370\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__37376\,
            I => \N__37367\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__37373\,
            I => \N__37364\
        );

    \I__8171\ : Span4Mux_h
    port map (
            O => \N__37370\,
            I => \N__37361\
        );

    \I__8170\ : Odrv12
    port map (
            O => \N__37367\,
            I => n31
        );

    \I__8169\ : Odrv4
    port map (
            O => \N__37364\,
            I => n31
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__37361\,
            I => n31
        );

    \I__8167\ : InMux
    port map (
            O => \N__37354\,
            I => \N__37350\
        );

    \I__8166\ : CascadeMux
    port map (
            O => \N__37353\,
            I => \N__37345\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__37350\,
            I => \N__37340\
        );

    \I__8164\ : InMux
    port map (
            O => \N__37349\,
            I => \N__37337\
        );

    \I__8163\ : InMux
    port map (
            O => \N__37348\,
            I => \N__37334\
        );

    \I__8162\ : InMux
    port map (
            O => \N__37345\,
            I => \N__37329\
        );

    \I__8161\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37329\
        );

    \I__8160\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37326\
        );

    \I__8159\ : Span4Mux_v
    port map (
            O => \N__37340\,
            I => \N__37323\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__37337\,
            I => rand_data_4
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__37334\,
            I => rand_data_4
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__37329\,
            I => rand_data_4
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__37326\,
            I => rand_data_4
        );

    \I__8154\ : Odrv4
    port map (
            O => \N__37323\,
            I => rand_data_4
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__37312\,
            I => \n10197_cascade_\
        );

    \I__8152\ : InMux
    port map (
            O => \N__37309\,
            I => \N__37306\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__37306\,
            I => \N__37299\
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__37305\,
            I => \N__37296\
        );

    \I__8149\ : InMux
    port map (
            O => \N__37304\,
            I => \N__37293\
        );

    \I__8148\ : InMux
    port map (
            O => \N__37303\,
            I => \N__37290\
        );

    \I__8147\ : InMux
    port map (
            O => \N__37302\,
            I => \N__37287\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__37299\,
            I => \N__37284\
        );

    \I__8145\ : InMux
    port map (
            O => \N__37296\,
            I => \N__37281\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__37293\,
            I => \N__37276\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__37290\,
            I => \N__37276\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__37287\,
            I => data_out_frame2_9_3
        );

    \I__8141\ : Odrv4
    port map (
            O => \N__37284\,
            I => data_out_frame2_9_3
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__37281\,
            I => data_out_frame2_9_3
        );

    \I__8139\ : Odrv4
    port map (
            O => \N__37276\,
            I => data_out_frame2_9_3
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__37267\,
            I => \c0.n17085_cascade_\
        );

    \I__8137\ : InMux
    port map (
            O => \N__37264\,
            I => \N__37260\
        );

    \I__8136\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37257\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__37260\,
            I => \N__37254\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__37257\,
            I => \N__37251\
        );

    \I__8133\ : Span4Mux_h
    port map (
            O => \N__37254\,
            I => \N__37248\
        );

    \I__8132\ : Odrv12
    port map (
            O => \N__37251\,
            I => \c0.n17073\
        );

    \I__8131\ : Odrv4
    port map (
            O => \N__37248\,
            I => \c0.n17073\
        );

    \I__8130\ : InMux
    port map (
            O => \N__37243\,
            I => \N__37240\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__37240\,
            I => \N__37237\
        );

    \I__8128\ : Span4Mux_h
    port map (
            O => \N__37237\,
            I => \N__37233\
        );

    \I__8127\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37230\
        );

    \I__8126\ : Span4Mux_v
    port map (
            O => \N__37233\,
            I => \N__37227\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__37230\,
            I => data_out_frame2_18_4
        );

    \I__8124\ : Odrv4
    port map (
            O => \N__37227\,
            I => data_out_frame2_18_4
        );

    \I__8123\ : InMux
    port map (
            O => \N__37222\,
            I => \N__37219\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__37219\,
            I => \N__37216\
        );

    \I__8121\ : Odrv4
    port map (
            O => \N__37216\,
            I => \c0.data_out_frame2_19_4\
        );

    \I__8120\ : InMux
    port map (
            O => \N__37213\,
            I => \N__37210\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__37210\,
            I => \N__37207\
        );

    \I__8118\ : Span4Mux_h
    port map (
            O => \N__37207\,
            I => \N__37203\
        );

    \I__8117\ : InMux
    port map (
            O => \N__37206\,
            I => \N__37200\
        );

    \I__8116\ : Odrv4
    port map (
            O => \N__37203\,
            I => \c0.n9707\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__37200\,
            I => \c0.n9707\
        );

    \I__8114\ : InMux
    port map (
            O => \N__37195\,
            I => \N__37192\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__37192\,
            I => \N__37188\
        );

    \I__8112\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37185\
        );

    \I__8111\ : Span4Mux_v
    port map (
            O => \N__37188\,
            I => \N__37180\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__37185\,
            I => \N__37180\
        );

    \I__8109\ : Sp12to4
    port map (
            O => \N__37180\,
            I => \N__37177\
        );

    \I__8108\ : Odrv12
    port map (
            O => \N__37177\,
            I => \c0.n16963\
        );

    \I__8107\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37171\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__37171\,
            I => \c0.n9579\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__37168\,
            I => \c0.n9579_cascade_\
        );

    \I__8104\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37162\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__37162\,
            I => \N__37159\
        );

    \I__8102\ : Odrv12
    port map (
            O => \N__37159\,
            I => \c0.n10_adj_2307\
        );

    \I__8101\ : InMux
    port map (
            O => \N__37156\,
            I => \N__37153\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__37153\,
            I => \c0.n17957\
        );

    \I__8099\ : InMux
    port map (
            O => \N__37150\,
            I => \N__37144\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37149\,
            I => \N__37141\
        );

    \I__8097\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37138\
        );

    \I__8096\ : InMux
    port map (
            O => \N__37147\,
            I => \N__37135\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__37144\,
            I => data_out_frame2_6_0
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__37141\,
            I => data_out_frame2_6_0
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__37138\,
            I => data_out_frame2_6_0
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__37135\,
            I => data_out_frame2_6_0
        );

    \I__8091\ : CascadeMux
    port map (
            O => \N__37126\,
            I => \N__37123\
        );

    \I__8090\ : InMux
    port map (
            O => \N__37123\,
            I => \N__37120\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__37120\,
            I => \c0.n5_adj_2334\
        );

    \I__8088\ : InMux
    port map (
            O => \N__37117\,
            I => \N__37113\
        );

    \I__8087\ : CascadeMux
    port map (
            O => \N__37116\,
            I => \N__37110\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__37113\,
            I => \N__37106\
        );

    \I__8085\ : InMux
    port map (
            O => \N__37110\,
            I => \N__37102\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37099\
        );

    \I__8083\ : Sp12to4
    port map (
            O => \N__37106\,
            I => \N__37096\
        );

    \I__8082\ : InMux
    port map (
            O => \N__37105\,
            I => \N__37093\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__37102\,
            I => \N__37090\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__37099\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__8079\ : Odrv12
    port map (
            O => \N__37096\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__37093\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__8077\ : Odrv4
    port map (
            O => \N__37090\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__8076\ : InMux
    port map (
            O => \N__37081\,
            I => \N__37078\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__37078\,
            I => \N__37074\
        );

    \I__8074\ : CascadeMux
    port map (
            O => \N__37077\,
            I => \N__37071\
        );

    \I__8073\ : Span4Mux_h
    port map (
            O => \N__37074\,
            I => \N__37068\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37071\,
            I => \N__37065\
        );

    \I__8071\ : Odrv4
    port map (
            O => \N__37068\,
            I => \c0.n17124\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__37065\,
            I => \c0.n17124\
        );

    \I__8069\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37057\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__37057\,
            I => \c0.n14_adj_2264\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__37054\,
            I => \N__37050\
        );

    \I__8066\ : InMux
    port map (
            O => \N__37053\,
            I => \N__37047\
        );

    \I__8065\ : InMux
    port map (
            O => \N__37050\,
            I => \N__37044\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__37047\,
            I => \N__37036\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__37044\,
            I => \N__37036\
        );

    \I__8062\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37033\
        );

    \I__8061\ : InMux
    port map (
            O => \N__37042\,
            I => \N__37028\
        );

    \I__8060\ : InMux
    port map (
            O => \N__37041\,
            I => \N__37028\
        );

    \I__8059\ : Odrv4
    port map (
            O => \N__37036\,
            I => data_out_frame2_16_2
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__37033\,
            I => data_out_frame2_16_2
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__37028\,
            I => data_out_frame2_16_2
        );

    \I__8056\ : InMux
    port map (
            O => \N__37021\,
            I => \N__37018\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__37018\,
            I => \N__37015\
        );

    \I__8054\ : Span4Mux_v
    port map (
            O => \N__37015\,
            I => \N__37012\
        );

    \I__8053\ : Span4Mux_h
    port map (
            O => \N__37012\,
            I => \N__37009\
        );

    \I__8052\ : Span4Mux_h
    port map (
            O => \N__37009\,
            I => \N__37006\
        );

    \I__8051\ : Odrv4
    port map (
            O => \N__37006\,
            I => \c0.n17031\
        );

    \I__8050\ : InMux
    port map (
            O => \N__37003\,
            I => \N__37000\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__37000\,
            I => \N__36997\
        );

    \I__8048\ : Span4Mux_h
    port map (
            O => \N__36997\,
            I => \N__36994\
        );

    \I__8047\ : Odrv4
    port map (
            O => \N__36994\,
            I => \c0.n17091\
        );

    \I__8046\ : CascadeMux
    port map (
            O => \N__36991\,
            I => \c0.n17031_cascade_\
        );

    \I__8045\ : InMux
    port map (
            O => \N__36988\,
            I => \N__36984\
        );

    \I__8044\ : InMux
    port map (
            O => \N__36987\,
            I => \N__36981\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__36984\,
            I => \N__36978\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__36981\,
            I => \N__36975\
        );

    \I__8041\ : Span4Mux_h
    port map (
            O => \N__36978\,
            I => \N__36972\
        );

    \I__8040\ : Odrv4
    port map (
            O => \N__36975\,
            I => \c0.n9692\
        );

    \I__8039\ : Odrv4
    port map (
            O => \N__36972\,
            I => \c0.n9692\
        );

    \I__8038\ : InMux
    port map (
            O => \N__36967\,
            I => \N__36964\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__36964\,
            I => \c0.n17085\
        );

    \I__8036\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36958\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__36958\,
            I => \c0.n18_adj_2331\
        );

    \I__8034\ : CascadeMux
    port map (
            O => \N__36955\,
            I => \c0.n17100_cascade_\
        );

    \I__8033\ : CascadeMux
    port map (
            O => \N__36952\,
            I => \c0.n16_adj_2332_cascade_\
        );

    \I__8032\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36946\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__36946\,
            I => \c0.n20_adj_2333\
        );

    \I__8030\ : CascadeMux
    port map (
            O => \N__36943\,
            I => \N__36940\
        );

    \I__8029\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36937\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__36937\,
            I => \N__36934\
        );

    \I__8027\ : Span4Mux_h
    port map (
            O => \N__36934\,
            I => \N__36931\
        );

    \I__8026\ : Odrv4
    port map (
            O => \N__36931\,
            I => \c0.data_out_frame2_19_0\
        );

    \I__8025\ : InMux
    port map (
            O => \N__36928\,
            I => \N__36925\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__36925\,
            I => \c0.n9886\
        );

    \I__8023\ : CascadeMux
    port map (
            O => \N__36922\,
            I => \c0.n12_adj_2263_cascade_\
        );

    \I__8022\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36916\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__36916\,
            I => \N__36913\
        );

    \I__8020\ : Span4Mux_h
    port map (
            O => \N__36913\,
            I => \N__36910\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__36910\,
            I => \c0.data_out_frame2_20_2\
        );

    \I__8018\ : InMux
    port map (
            O => \N__36907\,
            I => \N__36904\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__36904\,
            I => \N__36901\
        );

    \I__8016\ : Span4Mux_v
    port map (
            O => \N__36901\,
            I => \N__36898\
        );

    \I__8015\ : Odrv4
    port map (
            O => \N__36898\,
            I => \c0.n17112\
        );

    \I__8014\ : CascadeMux
    port map (
            O => \N__36895\,
            I => \c0.n16_adj_2312_cascade_\
        );

    \I__8013\ : CascadeMux
    port map (
            O => \N__36892\,
            I => \N__36889\
        );

    \I__8012\ : InMux
    port map (
            O => \N__36889\,
            I => \N__36885\
        );

    \I__8011\ : InMux
    port map (
            O => \N__36888\,
            I => \N__36882\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__36885\,
            I => \c0.n17097\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__36882\,
            I => \c0.n17097\
        );

    \I__8008\ : InMux
    port map (
            O => \N__36877\,
            I => n15586
        );

    \I__8007\ : InMux
    port map (
            O => \N__36874\,
            I => n15587
        );

    \I__8006\ : CascadeMux
    port map (
            O => \N__36871\,
            I => \N__36867\
        );

    \I__8005\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36864\
        );

    \I__8004\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36861\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__36864\,
            I => rand_setpoint_30
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__36861\,
            I => rand_setpoint_30
        );

    \I__8001\ : InMux
    port map (
            O => \N__36856\,
            I => n15588
        );

    \I__8000\ : InMux
    port map (
            O => \N__36853\,
            I => n15589
        );

    \I__7999\ : InMux
    port map (
            O => \N__36850\,
            I => \N__36846\
        );

    \I__7998\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36843\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__36846\,
            I => rand_setpoint_31
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__36843\,
            I => rand_setpoint_31
        );

    \I__7995\ : InMux
    port map (
            O => \N__36838\,
            I => \N__36835\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__36835\,
            I => \N__36832\
        );

    \I__7993\ : Span4Mux_v
    port map (
            O => \N__36832\,
            I => \N__36829\
        );

    \I__7992\ : Span4Mux_h
    port map (
            O => \N__36829\,
            I => \N__36824\
        );

    \I__7991\ : CascadeMux
    port map (
            O => \N__36828\,
            I => \N__36821\
        );

    \I__7990\ : InMux
    port map (
            O => \N__36827\,
            I => \N__36817\
        );

    \I__7989\ : Span4Mux_v
    port map (
            O => \N__36824\,
            I => \N__36814\
        );

    \I__7988\ : InMux
    port map (
            O => \N__36821\,
            I => \N__36811\
        );

    \I__7987\ : InMux
    port map (
            O => \N__36820\,
            I => \N__36808\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__36817\,
            I => \N__36803\
        );

    \I__7985\ : Span4Mux_v
    port map (
            O => \N__36814\,
            I => \N__36803\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__36811\,
            I => \c0.data_out_7_4\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__36808\,
            I => \c0.data_out_7_4\
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__36803\,
            I => \c0.data_out_7_4\
        );

    \I__7981\ : CascadeMux
    port map (
            O => \N__36796\,
            I => \c0.n22_adj_2357_cascade_\
        );

    \I__7980\ : InMux
    port map (
            O => \N__36793\,
            I => \N__36790\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__36790\,
            I => \N__36787\
        );

    \I__7978\ : Span12Mux_v
    port map (
            O => \N__36787\,
            I => \N__36784\
        );

    \I__7977\ : Odrv12
    port map (
            O => \N__36784\,
            I => \c0.tx2.r_Tx_Data_3\
        );

    \I__7976\ : InMux
    port map (
            O => \N__36781\,
            I => \N__36778\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__36778\,
            I => \N__36775\
        );

    \I__7974\ : Span4Mux_h
    port map (
            O => \N__36775\,
            I => \N__36772\
        );

    \I__7973\ : Odrv4
    port map (
            O => \N__36772\,
            I => \c0.n6_adj_2187\
        );

    \I__7972\ : InMux
    port map (
            O => \N__36769\,
            I => \N__36766\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__36766\,
            I => \c0.n18128\
        );

    \I__7970\ : CascadeMux
    port map (
            O => \N__36763\,
            I => \N__36760\
        );

    \I__7969\ : InMux
    port map (
            O => \N__36760\,
            I => \N__36757\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__36757\,
            I => \N__36753\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__36756\,
            I => \N__36750\
        );

    \I__7966\ : Span4Mux_h
    port map (
            O => \N__36753\,
            I => \N__36747\
        );

    \I__7965\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36744\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__36747\,
            I => \N__36741\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__36744\,
            I => \c0.n16936\
        );

    \I__7962\ : Odrv4
    port map (
            O => \N__36741\,
            I => \c0.n16936\
        );

    \I__7961\ : InMux
    port map (
            O => \N__36736\,
            I => \N__36732\
        );

    \I__7960\ : CascadeMux
    port map (
            O => \N__36735\,
            I => \N__36728\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__36732\,
            I => \N__36725\
        );

    \I__7958\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36722\
        );

    \I__7957\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36719\
        );

    \I__7956\ : Span4Mux_h
    port map (
            O => \N__36725\,
            I => \N__36715\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__36722\,
            I => \N__36712\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__36719\,
            I => \N__36709\
        );

    \I__7953\ : InMux
    port map (
            O => \N__36718\,
            I => \N__36705\
        );

    \I__7952\ : Span4Mux_v
    port map (
            O => \N__36715\,
            I => \N__36702\
        );

    \I__7951\ : Span4Mux_h
    port map (
            O => \N__36712\,
            I => \N__36699\
        );

    \I__7950\ : Span4Mux_v
    port map (
            O => \N__36709\,
            I => \N__36696\
        );

    \I__7949\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36693\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__36705\,
            I => \N__36690\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__36702\,
            I => rand_data_19
        );

    \I__7946\ : Odrv4
    port map (
            O => \N__36699\,
            I => rand_data_19
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__36696\,
            I => rand_data_19
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__36693\,
            I => rand_data_19
        );

    \I__7943\ : Odrv12
    port map (
            O => \N__36690\,
            I => rand_data_19
        );

    \I__7942\ : InMux
    port map (
            O => \N__36679\,
            I => n15577
        );

    \I__7941\ : InMux
    port map (
            O => \N__36676\,
            I => n15578
        );

    \I__7940\ : InMux
    port map (
            O => \N__36673\,
            I => n15579
        );

    \I__7939\ : CascadeMux
    port map (
            O => \N__36670\,
            I => \N__36666\
        );

    \I__7938\ : InMux
    port map (
            O => \N__36669\,
            I => \N__36663\
        );

    \I__7937\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36660\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__36663\,
            I => rand_setpoint_22
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__36660\,
            I => rand_setpoint_22
        );

    \I__7934\ : InMux
    port map (
            O => \N__36655\,
            I => n15580
        );

    \I__7933\ : InMux
    port map (
            O => \N__36652\,
            I => n15581
        );

    \I__7932\ : InMux
    port map (
            O => \N__36649\,
            I => \bfn_13_32_0_\
        );

    \I__7931\ : CascadeMux
    port map (
            O => \N__36646\,
            I => \N__36642\
        );

    \I__7930\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36639\
        );

    \I__7929\ : InMux
    port map (
            O => \N__36642\,
            I => \N__36636\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__36639\,
            I => rand_setpoint_25
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__36636\,
            I => rand_setpoint_25
        );

    \I__7926\ : InMux
    port map (
            O => \N__36631\,
            I => n15583
        );

    \I__7925\ : InMux
    port map (
            O => \N__36628\,
            I => n15584
        );

    \I__7924\ : InMux
    port map (
            O => \N__36625\,
            I => n15585
        );

    \I__7923\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36616\
        );

    \I__7922\ : CascadeMux
    port map (
            O => \N__36621\,
            I => \N__36613\
        );

    \I__7921\ : InMux
    port map (
            O => \N__36620\,
            I => \N__36610\
        );

    \I__7920\ : InMux
    port map (
            O => \N__36619\,
            I => \N__36606\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__36616\,
            I => \N__36603\
        );

    \I__7918\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36600\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__36610\,
            I => \N__36597\
        );

    \I__7916\ : InMux
    port map (
            O => \N__36609\,
            I => \N__36593\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__36606\,
            I => \N__36590\
        );

    \I__7914\ : Span4Mux_v
    port map (
            O => \N__36603\,
            I => \N__36587\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__36600\,
            I => \N__36582\
        );

    \I__7912\ : Sp12to4
    port map (
            O => \N__36597\,
            I => \N__36582\
        );

    \I__7911\ : InMux
    port map (
            O => \N__36596\,
            I => \N__36579\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__36593\,
            I => \N__36576\
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__36590\,
            I => rand_data_10
        );

    \I__7908\ : Odrv4
    port map (
            O => \N__36587\,
            I => rand_data_10
        );

    \I__7907\ : Odrv12
    port map (
            O => \N__36582\,
            I => rand_data_10
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__36579\,
            I => rand_data_10
        );

    \I__7905\ : Odrv12
    port map (
            O => \N__36576\,
            I => rand_data_10
        );

    \I__7904\ : InMux
    port map (
            O => \N__36565\,
            I => n15568
        );

    \I__7903\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36559\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__36559\,
            I => \N__36556\
        );

    \I__7901\ : Span4Mux_s2_v
    port map (
            O => \N__36556\,
            I => \N__36552\
        );

    \I__7900\ : CascadeMux
    port map (
            O => \N__36555\,
            I => \N__36549\
        );

    \I__7899\ : Sp12to4
    port map (
            O => \N__36552\,
            I => \N__36546\
        );

    \I__7898\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36543\
        );

    \I__7897\ : Odrv12
    port map (
            O => \N__36546\,
            I => rand_setpoint_11
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__36543\,
            I => rand_setpoint_11
        );

    \I__7895\ : InMux
    port map (
            O => \N__36538\,
            I => n15569
        );

    \I__7894\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36532\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__36532\,
            I => \N__36529\
        );

    \I__7892\ : Span4Mux_h
    port map (
            O => \N__36529\,
            I => \N__36525\
        );

    \I__7891\ : InMux
    port map (
            O => \N__36528\,
            I => \N__36522\
        );

    \I__7890\ : Odrv4
    port map (
            O => \N__36525\,
            I => rand_setpoint_12
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__36522\,
            I => rand_setpoint_12
        );

    \I__7888\ : InMux
    port map (
            O => \N__36517\,
            I => n15570
        );

    \I__7887\ : InMux
    port map (
            O => \N__36514\,
            I => \N__36511\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__36511\,
            I => \N__36508\
        );

    \I__7885\ : Span4Mux_h
    port map (
            O => \N__36508\,
            I => \N__36504\
        );

    \I__7884\ : InMux
    port map (
            O => \N__36507\,
            I => \N__36501\
        );

    \I__7883\ : Odrv4
    port map (
            O => \N__36504\,
            I => rand_setpoint_13
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__36501\,
            I => rand_setpoint_13
        );

    \I__7881\ : InMux
    port map (
            O => \N__36496\,
            I => n15571
        );

    \I__7880\ : InMux
    port map (
            O => \N__36493\,
            I => \N__36489\
        );

    \I__7879\ : CascadeMux
    port map (
            O => \N__36492\,
            I => \N__36486\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__36489\,
            I => \N__36483\
        );

    \I__7877\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36480\
        );

    \I__7876\ : Odrv4
    port map (
            O => \N__36483\,
            I => rand_setpoint_14
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__36480\,
            I => rand_setpoint_14
        );

    \I__7874\ : InMux
    port map (
            O => \N__36475\,
            I => n15572
        );

    \I__7873\ : InMux
    port map (
            O => \N__36472\,
            I => \N__36469\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__36469\,
            I => \N__36466\
        );

    \I__7871\ : Span4Mux_s2_v
    port map (
            O => \N__36466\,
            I => \N__36462\
        );

    \I__7870\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36459\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__36462\,
            I => rand_setpoint_15
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__36459\,
            I => rand_setpoint_15
        );

    \I__7867\ : InMux
    port map (
            O => \N__36454\,
            I => n15573
        );

    \I__7866\ : InMux
    port map (
            O => \N__36451\,
            I => \bfn_13_31_0_\
        );

    \I__7865\ : InMux
    port map (
            O => \N__36448\,
            I => n15575
        );

    \I__7864\ : InMux
    port map (
            O => \N__36445\,
            I => n15576
        );

    \I__7863\ : InMux
    port map (
            O => \N__36442\,
            I => \N__36436\
        );

    \I__7862\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36433\
        );

    \I__7861\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36428\
        );

    \I__7860\ : InMux
    port map (
            O => \N__36439\,
            I => \N__36428\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__36436\,
            I => \N__36425\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__36433\,
            I => \N__36419\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__36428\,
            I => \N__36419\
        );

    \I__7856\ : Span4Mux_h
    port map (
            O => \N__36425\,
            I => \N__36415\
        );

    \I__7855\ : InMux
    port map (
            O => \N__36424\,
            I => \N__36412\
        );

    \I__7854\ : Span4Mux_v
    port map (
            O => \N__36419\,
            I => \N__36409\
        );

    \I__7853\ : InMux
    port map (
            O => \N__36418\,
            I => \N__36406\
        );

    \I__7852\ : Sp12to4
    port map (
            O => \N__36415\,
            I => \N__36401\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36401\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__36409\,
            I => rand_data_2
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__36406\,
            I => rand_data_2
        );

    \I__7848\ : Odrv12
    port map (
            O => \N__36401\,
            I => rand_data_2
        );

    \I__7847\ : InMux
    port map (
            O => \N__36394\,
            I => n15560
        );

    \I__7846\ : CascadeMux
    port map (
            O => \N__36391\,
            I => \N__36387\
        );

    \I__7845\ : InMux
    port map (
            O => \N__36390\,
            I => \N__36384\
        );

    \I__7844\ : InMux
    port map (
            O => \N__36387\,
            I => \N__36381\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__36384\,
            I => rand_setpoint_3
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__36381\,
            I => rand_setpoint_3
        );

    \I__7841\ : InMux
    port map (
            O => \N__36376\,
            I => n15561
        );

    \I__7840\ : CascadeMux
    port map (
            O => \N__36373\,
            I => \N__36369\
        );

    \I__7839\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36366\
        );

    \I__7838\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36363\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__36366\,
            I => rand_setpoint_4
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__36363\,
            I => rand_setpoint_4
        );

    \I__7835\ : InMux
    port map (
            O => \N__36358\,
            I => n15562
        );

    \I__7834\ : InMux
    port map (
            O => \N__36355\,
            I => n15563
        );

    \I__7833\ : InMux
    port map (
            O => \N__36352\,
            I => n15564
        );

    \I__7832\ : InMux
    port map (
            O => \N__36349\,
            I => n15565
        );

    \I__7831\ : CascadeMux
    port map (
            O => \N__36346\,
            I => \N__36343\
        );

    \I__7830\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36340\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__36340\,
            I => \N__36336\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__36339\,
            I => \N__36333\
        );

    \I__7827\ : Span4Mux_s2_v
    port map (
            O => \N__36336\,
            I => \N__36330\
        );

    \I__7826\ : InMux
    port map (
            O => \N__36333\,
            I => \N__36327\
        );

    \I__7825\ : Odrv4
    port map (
            O => \N__36330\,
            I => rand_setpoint_8
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__36327\,
            I => rand_setpoint_8
        );

    \I__7823\ : InMux
    port map (
            O => \N__36322\,
            I => \bfn_13_30_0_\
        );

    \I__7822\ : CascadeMux
    port map (
            O => \N__36319\,
            I => \N__36316\
        );

    \I__7821\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36313\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__36313\,
            I => \N__36309\
        );

    \I__7819\ : CascadeMux
    port map (
            O => \N__36312\,
            I => \N__36306\
        );

    \I__7818\ : Span4Mux_h
    port map (
            O => \N__36309\,
            I => \N__36303\
        );

    \I__7817\ : InMux
    port map (
            O => \N__36306\,
            I => \N__36300\
        );

    \I__7816\ : Odrv4
    port map (
            O => \N__36303\,
            I => rand_setpoint_9
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__36300\,
            I => rand_setpoint_9
        );

    \I__7814\ : InMux
    port map (
            O => \N__36295\,
            I => n15567
        );

    \I__7813\ : InMux
    port map (
            O => \N__36292\,
            I => n15552
        );

    \I__7812\ : InMux
    port map (
            O => \N__36289\,
            I => n15553
        );

    \I__7811\ : InMux
    port map (
            O => \N__36286\,
            I => n15554
        );

    \I__7810\ : InMux
    port map (
            O => \N__36283\,
            I => n15555
        );

    \I__7809\ : InMux
    port map (
            O => \N__36280\,
            I => n15556
        );

    \I__7808\ : InMux
    port map (
            O => \N__36277\,
            I => n15557
        );

    \I__7807\ : InMux
    port map (
            O => \N__36274\,
            I => n15558
        );

    \I__7806\ : InMux
    port map (
            O => \N__36271\,
            I => \N__36268\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__36268\,
            I => \N__36264\
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__36267\,
            I => \N__36261\
        );

    \I__7803\ : Span4Mux_h
    port map (
            O => \N__36264\,
            I => \N__36258\
        );

    \I__7802\ : InMux
    port map (
            O => \N__36261\,
            I => \N__36255\
        );

    \I__7801\ : Odrv4
    port map (
            O => \N__36258\,
            I => rand_setpoint_0
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__36255\,
            I => rand_setpoint_0
        );

    \I__7799\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36246\
        );

    \I__7798\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36242\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__36246\,
            I => \N__36239\
        );

    \I__7796\ : InMux
    port map (
            O => \N__36245\,
            I => \N__36236\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__36242\,
            I => \N__36233\
        );

    \I__7794\ : Span4Mux_v
    port map (
            O => \N__36239\,
            I => \N__36228\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__36236\,
            I => \N__36225\
        );

    \I__7792\ : Sp12to4
    port map (
            O => \N__36233\,
            I => \N__36221\
        );

    \I__7791\ : InMux
    port map (
            O => \N__36232\,
            I => \N__36218\
        );

    \I__7790\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36215\
        );

    \I__7789\ : Sp12to4
    port map (
            O => \N__36228\,
            I => \N__36212\
        );

    \I__7788\ : Span4Mux_h
    port map (
            O => \N__36225\,
            I => \N__36209\
        );

    \I__7787\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36206\
        );

    \I__7786\ : Span12Mux_h
    port map (
            O => \N__36221\,
            I => \N__36201\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__36218\,
            I => \N__36201\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__36215\,
            I => rand_data_1
        );

    \I__7783\ : Odrv12
    port map (
            O => \N__36212\,
            I => rand_data_1
        );

    \I__7782\ : Odrv4
    port map (
            O => \N__36209\,
            I => rand_data_1
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__36206\,
            I => rand_data_1
        );

    \I__7780\ : Odrv12
    port map (
            O => \N__36201\,
            I => rand_data_1
        );

    \I__7779\ : InMux
    port map (
            O => \N__36190\,
            I => n15559
        );

    \I__7778\ : InMux
    port map (
            O => \N__36187\,
            I => \bfn_13_27_0_\
        );

    \I__7777\ : InMux
    port map (
            O => \N__36184\,
            I => n15544
        );

    \I__7776\ : InMux
    port map (
            O => \N__36181\,
            I => n15545
        );

    \I__7775\ : InMux
    port map (
            O => \N__36178\,
            I => n15546
        );

    \I__7774\ : InMux
    port map (
            O => \N__36175\,
            I => n15547
        );

    \I__7773\ : InMux
    port map (
            O => \N__36172\,
            I => n15548
        );

    \I__7772\ : InMux
    port map (
            O => \N__36169\,
            I => n15549
        );

    \I__7771\ : InMux
    port map (
            O => \N__36166\,
            I => n15550
        );

    \I__7770\ : InMux
    port map (
            O => \N__36163\,
            I => \bfn_13_28_0_\
        );

    \I__7769\ : InMux
    port map (
            O => \N__36160\,
            I => n15533
        );

    \I__7768\ : InMux
    port map (
            O => \N__36157\,
            I => n15534
        );

    \I__7767\ : InMux
    port map (
            O => \N__36154\,
            I => \bfn_13_26_0_\
        );

    \I__7766\ : InMux
    port map (
            O => \N__36151\,
            I => n15536
        );

    \I__7765\ : InMux
    port map (
            O => \N__36148\,
            I => n15537
        );

    \I__7764\ : InMux
    port map (
            O => \N__36145\,
            I => n15538
        );

    \I__7763\ : InMux
    port map (
            O => \N__36142\,
            I => n15539
        );

    \I__7762\ : InMux
    port map (
            O => \N__36139\,
            I => n15540
        );

    \I__7761\ : InMux
    port map (
            O => \N__36136\,
            I => n15541
        );

    \I__7760\ : InMux
    port map (
            O => \N__36133\,
            I => n15542
        );

    \I__7759\ : InMux
    port map (
            O => \N__36130\,
            I => \N__36127\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__36127\,
            I => \N__36124\
        );

    \I__7757\ : Span4Mux_v
    port map (
            O => \N__36124\,
            I => \N__36121\
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__36121\,
            I => \c0.n17981\
        );

    \I__7755\ : CascadeMux
    port map (
            O => \N__36118\,
            I => \c0.n17984_cascade_\
        );

    \I__7754\ : InMux
    port map (
            O => \N__36115\,
            I => \N__36112\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__36112\,
            I => \c0.n22_adj_2354\
        );

    \I__7752\ : CascadeMux
    port map (
            O => \N__36109\,
            I => \N__36105\
        );

    \I__7751\ : CascadeMux
    port map (
            O => \N__36108\,
            I => \N__36102\
        );

    \I__7750\ : InMux
    port map (
            O => \N__36105\,
            I => \N__36097\
        );

    \I__7749\ : InMux
    port map (
            O => \N__36102\,
            I => \N__36097\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__36097\,
            I => data_out_frame2_17_5
        );

    \I__7747\ : InMux
    port map (
            O => \N__36094\,
            I => \bfn_13_25_0_\
        );

    \I__7746\ : InMux
    port map (
            O => \N__36091\,
            I => n15528
        );

    \I__7745\ : InMux
    port map (
            O => \N__36088\,
            I => n15529
        );

    \I__7744\ : InMux
    port map (
            O => \N__36085\,
            I => n15530
        );

    \I__7743\ : InMux
    port map (
            O => \N__36082\,
            I => n15531
        );

    \I__7742\ : InMux
    port map (
            O => \N__36079\,
            I => n15532
        );

    \I__7741\ : InMux
    port map (
            O => \N__36076\,
            I => \N__36070\
        );

    \I__7740\ : InMux
    port map (
            O => \N__36075\,
            I => \N__36066\
        );

    \I__7739\ : InMux
    port map (
            O => \N__36074\,
            I => \N__36061\
        );

    \I__7738\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36061\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36070\,
            I => \N__36058\
        );

    \I__7736\ : InMux
    port map (
            O => \N__36069\,
            I => \N__36055\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__36066\,
            I => \N__36052\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__36061\,
            I => data_out_frame2_15_3
        );

    \I__7733\ : Odrv4
    port map (
            O => \N__36058\,
            I => data_out_frame2_15_3
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__36055\,
            I => data_out_frame2_15_3
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__36052\,
            I => data_out_frame2_15_3
        );

    \I__7730\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36038\
        );

    \I__7729\ : InMux
    port map (
            O => \N__36042\,
            I => \N__36033\
        );

    \I__7728\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36033\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__36038\,
            I => data_out_frame2_13_4
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__36033\,
            I => data_out_frame2_13_4
        );

    \I__7725\ : InMux
    port map (
            O => \N__36028\,
            I => \N__36025\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__36025\,
            I => \N__36022\
        );

    \I__7723\ : Span4Mux_h
    port map (
            O => \N__36022\,
            I => \N__36019\
        );

    \I__7722\ : Odrv4
    port map (
            O => \N__36019\,
            I => \c0.n11\
        );

    \I__7721\ : InMux
    port map (
            O => \N__36016\,
            I => \N__36013\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__36013\,
            I => \N__36010\
        );

    \I__7719\ : Odrv12
    port map (
            O => \N__36010\,
            I => \c0.n9810\
        );

    \I__7718\ : InMux
    port map (
            O => \N__36007\,
            I => \N__36004\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__36004\,
            I => \N__36001\
        );

    \I__7716\ : Span4Mux_h
    port map (
            O => \N__36001\,
            I => \N__35998\
        );

    \I__7715\ : Odrv4
    port map (
            O => \N__35998\,
            I => \c0.n17_adj_2193\
        );

    \I__7714\ : CascadeMux
    port map (
            O => \N__35995\,
            I => \c0.n16_cascade_\
        );

    \I__7713\ : CascadeMux
    port map (
            O => \N__35992\,
            I => \c0.n17112_cascade_\
        );

    \I__7712\ : CascadeMux
    port map (
            O => \N__35989\,
            I => \c0.n14_adj_2308_cascade_\
        );

    \I__7711\ : CascadeMux
    port map (
            O => \N__35986\,
            I => \N__35983\
        );

    \I__7710\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35980\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__35980\,
            I => \N__35977\
        );

    \I__7708\ : Span12Mux_h
    port map (
            O => \N__35977\,
            I => \N__35974\
        );

    \I__7707\ : Odrv12
    port map (
            O => \N__35974\,
            I => \c0.data_out_frame2_19_5\
        );

    \I__7706\ : InMux
    port map (
            O => \N__35971\,
            I => \N__35968\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__35968\,
            I => \N__35965\
        );

    \I__7704\ : Span4Mux_v
    port map (
            O => \N__35965\,
            I => \N__35962\
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__35962\,
            I => \c0.n17933\
        );

    \I__7702\ : InMux
    port map (
            O => \N__35959\,
            I => \N__35956\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__35956\,
            I => \N__35953\
        );

    \I__7700\ : Odrv4
    port map (
            O => \N__35953\,
            I => \c0.n5_adj_2317\
        );

    \I__7699\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35947\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__35947\,
            I => \N__35944\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__35944\,
            I => \c0.n16957\
        );

    \I__7696\ : CascadeMux
    port map (
            O => \N__35941\,
            I => \N__35938\
        );

    \I__7695\ : InMux
    port map (
            O => \N__35938\,
            I => \N__35934\
        );

    \I__7694\ : InMux
    port map (
            O => \N__35937\,
            I => \N__35931\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__35934\,
            I => \N__35928\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__35931\,
            I => \N__35925\
        );

    \I__7691\ : Span4Mux_h
    port map (
            O => \N__35928\,
            I => \N__35922\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__35925\,
            I => \c0.n17106\
        );

    \I__7689\ : Odrv4
    port map (
            O => \N__35922\,
            I => \c0.n17106\
        );

    \I__7688\ : CascadeMux
    port map (
            O => \N__35917\,
            I => \c0.n16957_cascade_\
        );

    \I__7687\ : InMux
    port map (
            O => \N__35914\,
            I => \N__35911\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__35911\,
            I => \c0.n15_adj_2269\
        );

    \I__7685\ : CascadeMux
    port map (
            O => \N__35908\,
            I => \N__35905\
        );

    \I__7684\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35902\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__35902\,
            I => \N__35899\
        );

    \I__7682\ : Span4Mux_v
    port map (
            O => \N__35899\,
            I => \N__35896\
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__35896\,
            I => \c0.data_out_frame2_20_1\
        );

    \I__7680\ : InMux
    port map (
            O => \N__35893\,
            I => \N__35887\
        );

    \I__7679\ : InMux
    port map (
            O => \N__35892\,
            I => \N__35887\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__35887\,
            I => \c0.n17061\
        );

    \I__7677\ : InMux
    port map (
            O => \N__35884\,
            I => \N__35881\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__35881\,
            I => \N__35878\
        );

    \I__7675\ : Odrv4
    port map (
            O => \N__35878\,
            I => \c0.data_out_frame2_20_0\
        );

    \I__7674\ : InMux
    port map (
            O => \N__35875\,
            I => \N__35870\
        );

    \I__7673\ : InMux
    port map (
            O => \N__35874\,
            I => \N__35866\
        );

    \I__7672\ : InMux
    port map (
            O => \N__35873\,
            I => \N__35863\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__35870\,
            I => \N__35860\
        );

    \I__7670\ : InMux
    port map (
            O => \N__35869\,
            I => \N__35857\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__35866\,
            I => \N__35854\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__35863\,
            I => \N__35846\
        );

    \I__7667\ : Span4Mux_h
    port map (
            O => \N__35860\,
            I => \N__35846\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__35857\,
            I => \N__35846\
        );

    \I__7665\ : Span4Mux_v
    port map (
            O => \N__35854\,
            I => \N__35843\
        );

    \I__7664\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35840\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__35846\,
            I => \N__35837\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__35843\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__35840\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__7660\ : Odrv4
    port map (
            O => \N__35837\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__7659\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35827\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__35827\,
            I => \N__35824\
        );

    \I__7657\ : Span4Mux_h
    port map (
            O => \N__35824\,
            I => \N__35821\
        );

    \I__7656\ : Odrv4
    port map (
            O => \N__35821\,
            I => \c0.n17578\
        );

    \I__7655\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35815\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__35815\,
            I => \N__35811\
        );

    \I__7653\ : CascadeMux
    port map (
            O => \N__35814\,
            I => \N__35806\
        );

    \I__7652\ : Span4Mux_v
    port map (
            O => \N__35811\,
            I => \N__35803\
        );

    \I__7651\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35800\
        );

    \I__7650\ : InMux
    port map (
            O => \N__35809\,
            I => \N__35797\
        );

    \I__7649\ : InMux
    port map (
            O => \N__35806\,
            I => \N__35794\
        );

    \I__7648\ : Span4Mux_h
    port map (
            O => \N__35803\,
            I => \N__35791\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35788\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__35797\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__35794\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__7644\ : Odrv4
    port map (
            O => \N__35791\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__35788\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__7642\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35776\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__35776\,
            I => \c0.n6_adj_2335\
        );

    \I__7640\ : CascadeMux
    port map (
            O => \N__35773\,
            I => \N__35769\
        );

    \I__7639\ : CascadeMux
    port map (
            O => \N__35772\,
            I => \N__35764\
        );

    \I__7638\ : InMux
    port map (
            O => \N__35769\,
            I => \N__35753\
        );

    \I__7637\ : InMux
    port map (
            O => \N__35768\,
            I => \N__35753\
        );

    \I__7636\ : InMux
    port map (
            O => \N__35767\,
            I => \N__35753\
        );

    \I__7635\ : InMux
    port map (
            O => \N__35764\,
            I => \N__35746\
        );

    \I__7634\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35746\
        );

    \I__7633\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35746\
        );

    \I__7632\ : InMux
    port map (
            O => \N__35761\,
            I => \N__35742\
        );

    \I__7631\ : CascadeMux
    port map (
            O => \N__35760\,
            I => \N__35739\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__35753\,
            I => \N__35734\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__35746\,
            I => \N__35734\
        );

    \I__7628\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35731\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__35742\,
            I => \N__35728\
        );

    \I__7626\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35725\
        );

    \I__7625\ : Span4Mux_s3_v
    port map (
            O => \N__35734\,
            I => \N__35722\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__35731\,
            I => \N__35717\
        );

    \I__7623\ : Span4Mux_v
    port map (
            O => \N__35728\,
            I => \N__35717\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__35725\,
            I => \N__35714\
        );

    \I__7621\ : Span4Mux_h
    port map (
            O => \N__35722\,
            I => \N__35711\
        );

    \I__7620\ : Span4Mux_h
    port map (
            O => \N__35717\,
            I => \N__35708\
        );

    \I__7619\ : Odrv12
    port map (
            O => \N__35714\,
            I => \c0.n10181\
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__35711\,
            I => \c0.n10181\
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__35708\,
            I => \c0.n10181\
        );

    \I__7616\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35697\
        );

    \I__7615\ : InMux
    port map (
            O => \N__35700\,
            I => \N__35694\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__35697\,
            I => \N__35691\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__35694\,
            I => \c0.data_out_6_6\
        );

    \I__7612\ : Odrv4
    port map (
            O => \N__35691\,
            I => \c0.data_out_6_6\
        );

    \I__7611\ : InMux
    port map (
            O => \N__35686\,
            I => \N__35683\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__35683\,
            I => \c0.n5_adj_2300\
        );

    \I__7609\ : CascadeMux
    port map (
            O => \N__35680\,
            I => \c0.n17555_cascade_\
        );

    \I__7608\ : InMux
    port map (
            O => \N__35677\,
            I => \N__35674\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__35674\,
            I => \N__35671\
        );

    \I__7606\ : Odrv4
    port map (
            O => \N__35671\,
            I => \c0.n18035\
        );

    \I__7605\ : InMux
    port map (
            O => \N__35668\,
            I => \N__35665\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__35665\,
            I => \N__35662\
        );

    \I__7603\ : Odrv4
    port map (
            O => \N__35662\,
            I => \c0.n17569\
        );

    \I__7602\ : InMux
    port map (
            O => \N__35659\,
            I => \N__35656\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__35656\,
            I => \c0.n16912\
        );

    \I__7600\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35650\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__35650\,
            I => \N__35647\
        );

    \I__7598\ : Span4Mux_h
    port map (
            O => \N__35647\,
            I => \N__35644\
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__35644\,
            I => \c0.n21\
        );

    \I__7596\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35638\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__35638\,
            I => \c0.n17588\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__35635\,
            I => \N__35632\
        );

    \I__7593\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35629\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__35629\,
            I => \N__35626\
        );

    \I__7591\ : Span4Mux_s3_v
    port map (
            O => \N__35626\,
            I => \N__35623\
        );

    \I__7590\ : Odrv4
    port map (
            O => \N__35623\,
            I => \c0.n1\
        );

    \I__7589\ : CascadeMux
    port map (
            O => \N__35620\,
            I => \n18038_cascade_\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__35617\,
            I => \N__35612\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__35616\,
            I => \N__35609\
        );

    \I__7586\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35606\
        );

    \I__7585\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35599\
        );

    \I__7584\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35596\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__35606\,
            I => \N__35593\
        );

    \I__7582\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35590\
        );

    \I__7581\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35587\
        );

    \I__7580\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35584\
        );

    \I__7579\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35581\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__35599\,
            I => \N__35576\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__35596\,
            I => \N__35576\
        );

    \I__7576\ : Span4Mux_s3_v
    port map (
            O => \N__35593\,
            I => \N__35571\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__35590\,
            I => \N__35571\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__35587\,
            I => \N__35568\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__35584\,
            I => \N__35565\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__35581\,
            I => \N__35561\
        );

    \I__7571\ : Span4Mux_h
    port map (
            O => \N__35576\,
            I => \N__35556\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__35571\,
            I => \N__35556\
        );

    \I__7569\ : Span4Mux_v
    port map (
            O => \N__35568\,
            I => \N__35551\
        );

    \I__7568\ : Span4Mux_s1_v
    port map (
            O => \N__35565\,
            I => \N__35551\
        );

    \I__7567\ : InMux
    port map (
            O => \N__35564\,
            I => \N__35548\
        );

    \I__7566\ : Span4Mux_v
    port map (
            O => \N__35561\,
            I => \N__35545\
        );

    \I__7565\ : Span4Mux_h
    port map (
            O => \N__35556\,
            I => \N__35542\
        );

    \I__7564\ : Span4Mux_h
    port map (
            O => \N__35551\,
            I => \N__35539\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35534\
        );

    \I__7562\ : Sp12to4
    port map (
            O => \N__35545\,
            I => \N__35534\
        );

    \I__7561\ : Odrv4
    port map (
            O => \N__35542\,
            I => n8730
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__35539\,
            I => n8730
        );

    \I__7559\ : Odrv12
    port map (
            O => \N__35534\,
            I => n8730
        );

    \I__7558\ : CascadeMux
    port map (
            O => \N__35527\,
            I => \n10_adj_2413_cascade_\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__35524\,
            I => \N__35515\
        );

    \I__7556\ : InMux
    port map (
            O => \N__35523\,
            I => \N__35512\
        );

    \I__7555\ : InMux
    port map (
            O => \N__35522\,
            I => \N__35508\
        );

    \I__7554\ : InMux
    port map (
            O => \N__35521\,
            I => \N__35505\
        );

    \I__7553\ : InMux
    port map (
            O => \N__35520\,
            I => \N__35500\
        );

    \I__7552\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35500\
        );

    \I__7551\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35497\
        );

    \I__7550\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35494\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__35512\,
            I => \N__35491\
        );

    \I__7548\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35487\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__35508\,
            I => \N__35484\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__35505\,
            I => \N__35479\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35479\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__35497\,
            I => \N__35472\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__35494\,
            I => \N__35472\
        );

    \I__7542\ : Span4Mux_h
    port map (
            O => \N__35491\,
            I => \N__35472\
        );

    \I__7541\ : InMux
    port map (
            O => \N__35490\,
            I => \N__35468\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__35487\,
            I => \N__35465\
        );

    \I__7539\ : Span4Mux_s1_v
    port map (
            O => \N__35484\,
            I => \N__35460\
        );

    \I__7538\ : Span4Mux_v
    port map (
            O => \N__35479\,
            I => \N__35460\
        );

    \I__7537\ : Span4Mux_h
    port map (
            O => \N__35472\,
            I => \N__35457\
        );

    \I__7536\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35454\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__35468\,
            I => byte_transmit_counter_4
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__35465\,
            I => byte_transmit_counter_4
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__35460\,
            I => byte_transmit_counter_4
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__35457\,
            I => byte_transmit_counter_4
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__35454\,
            I => byte_transmit_counter_4
        );

    \I__7530\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35440\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__35440\,
            I => \N__35437\
        );

    \I__7528\ : Span4Mux_s3_h
    port map (
            O => \N__35437\,
            I => \N__35434\
        );

    \I__7527\ : Span4Mux_h
    port map (
            O => \N__35434\,
            I => \N__35430\
        );

    \I__7526\ : InMux
    port map (
            O => \N__35433\,
            I => \N__35427\
        );

    \I__7525\ : Span4Mux_h
    port map (
            O => \N__35430\,
            I => \N__35424\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__35427\,
            I => \r_Tx_Data_6\
        );

    \I__7523\ : Odrv4
    port map (
            O => \N__35424\,
            I => \r_Tx_Data_6\
        );

    \I__7522\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35416\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__35416\,
            I => \N__35413\
        );

    \I__7520\ : Span4Mux_s1_v
    port map (
            O => \N__35413\,
            I => \N__35410\
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__35410\,
            I => \c0.data_out_1_1\
        );

    \I__7518\ : CascadeMux
    port map (
            O => \N__35407\,
            I => \c0.n8_adj_2348_cascade_\
        );

    \I__7517\ : InMux
    port map (
            O => \N__35404\,
            I => \N__35401\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__35401\,
            I => \N__35398\
        );

    \I__7515\ : Span4Mux_h
    port map (
            O => \N__35398\,
            I => \N__35395\
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__35395\,
            I => \c0.n17900\
        );

    \I__7513\ : CascadeMux
    port map (
            O => \N__35392\,
            I => \N__35387\
        );

    \I__7512\ : CascadeMux
    port map (
            O => \N__35391\,
            I => \N__35382\
        );

    \I__7511\ : CascadeMux
    port map (
            O => \N__35390\,
            I => \N__35377\
        );

    \I__7510\ : InMux
    port map (
            O => \N__35387\,
            I => \N__35374\
        );

    \I__7509\ : InMux
    port map (
            O => \N__35386\,
            I => \N__35369\
        );

    \I__7508\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35369\
        );

    \I__7507\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35360\
        );

    \I__7506\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35360\
        );

    \I__7505\ : InMux
    port map (
            O => \N__35380\,
            I => \N__35360\
        );

    \I__7504\ : InMux
    port map (
            O => \N__35377\,
            I => \N__35360\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__35374\,
            I => \N__35357\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__35369\,
            I => \r_Bit_Index_1_adj_2456\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__35360\,
            I => \r_Bit_Index_1_adj_2456\
        );

    \I__7500\ : Odrv4
    port map (
            O => \N__35357\,
            I => \r_Bit_Index_1_adj_2456\
        );

    \I__7499\ : InMux
    port map (
            O => \N__35350\,
            I => \N__35344\
        );

    \I__7498\ : InMux
    port map (
            O => \N__35349\,
            I => \N__35335\
        );

    \I__7497\ : InMux
    port map (
            O => \N__35348\,
            I => \N__35335\
        );

    \I__7496\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35335\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__35344\,
            I => \N__35332\
        );

    \I__7494\ : InMux
    port map (
            O => \N__35343\,
            I => \N__35329\
        );

    \I__7493\ : InMux
    port map (
            O => \N__35342\,
            I => \N__35326\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__35335\,
            I => \N__35321\
        );

    \I__7491\ : Span4Mux_v
    port map (
            O => \N__35332\,
            I => \N__35321\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__35329\,
            I => \r_Bit_Index_0_adj_2457\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__35326\,
            I => \r_Bit_Index_0_adj_2457\
        );

    \I__7488\ : Odrv4
    port map (
            O => \N__35321\,
            I => \r_Bit_Index_0_adj_2457\
        );

    \I__7487\ : InMux
    port map (
            O => \N__35314\,
            I => \N__35311\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__35311\,
            I => \N__35308\
        );

    \I__7485\ : Odrv4
    port map (
            O => \N__35308\,
            I => \c0.tx2.n17903\
        );

    \I__7484\ : InMux
    port map (
            O => \N__35305\,
            I => \N__35301\
        );

    \I__7483\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35298\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__35301\,
            I => \c0.n16975\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__35298\,
            I => \c0.n16975\
        );

    \I__7480\ : CascadeMux
    port map (
            O => \N__35293\,
            I => \c0.n16978_cascade_\
        );

    \I__7479\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35287\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__35287\,
            I => \N__35283\
        );

    \I__7477\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35280\
        );

    \I__7476\ : Span4Mux_v
    port map (
            O => \N__35283\,
            I => \N__35277\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__35280\,
            I => data_out_0_3
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__35277\,
            I => data_out_0_3
        );

    \I__7473\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35268\
        );

    \I__7472\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35265\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__35268\,
            I => data_out_2_2
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__35265\,
            I => data_out_2_2
        );

    \I__7469\ : InMux
    port map (
            O => \N__35260\,
            I => \N__35257\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__35257\,
            I => \N__35254\
        );

    \I__7467\ : Span4Mux_v
    port map (
            O => \N__35254\,
            I => \N__35251\
        );

    \I__7466\ : Odrv4
    port map (
            O => \N__35251\,
            I => \c0.n2_adj_2291\
        );

    \I__7465\ : InMux
    port map (
            O => \N__35248\,
            I => \N__35242\
        );

    \I__7464\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35242\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__35242\,
            I => data_out_3_2
        );

    \I__7462\ : CascadeMux
    port map (
            O => \N__35239\,
            I => \N__35233\
        );

    \I__7461\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35227\
        );

    \I__7460\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35227\
        );

    \I__7459\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35224\
        );

    \I__7458\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35219\
        );

    \I__7457\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35219\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__35227\,
            I => \N__35216\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__35224\,
            I => \N__35212\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__35219\,
            I => \N__35209\
        );

    \I__7453\ : Span4Mux_v
    port map (
            O => \N__35216\,
            I => \N__35206\
        );

    \I__7452\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35203\
        );

    \I__7451\ : Span4Mux_h
    port map (
            O => \N__35212\,
            I => \N__35200\
        );

    \I__7450\ : Span4Mux_v
    port map (
            O => \N__35209\,
            I => \N__35197\
        );

    \I__7449\ : Span4Mux_h
    port map (
            O => \N__35206\,
            I => \N__35194\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__35203\,
            I => data_out_frame2_9_4
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__35200\,
            I => data_out_frame2_9_4
        );

    \I__7446\ : Odrv4
    port map (
            O => \N__35197\,
            I => data_out_frame2_9_4
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__35194\,
            I => data_out_frame2_9_4
        );

    \I__7444\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35182\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__35182\,
            I => \N__35179\
        );

    \I__7442\ : Sp12to4
    port map (
            O => \N__35179\,
            I => \N__35176\
        );

    \I__7441\ : Odrv12
    port map (
            O => \N__35176\,
            I => \c0.n9_adj_2347\
        );

    \I__7440\ : InMux
    port map (
            O => \N__35173\,
            I => \N__35170\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__35170\,
            I => \c0.n17897\
        );

    \I__7438\ : InMux
    port map (
            O => \N__35167\,
            I => \N__35160\
        );

    \I__7437\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35160\
        );

    \I__7436\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35156\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__35160\,
            I => \N__35153\
        );

    \I__7434\ : InMux
    port map (
            O => \N__35159\,
            I => \N__35150\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__35156\,
            I => data_out_frame2_10_2
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__35153\,
            I => data_out_frame2_10_2
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__35150\,
            I => data_out_frame2_10_2
        );

    \I__7430\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35140\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__35140\,
            I => \N__35137\
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__35137\,
            I => \c0.n12_adj_2305\
        );

    \I__7427\ : InMux
    port map (
            O => \N__35134\,
            I => \N__35131\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__35131\,
            I => \c0.n17990\
        );

    \I__7425\ : CascadeMux
    port map (
            O => \N__35128\,
            I => \c0.n17993_cascade_\
        );

    \I__7424\ : InMux
    port map (
            O => \N__35125\,
            I => \N__35122\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__35122\,
            I => \c0.n17894\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__35119\,
            I => \c0.n17393_cascade_\
        );

    \I__7421\ : InMux
    port map (
            O => \N__35116\,
            I => \N__35113\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__35113\,
            I => \N__35110\
        );

    \I__7419\ : Odrv4
    port map (
            O => \N__35110\,
            I => \c0.n17571\
        );

    \I__7418\ : CascadeMux
    port map (
            O => \N__35107\,
            I => \c0.n17963_cascade_\
        );

    \I__7417\ : CascadeMux
    port map (
            O => \N__35104\,
            I => \c0.n17966_cascade_\
        );

    \I__7416\ : InMux
    port map (
            O => \N__35101\,
            I => \N__35098\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__35098\,
            I => \N__35095\
        );

    \I__7414\ : Span4Mux_v
    port map (
            O => \N__35095\,
            I => \N__35092\
        );

    \I__7413\ : Odrv4
    port map (
            O => \N__35092\,
            I => \c0.tx2.r_Tx_Data_5\
        );

    \I__7412\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35086\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__35086\,
            I => \N__35082\
        );

    \I__7410\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35079\
        );

    \I__7409\ : Span4Mux_v
    port map (
            O => \N__35082\,
            I => \N__35076\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__35079\,
            I => data_out_0_5
        );

    \I__7407\ : Odrv4
    port map (
            O => \N__35076\,
            I => data_out_0_5
        );

    \I__7406\ : CascadeMux
    port map (
            O => \N__35071\,
            I => \N__35068\
        );

    \I__7405\ : InMux
    port map (
            O => \N__35068\,
            I => \N__35065\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__35065\,
            I => \N__35059\
        );

    \I__7403\ : InMux
    port map (
            O => \N__35064\,
            I => \N__35056\
        );

    \I__7402\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35053\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35062\,
            I => \N__35050\
        );

    \I__7400\ : Span4Mux_h
    port map (
            O => \N__35059\,
            I => \N__35047\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__35056\,
            I => data_out_frame2_5_3
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__35053\,
            I => data_out_frame2_5_3
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__35050\,
            I => data_out_frame2_5_3
        );

    \I__7396\ : Odrv4
    port map (
            O => \N__35047\,
            I => data_out_frame2_5_3
        );

    \I__7395\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35031\
        );

    \I__7394\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35028\
        );

    \I__7393\ : InMux
    port map (
            O => \N__35036\,
            I => \N__35025\
        );

    \I__7392\ : InMux
    port map (
            O => \N__35035\,
            I => \N__35022\
        );

    \I__7391\ : InMux
    port map (
            O => \N__35034\,
            I => \N__35019\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__35014\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__35028\,
            I => \N__35005\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__35025\,
            I => \N__35005\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__35022\,
            I => \N__35005\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__35019\,
            I => \N__35005\
        );

    \I__7385\ : InMux
    port map (
            O => \N__35018\,
            I => \N__35001\
        );

    \I__7384\ : InMux
    port map (
            O => \N__35017\,
            I => \N__34998\
        );

    \I__7383\ : Span4Mux_h
    port map (
            O => \N__35014\,
            I => \N__34993\
        );

    \I__7382\ : Span4Mux_v
    port map (
            O => \N__35005\,
            I => \N__34993\
        );

    \I__7381\ : InMux
    port map (
            O => \N__35004\,
            I => \N__34990\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__35001\,
            I => \c0.n16148\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__34998\,
            I => \c0.n16148\
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__34993\,
            I => \c0.n16148\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__34990\,
            I => \c0.n16148\
        );

    \I__7376\ : CascadeMux
    port map (
            O => \N__34981\,
            I => \c0.n17331_cascade_\
        );

    \I__7375\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34973\
        );

    \I__7374\ : InMux
    port map (
            O => \N__34977\,
            I => \N__34970\
        );

    \I__7373\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34967\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__34973\,
            I => \N__34964\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__34970\,
            I => \N__34961\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__34967\,
            I => \N__34958\
        );

    \I__7369\ : Span4Mux_v
    port map (
            O => \N__34964\,
            I => \N__34953\
        );

    \I__7368\ : Span4Mux_h
    port map (
            O => \N__34961\,
            I => \N__34950\
        );

    \I__7367\ : Span4Mux_h
    port map (
            O => \N__34958\,
            I => \N__34947\
        );

    \I__7366\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34944\
        );

    \I__7365\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34941\
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__34953\,
            I => \c0.n15846\
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__34950\,
            I => \c0.n15846\
        );

    \I__7362\ : Odrv4
    port map (
            O => \N__34947\,
            I => \c0.n15846\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__34944\,
            I => \c0.n15846\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__34941\,
            I => \c0.n15846\
        );

    \I__7359\ : InMux
    port map (
            O => \N__34930\,
            I => \N__34927\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__34927\,
            I => \c0.n17891\
        );

    \I__7357\ : InMux
    port map (
            O => \N__34924\,
            I => \N__34921\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__34921\,
            I => \N__34918\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__34918\,
            I => \c0.n17939\
        );

    \I__7354\ : InMux
    port map (
            O => \N__34915\,
            I => \N__34909\
        );

    \I__7353\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34906\
        );

    \I__7352\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34903\
        );

    \I__7351\ : InMux
    port map (
            O => \N__34912\,
            I => \N__34900\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__34909\,
            I => data_out_frame2_6_3
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__34906\,
            I => data_out_frame2_6_3
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__34903\,
            I => data_out_frame2_6_3
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__34900\,
            I => data_out_frame2_6_3
        );

    \I__7346\ : CascadeMux
    port map (
            O => \N__34891\,
            I => \N__34888\
        );

    \I__7345\ : InMux
    port map (
            O => \N__34888\,
            I => \N__34885\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__34885\,
            I => \N__34882\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__34882\,
            I => \N__34879\
        );

    \I__7342\ : Odrv4
    port map (
            O => \N__34879\,
            I => \c0.n16_adj_2197\
        );

    \I__7341\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34873\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__34873\,
            I => \N__34870\
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__34870\,
            I => \c0.n22_adj_2194\
        );

    \I__7338\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34864\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__34864\,
            I => \N__34861\
        );

    \I__7336\ : Odrv4
    port map (
            O => \N__34861\,
            I => \c0.n9754\
        );

    \I__7335\ : CascadeMux
    port map (
            O => \N__34858\,
            I => \c0.n9901_cascade_\
        );

    \I__7334\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34852\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__34852\,
            I => \c0.n6_adj_2201\
        );

    \I__7332\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34846\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__34846\,
            I => \c0.n17942\
        );

    \I__7330\ : CascadeMux
    port map (
            O => \N__34843\,
            I => \N__34840\
        );

    \I__7329\ : InMux
    port map (
            O => \N__34840\,
            I => \N__34837\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__34837\,
            I => \N__34834\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__34834\,
            I => \N__34831\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__34831\,
            I => \c0.n17560\
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__34828\,
            I => \c0.n17301_cascade_\
        );

    \I__7324\ : CascadeMux
    port map (
            O => \N__34825\,
            I => \c0.n17303_cascade_\
        );

    \I__7323\ : InMux
    port map (
            O => \N__34822\,
            I => \N__34819\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__34819\,
            I => \N__34816\
        );

    \I__7321\ : Span4Mux_h
    port map (
            O => \N__34816\,
            I => \N__34813\
        );

    \I__7320\ : Span4Mux_v
    port map (
            O => \N__34813\,
            I => \N__34810\
        );

    \I__7319\ : Odrv4
    port map (
            O => \N__34810\,
            I => \c0.tx2.r_Tx_Data_0\
        );

    \I__7318\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34803\
        );

    \I__7317\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34800\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34797\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__34800\,
            I => data_out_frame2_18_0
        );

    \I__7314\ : Odrv4
    port map (
            O => \N__34797\,
            I => data_out_frame2_18_0
        );

    \I__7313\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34789\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__34789\,
            I => \N__34786\
        );

    \I__7311\ : Span4Mux_v
    port map (
            O => \N__34786\,
            I => \N__34782\
        );

    \I__7310\ : InMux
    port map (
            O => \N__34785\,
            I => \N__34779\
        );

    \I__7309\ : Span4Mux_h
    port map (
            O => \N__34782\,
            I => \N__34776\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__34779\,
            I => data_out_frame2_17_0
        );

    \I__7307\ : Odrv4
    port map (
            O => \N__34776\,
            I => data_out_frame2_17_0
        );

    \I__7306\ : CascadeMux
    port map (
            O => \N__34771\,
            I => \c0.n18101_cascade_\
        );

    \I__7305\ : CascadeMux
    port map (
            O => \N__34768\,
            I => \c0.n18104_cascade_\
        );

    \I__7304\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34762\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__34762\,
            I => \c0.n22_adj_2337\
        );

    \I__7302\ : InMux
    port map (
            O => \N__34759\,
            I => \c0.n15618\
        );

    \I__7301\ : InMux
    port map (
            O => \N__34756\,
            I => \N__34753\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__34753\,
            I => \N__34749\
        );

    \I__7299\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34746\
        );

    \I__7298\ : Span4Mux_h
    port map (
            O => \N__34749\,
            I => \N__34743\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__34746\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__7296\ : Odrv4
    port map (
            O => \N__34743\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__7295\ : InMux
    port map (
            O => \N__34738\,
            I => \c0.n15619\
        );

    \I__7294\ : CascadeMux
    port map (
            O => \N__34735\,
            I => \N__34732\
        );

    \I__7293\ : InMux
    port map (
            O => \N__34732\,
            I => \N__34729\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__34729\,
            I => \N__34725\
        );

    \I__7291\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34722\
        );

    \I__7290\ : Span4Mux_h
    port map (
            O => \N__34725\,
            I => \N__34719\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__34722\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__34719\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__7287\ : InMux
    port map (
            O => \N__34714\,
            I => \c0.n15620\
        );

    \I__7286\ : InMux
    port map (
            O => \N__34711\,
            I => \c0.n15621\
        );

    \I__7285\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34705\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__34705\,
            I => \N__34701\
        );

    \I__7283\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34698\
        );

    \I__7282\ : Span4Mux_h
    port map (
            O => \N__34701\,
            I => \N__34695\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__34698\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__34695\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__7279\ : CEMux
    port map (
            O => \N__34690\,
            I => \N__34687\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__34687\,
            I => \N__34684\
        );

    \I__7277\ : Span4Mux_h
    port map (
            O => \N__34684\,
            I => \N__34680\
        );

    \I__7276\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34677\
        );

    \I__7275\ : Odrv4
    port map (
            O => \N__34680\,
            I => \c0.n10052\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__34677\,
            I => \c0.n10052\
        );

    \I__7273\ : SRMux
    port map (
            O => \N__34672\,
            I => \N__34669\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34666\
        );

    \I__7271\ : Odrv12
    port map (
            O => \N__34666\,
            I => \c0.n10297\
        );

    \I__7270\ : InMux
    port map (
            O => \N__34663\,
            I => \N__34656\
        );

    \I__7269\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34638\
        );

    \I__7268\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34635\
        );

    \I__7267\ : InMux
    port map (
            O => \N__34660\,
            I => \N__34632\
        );

    \I__7266\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34629\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__34656\,
            I => \N__34626\
        );

    \I__7264\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34623\
        );

    \I__7263\ : InMux
    port map (
            O => \N__34654\,
            I => \N__34620\
        );

    \I__7262\ : InMux
    port map (
            O => \N__34653\,
            I => \N__34617\
        );

    \I__7261\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34614\
        );

    \I__7260\ : InMux
    port map (
            O => \N__34651\,
            I => \N__34610\
        );

    \I__7259\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34607\
        );

    \I__7258\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34604\
        );

    \I__7257\ : InMux
    port map (
            O => \N__34648\,
            I => \N__34601\
        );

    \I__7256\ : InMux
    port map (
            O => \N__34647\,
            I => \N__34598\
        );

    \I__7255\ : InMux
    port map (
            O => \N__34646\,
            I => \N__34595\
        );

    \I__7254\ : InMux
    port map (
            O => \N__34645\,
            I => \N__34592\
        );

    \I__7253\ : InMux
    port map (
            O => \N__34644\,
            I => \N__34589\
        );

    \I__7252\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34586\
        );

    \I__7251\ : InMux
    port map (
            O => \N__34642\,
            I => \N__34583\
        );

    \I__7250\ : InMux
    port map (
            O => \N__34641\,
            I => \N__34580\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__34638\,
            I => \N__34577\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__34635\,
            I => \N__34574\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__34632\,
            I => \N__34565\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__34629\,
            I => \N__34565\
        );

    \I__7245\ : Span4Mux_s1_h
    port map (
            O => \N__34626\,
            I => \N__34565\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__34623\,
            I => \N__34565\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__34620\,
            I => \N__34555\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__34617\,
            I => \N__34550\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__34614\,
            I => \N__34550\
        );

    \I__7240\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34547\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__34610\,
            I => \N__34544\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__34607\,
            I => \N__34537\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__34604\,
            I => \N__34537\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__34601\,
            I => \N__34537\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__34598\,
            I => \N__34530\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__34595\,
            I => \N__34530\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__34592\,
            I => \N__34530\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34527\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__34586\,
            I => \N__34524\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__34583\,
            I => \N__34521\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__34580\,
            I => \N__34516\
        );

    \I__7228\ : Span4Mux_v
    port map (
            O => \N__34577\,
            I => \N__34516\
        );

    \I__7227\ : Span4Mux_v
    port map (
            O => \N__34574\,
            I => \N__34511\
        );

    \I__7226\ : Span4Mux_v
    port map (
            O => \N__34565\,
            I => \N__34511\
        );

    \I__7225\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34508\
        );

    \I__7224\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34505\
        );

    \I__7223\ : InMux
    port map (
            O => \N__34562\,
            I => \N__34502\
        );

    \I__7222\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34499\
        );

    \I__7221\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34496\
        );

    \I__7220\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34493\
        );

    \I__7219\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34490\
        );

    \I__7218\ : Span4Mux_h
    port map (
            O => \N__34555\,
            I => \N__34485\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__34550\,
            I => \N__34485\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__34547\,
            I => \N__34476\
        );

    \I__7215\ : Span4Mux_h
    port map (
            O => \N__34544\,
            I => \N__34476\
        );

    \I__7214\ : Span4Mux_v
    port map (
            O => \N__34537\,
            I => \N__34476\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__34530\,
            I => \N__34476\
        );

    \I__7212\ : Span4Mux_v
    port map (
            O => \N__34527\,
            I => \N__34467\
        );

    \I__7211\ : Span4Mux_v
    port map (
            O => \N__34524\,
            I => \N__34467\
        );

    \I__7210\ : Span4Mux_v
    port map (
            O => \N__34521\,
            I => \N__34467\
        );

    \I__7209\ : Span4Mux_h
    port map (
            O => \N__34516\,
            I => \N__34467\
        );

    \I__7208\ : Span4Mux_h
    port map (
            O => \N__34511\,
            I => \N__34464\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__34508\,
            I => \c0.n7\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__34505\,
            I => \c0.n7\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__34502\,
            I => \c0.n7\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__34499\,
            I => \c0.n7\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__34496\,
            I => \c0.n7\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__34493\,
            I => \c0.n7\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__34490\,
            I => \c0.n7\
        );

    \I__7200\ : Odrv4
    port map (
            O => \N__34485\,
            I => \c0.n7\
        );

    \I__7199\ : Odrv4
    port map (
            O => \N__34476\,
            I => \c0.n7\
        );

    \I__7198\ : Odrv4
    port map (
            O => \N__34467\,
            I => \c0.n7\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__34464\,
            I => \c0.n7\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__34441\,
            I => \N__34438\
        );

    \I__7195\ : InMux
    port map (
            O => \N__34438\,
            I => \N__34435\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__34435\,
            I => \N__34432\
        );

    \I__7193\ : Span4Mux_h
    port map (
            O => \N__34432\,
            I => \N__34427\
        );

    \I__7192\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34424\
        );

    \I__7191\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34421\
        );

    \I__7190\ : Span4Mux_h
    port map (
            O => \N__34427\,
            I => \N__34418\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__34424\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__34421\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__34418\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__7186\ : SRMux
    port map (
            O => \N__34411\,
            I => \N__34408\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__34408\,
            I => \c0.n16455\
        );

    \I__7184\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34402\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__34402\,
            I => \c0.n17927\
        );

    \I__7182\ : CascadeMux
    port map (
            O => \N__34399\,
            I => \N__34396\
        );

    \I__7181\ : InMux
    port map (
            O => \N__34396\,
            I => \N__34393\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__34393\,
            I => \N__34389\
        );

    \I__7179\ : InMux
    port map (
            O => \N__34392\,
            I => \N__34386\
        );

    \I__7178\ : Span4Mux_v
    port map (
            O => \N__34389\,
            I => \N__34383\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__34386\,
            I => data_out_frame2_17_2
        );

    \I__7176\ : Odrv4
    port map (
            O => \N__34383\,
            I => data_out_frame2_17_2
        );

    \I__7175\ : CascadeMux
    port map (
            O => \N__34378\,
            I => \c0.n17930_cascade_\
        );

    \I__7174\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34372\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__34372\,
            I => \c0.n22_adj_2358\
        );

    \I__7172\ : CascadeMux
    port map (
            O => \N__34369\,
            I => \N__34366\
        );

    \I__7171\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34363\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__34363\,
            I => \c0.n17936\
        );

    \I__7169\ : CascadeMux
    port map (
            O => \N__34360\,
            I => \c0.n17456_cascade_\
        );

    \I__7168\ : CEMux
    port map (
            O => \N__34357\,
            I => \N__34352\
        );

    \I__7167\ : CascadeMux
    port map (
            O => \N__34356\,
            I => \N__34349\
        );

    \I__7166\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34345\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__34352\,
            I => \N__34342\
        );

    \I__7164\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34339\
        );

    \I__7163\ : InMux
    port map (
            O => \N__34348\,
            I => \N__34336\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__34345\,
            I => \N__34333\
        );

    \I__7161\ : Span4Mux_s2_v
    port map (
            O => \N__34342\,
            I => \N__34330\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__34339\,
            I => \c0.n10054\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__34336\,
            I => \c0.n10054\
        );

    \I__7158\ : Odrv4
    port map (
            O => \N__34333\,
            I => \c0.n10054\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__34330\,
            I => \c0.n10054\
        );

    \I__7156\ : InMux
    port map (
            O => \N__34321\,
            I => \N__34318\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__34318\,
            I => \N__34314\
        );

    \I__7154\ : InMux
    port map (
            O => \N__34317\,
            I => \N__34311\
        );

    \I__7153\ : Span4Mux_h
    port map (
            O => \N__34314\,
            I => \N__34304\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__34311\,
            I => \N__34304\
        );

    \I__7151\ : InMux
    port map (
            O => \N__34310\,
            I => \N__34299\
        );

    \I__7150\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34299\
        );

    \I__7149\ : Span4Mux_h
    port map (
            O => \N__34304\,
            I => \N__34294\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__34299\,
            I => \N__34294\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__34294\,
            I => n9361
        );

    \I__7146\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34288\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__34288\,
            I => \N__34285\
        );

    \I__7144\ : Odrv12
    port map (
            O => \N__34285\,
            I => n17154
        );

    \I__7143\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34277\
        );

    \I__7142\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34272\
        );

    \I__7141\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34269\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34266\
        );

    \I__7139\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34263\
        );

    \I__7138\ : InMux
    port map (
            O => \N__34275\,
            I => \N__34259\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__34272\,
            I => \N__34256\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__34269\,
            I => \N__34249\
        );

    \I__7135\ : Span4Mux_v
    port map (
            O => \N__34266\,
            I => \N__34249\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__34263\,
            I => \N__34249\
        );

    \I__7133\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34243\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__34259\,
            I => \N__34238\
        );

    \I__7131\ : Span12Mux_v
    port map (
            O => \N__34256\,
            I => \N__34238\
        );

    \I__7130\ : Span4Mux_v
    port map (
            O => \N__34249\,
            I => \N__34235\
        );

    \I__7129\ : InMux
    port map (
            O => \N__34248\,
            I => \N__34228\
        );

    \I__7128\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34228\
        );

    \I__7127\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34228\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__34243\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__7125\ : Odrv12
    port map (
            O => \N__34238\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__34235\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__34228\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__7122\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34216\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__34216\,
            I => \N__34213\
        );

    \I__7120\ : Span4Mux_h
    port map (
            O => \N__34213\,
            I => \N__34210\
        );

    \I__7119\ : Odrv4
    port map (
            O => \N__34210\,
            I => \c0.tx2_transmit_N_1997\
        );

    \I__7118\ : InMux
    port map (
            O => \N__34207\,
            I => \c0.n15615\
        );

    \I__7117\ : InMux
    port map (
            O => \N__34204\,
            I => \c0.n15616\
        );

    \I__7116\ : InMux
    port map (
            O => \N__34201\,
            I => \c0.n15617\
        );

    \I__7115\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34189\
        );

    \I__7114\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34189\
        );

    \I__7113\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34186\
        );

    \I__7112\ : InMux
    port map (
            O => \N__34195\,
            I => \N__34181\
        );

    \I__7111\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34181\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__34189\,
            I => \N__34176\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__34186\,
            I => \N__34176\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__34181\,
            I => \c0.data_out_7_7\
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__34176\,
            I => \c0.data_out_7_7\
        );

    \I__7106\ : CascadeMux
    port map (
            O => \N__34171\,
            I => \c0.n5_adj_2188_cascade_\
        );

    \I__7105\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34165\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__34165\,
            I => \c0.n18041\
        );

    \I__7103\ : InMux
    port map (
            O => \N__34162\,
            I => \N__34159\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__34159\,
            I => \c0.n5_adj_2208\
        );

    \I__7101\ : CascadeMux
    port map (
            O => \N__34156\,
            I => \c0.n17543_cascade_\
        );

    \I__7100\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34150\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__34150\,
            I => \c0.n18011\
        );

    \I__7098\ : InMux
    port map (
            O => \N__34147\,
            I => \N__34144\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__34144\,
            I => \c0.n17445\
        );

    \I__7096\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34137\
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__34140\,
            I => \N__34134\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__34137\,
            I => \N__34130\
        );

    \I__7093\ : InMux
    port map (
            O => \N__34134\,
            I => \N__34127\
        );

    \I__7092\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34124\
        );

    \I__7091\ : Span4Mux_h
    port map (
            O => \N__34130\,
            I => \N__34121\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__34127\,
            I => \c0.data_out_7_5\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__34124\,
            I => \c0.data_out_7_5\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__34121\,
            I => \c0.data_out_7_5\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__34114\,
            I => \N__34111\
        );

    \I__7086\ : InMux
    port map (
            O => \N__34111\,
            I => \N__34108\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__34108\,
            I => \N__34105\
        );

    \I__7084\ : Odrv4
    port map (
            O => \N__34105\,
            I => \c0.n26\
        );

    \I__7083\ : InMux
    port map (
            O => \N__34102\,
            I => \N__34099\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__34099\,
            I => \N__34096\
        );

    \I__7081\ : Odrv12
    port map (
            O => \N__34096\,
            I => n18032
        );

    \I__7080\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34090\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__34090\,
            I => n10
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__34087\,
            I => \N__34084\
        );

    \I__7077\ : InMux
    port map (
            O => \N__34084\,
            I => \N__34081\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__34081\,
            I => \N__34078\
        );

    \I__7075\ : Odrv4
    port map (
            O => \N__34078\,
            I => \c0.n5_adj_2142\
        );

    \I__7074\ : InMux
    port map (
            O => \N__34075\,
            I => \N__34071\
        );

    \I__7073\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34068\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__34071\,
            I => \N__34065\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__34068\,
            I => data_out_3_0
        );

    \I__7070\ : Odrv4
    port map (
            O => \N__34065\,
            I => data_out_3_0
        );

    \I__7069\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34057\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__34057\,
            I => \N__34054\
        );

    \I__7067\ : Span4Mux_v
    port map (
            O => \N__34054\,
            I => \N__34050\
        );

    \I__7066\ : InMux
    port map (
            O => \N__34053\,
            I => \N__34047\
        );

    \I__7065\ : Span4Mux_h
    port map (
            O => \N__34050\,
            I => \N__34044\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__34047\,
            I => \c0.data_out_3_6\
        );

    \I__7063\ : Odrv4
    port map (
            O => \N__34044\,
            I => \c0.data_out_3_6\
        );

    \I__7062\ : CascadeMux
    port map (
            O => \N__34039\,
            I => \c0.n10054_cascade_\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34032\
        );

    \I__7060\ : InMux
    port map (
            O => \N__34035\,
            I => \N__34029\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__34032\,
            I => data_out_3_5
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__34029\,
            I => data_out_3_5
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__34024\,
            I => \N__34021\
        );

    \I__7056\ : InMux
    port map (
            O => \N__34021\,
            I => \N__34017\
        );

    \I__7055\ : InMux
    port map (
            O => \N__34020\,
            I => \N__34014\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__34017\,
            I => data_out_2_5
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__34014\,
            I => data_out_2_5
        );

    \I__7052\ : CascadeMux
    port map (
            O => \N__34009\,
            I => \N__34006\
        );

    \I__7051\ : InMux
    port map (
            O => \N__34006\,
            I => \N__34003\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__34003\,
            I => \N__34000\
        );

    \I__7049\ : Span4Mux_h
    port map (
            O => \N__34000\,
            I => \N__33997\
        );

    \I__7048\ : Span4Mux_h
    port map (
            O => \N__33997\,
            I => \N__33994\
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__33994\,
            I => \c0.n9530\
        );

    \I__7046\ : CascadeMux
    port map (
            O => \N__33991\,
            I => \N__33988\
        );

    \I__7045\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33984\
        );

    \I__7044\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33981\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__33984\,
            I => data_out_1_6
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__33981\,
            I => data_out_1_6
        );

    \I__7041\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33973\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__33973\,
            I => \N__33969\
        );

    \I__7039\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33966\
        );

    \I__7038\ : Span4Mux_h
    port map (
            O => \N__33969\,
            I => \N__33963\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__33966\,
            I => data_out_2_0
        );

    \I__7036\ : Odrv4
    port map (
            O => \N__33963\,
            I => data_out_2_0
        );

    \I__7035\ : InMux
    port map (
            O => \N__33958\,
            I => \N__33955\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__33955\,
            I => \N__33952\
        );

    \I__7033\ : Odrv12
    port map (
            O => \N__33952\,
            I => \c0.n9509\
        );

    \I__7032\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33946\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__33946\,
            I => \N__33943\
        );

    \I__7030\ : Span4Mux_h
    port map (
            O => \N__33943\,
            I => \N__33940\
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__33940\,
            I => \c0.tx2.r_Tx_Data_1\
        );

    \I__7028\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33934\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__33934\,
            I => \N__33931\
        );

    \I__7026\ : Span4Mux_v
    port map (
            O => \N__33931\,
            I => \N__33928\
        );

    \I__7025\ : Odrv4
    port map (
            O => \N__33928\,
            I => \c0.n17548\
        );

    \I__7024\ : InMux
    port map (
            O => \N__33925\,
            I => \N__33922\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__33922\,
            I => \N__33919\
        );

    \I__7022\ : Odrv12
    port map (
            O => \N__33919\,
            I => \c0.n17589\
        );

    \I__7021\ : InMux
    port map (
            O => \N__33916\,
            I => \N__33913\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__33913\,
            I => \N__33910\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__33910\,
            I => \c0.n2_adj_2298\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__33907\,
            I => \c0.n18029_cascade_\
        );

    \I__7017\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33901\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__33901\,
            I => \N__33898\
        );

    \I__7015\ : Odrv4
    port map (
            O => \N__33898\,
            I => \c0.n8_adj_2138\
        );

    \I__7014\ : CascadeMux
    port map (
            O => \N__33895\,
            I => \N__33892\
        );

    \I__7013\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33889\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__33889\,
            I => \c0.n5_adj_2299\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__33886\,
            I => \N__33882\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \N__33877\
        );

    \I__7009\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33871\
        );

    \I__7008\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33866\
        );

    \I__7007\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33866\
        );

    \I__7006\ : InMux
    port map (
            O => \N__33877\,
            I => \N__33863\
        );

    \I__7005\ : CascadeMux
    port map (
            O => \N__33876\,
            I => \N__33860\
        );

    \I__7004\ : CascadeMux
    port map (
            O => \N__33875\,
            I => \N__33855\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__33874\,
            I => \N__33852\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__33871\,
            I => \N__33849\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__33866\,
            I => \N__33844\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__33863\,
            I => \N__33844\
        );

    \I__6999\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33841\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__33859\,
            I => \N__33838\
        );

    \I__6997\ : InMux
    port map (
            O => \N__33858\,
            I => \N__33835\
        );

    \I__6996\ : InMux
    port map (
            O => \N__33855\,
            I => \N__33829\
        );

    \I__6995\ : InMux
    port map (
            O => \N__33852\,
            I => \N__33829\
        );

    \I__6994\ : Span4Mux_v
    port map (
            O => \N__33849\,
            I => \N__33822\
        );

    \I__6993\ : Span4Mux_s2_v
    port map (
            O => \N__33844\,
            I => \N__33822\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__33841\,
            I => \N__33822\
        );

    \I__6991\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33819\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__33835\,
            I => \N__33816\
        );

    \I__6989\ : InMux
    port map (
            O => \N__33834\,
            I => \N__33813\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__33829\,
            I => \N__33810\
        );

    \I__6987\ : Span4Mux_h
    port map (
            O => \N__33822\,
            I => \N__33807\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__33819\,
            I => \N__33798\
        );

    \I__6985\ : Span12Mux_s5_v
    port map (
            O => \N__33816\,
            I => \N__33798\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__33813\,
            I => \N__33798\
        );

    \I__6983\ : Span12Mux_s2_h
    port map (
            O => \N__33810\,
            I => \N__33798\
        );

    \I__6982\ : Span4Mux_h
    port map (
            O => \N__33807\,
            I => \N__33795\
        );

    \I__6981\ : Odrv12
    port map (
            O => \N__33798\,
            I => \r_SM_Main_0_adj_2441\
        );

    \I__6980\ : Odrv4
    port map (
            O => \N__33795\,
            I => \r_SM_Main_0_adj_2441\
        );

    \I__6979\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33787\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__33787\,
            I => \N__33784\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__33784\,
            I => \N__33781\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__33781\,
            I => \N__33777\
        );

    \I__6975\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33774\
        );

    \I__6974\ : Span4Mux_h
    port map (
            O => \N__33777\,
            I => \N__33771\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__33774\,
            I => \c0.rx.r_SM_Main_2_N_2096_0\
        );

    \I__6972\ : Odrv4
    port map (
            O => \N__33771\,
            I => \c0.rx.r_SM_Main_2_N_2096_0\
        );

    \I__6971\ : CascadeMux
    port map (
            O => \N__33766\,
            I => \N__33760\
        );

    \I__6970\ : CascadeMux
    port map (
            O => \N__33765\,
            I => \N__33755\
        );

    \I__6969\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33748\
        );

    \I__6968\ : InMux
    port map (
            O => \N__33763\,
            I => \N__33748\
        );

    \I__6967\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33741\
        );

    \I__6966\ : InMux
    port map (
            O => \N__33759\,
            I => \N__33741\
        );

    \I__6965\ : InMux
    port map (
            O => \N__33758\,
            I => \N__33738\
        );

    \I__6964\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33735\
        );

    \I__6963\ : InMux
    port map (
            O => \N__33754\,
            I => \N__33732\
        );

    \I__6962\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33728\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__33748\,
            I => \N__33725\
        );

    \I__6960\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33722\
        );

    \I__6959\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33719\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33716\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__33738\,
            I => \N__33713\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33710\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__33732\,
            I => \N__33707\
        );

    \I__6954\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33704\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__33728\,
            I => \N__33699\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__33725\,
            I => \N__33699\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__33722\,
            I => \N__33696\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__33719\,
            I => \N__33689\
        );

    \I__6949\ : Span4Mux_h
    port map (
            O => \N__33716\,
            I => \N__33689\
        );

    \I__6948\ : Span4Mux_v
    port map (
            O => \N__33713\,
            I => \N__33689\
        );

    \I__6947\ : Span4Mux_v
    port map (
            O => \N__33710\,
            I => \N__33684\
        );

    \I__6946\ : Span4Mux_s2_v
    port map (
            O => \N__33707\,
            I => \N__33684\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__33704\,
            I => \N__33681\
        );

    \I__6944\ : Span4Mux_v
    port map (
            O => \N__33699\,
            I => \N__33676\
        );

    \I__6943\ : Span4Mux_s2_v
    port map (
            O => \N__33696\,
            I => \N__33676\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__33689\,
            I => \N__33671\
        );

    \I__6941\ : Span4Mux_h
    port map (
            O => \N__33684\,
            I => \N__33671\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__33681\,
            I => \N__33666\
        );

    \I__6939\ : Span4Mux_h
    port map (
            O => \N__33676\,
            I => \N__33666\
        );

    \I__6938\ : Odrv4
    port map (
            O => \N__33671\,
            I => \r_Rx_Data\
        );

    \I__6937\ : Odrv4
    port map (
            O => \N__33666\,
            I => \r_Rx_Data\
        );

    \I__6936\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33658\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__33658\,
            I => n1
        );

    \I__6934\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33652\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__33652\,
            I => \N__33649\
        );

    \I__6932\ : Span4Mux_v
    port map (
            O => \N__33649\,
            I => \N__33646\
        );

    \I__6931\ : Odrv4
    port map (
            O => \N__33646\,
            I => \c0.n17915\
        );

    \I__6930\ : CascadeMux
    port map (
            O => \N__33643\,
            I => \N__33640\
        );

    \I__6929\ : InMux
    port map (
            O => \N__33640\,
            I => \N__33634\
        );

    \I__6928\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33634\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__33634\,
            I => data_out_frame2_18_1
        );

    \I__6926\ : CascadeMux
    port map (
            O => \N__33631\,
            I => \c0.n17909_cascade_\
        );

    \I__6925\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33625\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__33625\,
            I => \N__33622\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__33622\,
            I => \c0.n6\
        );

    \I__6922\ : InMux
    port map (
            O => \N__33619\,
            I => \N__33616\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__33616\,
            I => \c0.n18107\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__33613\,
            I => \N__33610\
        );

    \I__6919\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33604\
        );

    \I__6917\ : Odrv12
    port map (
            O => \N__33604\,
            I => \c0.n17579\
        );

    \I__6916\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33598\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__33598\,
            I => \c0.n17912\
        );

    \I__6914\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33592\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__33592\,
            I => \c0.n18110\
        );

    \I__6912\ : CascadeMux
    port map (
            O => \N__33589\,
            I => \c0.n22_adj_2359_cascade_\
        );

    \I__6911\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33583\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__33583\,
            I => \c0.n9758\
        );

    \I__6909\ : SRMux
    port map (
            O => \N__33580\,
            I => \N__33577\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__33577\,
            I => \N__33574\
        );

    \I__6907\ : Span4Mux_h
    port map (
            O => \N__33574\,
            I => \N__33571\
        );

    \I__6906\ : Odrv4
    port map (
            O => \N__33571\,
            I => \c0.n13496\
        );

    \I__6905\ : CascadeMux
    port map (
            O => \N__33568\,
            I => \N__33565\
        );

    \I__6904\ : InMux
    port map (
            O => \N__33565\,
            I => \N__33561\
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__33564\,
            I => \N__33558\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__33561\,
            I => \N__33553\
        );

    \I__6901\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33548\
        );

    \I__6900\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33548\
        );

    \I__6899\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33545\
        );

    \I__6898\ : Span4Mux_v
    port map (
            O => \N__33553\,
            I => \N__33538\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__33548\,
            I => \N__33538\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__33545\,
            I => \N__33538\
        );

    \I__6895\ : Odrv4
    port map (
            O => \N__33538\,
            I => data_out_frame2_7_3
        );

    \I__6894\ : InMux
    port map (
            O => \N__33535\,
            I => \N__33527\
        );

    \I__6893\ : InMux
    port map (
            O => \N__33534\,
            I => \N__33524\
        );

    \I__6892\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33518\
        );

    \I__6891\ : InMux
    port map (
            O => \N__33532\,
            I => \N__33512\
        );

    \I__6890\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33509\
        );

    \I__6889\ : InMux
    port map (
            O => \N__33530\,
            I => \N__33506\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__33527\,
            I => \N__33501\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__33524\,
            I => \N__33501\
        );

    \I__6886\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33494\
        );

    \I__6885\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33494\
        );

    \I__6884\ : InMux
    port map (
            O => \N__33521\,
            I => \N__33494\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__33518\,
            I => \N__33490\
        );

    \I__6882\ : InMux
    port map (
            O => \N__33517\,
            I => \N__33487\
        );

    \I__6881\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33482\
        );

    \I__6880\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33482\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__33512\,
            I => \N__33479\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__33509\,
            I => \N__33467\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__33506\,
            I => \N__33467\
        );

    \I__6876\ : Span4Mux_h
    port map (
            O => \N__33501\,
            I => \N__33467\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__33494\,
            I => \N__33467\
        );

    \I__6874\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33464\
        );

    \I__6873\ : Sp12to4
    port map (
            O => \N__33490\,
            I => \N__33455\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__33487\,
            I => \N__33455\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__33482\,
            I => \N__33455\
        );

    \I__6870\ : Span12Mux_v
    port map (
            O => \N__33479\,
            I => \N__33455\
        );

    \I__6869\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33450\
        );

    \I__6868\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33450\
        );

    \I__6867\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33447\
        );

    \I__6866\ : Span4Mux_v
    port map (
            O => \N__33467\,
            I => \N__33444\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__33464\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6864\ : Odrv12
    port map (
            O => \N__33455\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__33450\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__33447\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__33444\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__6860\ : CascadeMux
    port map (
            O => \N__33433\,
            I => \N__33430\
        );

    \I__6859\ : InMux
    port map (
            O => \N__33430\,
            I => \N__33426\
        );

    \I__6858\ : InMux
    port map (
            O => \N__33429\,
            I => \N__33422\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33419\
        );

    \I__6856\ : InMux
    port map (
            O => \N__33425\,
            I => \N__33416\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__33422\,
            I => \N__33413\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__33419\,
            I => \N__33409\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__33416\,
            I => \N__33406\
        );

    \I__6852\ : Span4Mux_h
    port map (
            O => \N__33413\,
            I => \N__33403\
        );

    \I__6851\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33398\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__33409\,
            I => \N__33392\
        );

    \I__6849\ : Span4Mux_v
    port map (
            O => \N__33406\,
            I => \N__33392\
        );

    \I__6848\ : Sp12to4
    port map (
            O => \N__33403\,
            I => \N__33389\
        );

    \I__6847\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33386\
        );

    \I__6846\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33383\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__33398\,
            I => \N__33380\
        );

    \I__6844\ : InMux
    port map (
            O => \N__33397\,
            I => \N__33377\
        );

    \I__6843\ : Sp12to4
    port map (
            O => \N__33392\,
            I => \N__33372\
        );

    \I__6842\ : Span12Mux_v
    port map (
            O => \N__33389\,
            I => \N__33372\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__33386\,
            I => \N__33365\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__33383\,
            I => \N__33365\
        );

    \I__6839\ : Span4Mux_v
    port map (
            O => \N__33380\,
            I => \N__33365\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__33377\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__6837\ : Odrv12
    port map (
            O => \N__33372\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__6836\ : Odrv4
    port map (
            O => \N__33365\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__6835\ : InMux
    port map (
            O => \N__33358\,
            I => \N__33353\
        );

    \I__6834\ : InMux
    port map (
            O => \N__33357\,
            I => \N__33349\
        );

    \I__6833\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33346\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__33353\,
            I => \N__33343\
        );

    \I__6831\ : InMux
    port map (
            O => \N__33352\,
            I => \N__33340\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__33349\,
            I => \N__33335\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__33346\,
            I => \N__33335\
        );

    \I__6828\ : Span4Mux_h
    port map (
            O => \N__33343\,
            I => \N__33328\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__33340\,
            I => \N__33328\
        );

    \I__6826\ : Span4Mux_v
    port map (
            O => \N__33335\,
            I => \N__33328\
        );

    \I__6825\ : Span4Mux_h
    port map (
            O => \N__33328\,
            I => \N__33325\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__33325\,
            I => \c0.n62\
        );

    \I__6823\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33316\
        );

    \I__6822\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33313\
        );

    \I__6821\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33310\
        );

    \I__6820\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33307\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__33316\,
            I => \N__33304\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__33313\,
            I => \c0.n13464\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__33310\,
            I => \c0.n13464\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__33307\,
            I => \c0.n13464\
        );

    \I__6815\ : Odrv12
    port map (
            O => \N__33304\,
            I => \c0.n13464\
        );

    \I__6814\ : CascadeMux
    port map (
            O => \N__33295\,
            I => \c0.n2_adj_2330_cascade_\
        );

    \I__6813\ : SRMux
    port map (
            O => \N__33292\,
            I => \N__33289\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__33289\,
            I => \N__33286\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__33286\,
            I => \N__33283\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__33283\,
            I => \c0.n16377\
        );

    \I__6809\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33273\
        );

    \I__6808\ : InMux
    port map (
            O => \N__33279\,
            I => \N__33270\
        );

    \I__6807\ : InMux
    port map (
            O => \N__33278\,
            I => \N__33262\
        );

    \I__6806\ : InMux
    port map (
            O => \N__33277\,
            I => \N__33251\
        );

    \I__6805\ : InMux
    port map (
            O => \N__33276\,
            I => \N__33248\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__33273\,
            I => \N__33242\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__33270\,
            I => \N__33242\
        );

    \I__6802\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33239\
        );

    \I__6801\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33236\
        );

    \I__6800\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33233\
        );

    \I__6799\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33230\
        );

    \I__6798\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33227\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__33262\,
            I => \N__33222\
        );

    \I__6796\ : InMux
    port map (
            O => \N__33261\,
            I => \N__33219\
        );

    \I__6795\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33216\
        );

    \I__6794\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33213\
        );

    \I__6793\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33210\
        );

    \I__6792\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33205\
        );

    \I__6791\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33202\
        );

    \I__6790\ : InMux
    port map (
            O => \N__33255\,
            I => \N__33199\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33254\,
            I => \N__33196\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__33251\,
            I => \N__33190\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__33248\,
            I => \N__33190\
        );

    \I__6786\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33187\
        );

    \I__6785\ : Span4Mux_v
    port map (
            O => \N__33242\,
            I => \N__33168\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__33239\,
            I => \N__33168\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__33236\,
            I => \N__33168\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__33233\,
            I => \N__33168\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__33230\,
            I => \N__33168\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__33227\,
            I => \N__33168\
        );

    \I__6779\ : InMux
    port map (
            O => \N__33226\,
            I => \N__33165\
        );

    \I__6778\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33162\
        );

    \I__6777\ : Span4Mux_v
    port map (
            O => \N__33222\,
            I => \N__33150\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__33219\,
            I => \N__33150\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__33216\,
            I => \N__33150\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__33213\,
            I => \N__33150\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__33210\,
            I => \N__33150\
        );

    \I__6772\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33147\
        );

    \I__6771\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33144\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__33205\,
            I => \N__33135\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__33202\,
            I => \N__33135\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__33199\,
            I => \N__33135\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__33196\,
            I => \N__33135\
        );

    \I__6766\ : InMux
    port map (
            O => \N__33195\,
            I => \N__33132\
        );

    \I__6765\ : Span4Mux_v
    port map (
            O => \N__33190\,
            I => \N__33127\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__33187\,
            I => \N__33127\
        );

    \I__6763\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33124\
        );

    \I__6762\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33121\
        );

    \I__6761\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33118\
        );

    \I__6760\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33115\
        );

    \I__6759\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33112\
        );

    \I__6758\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33109\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__33168\,
            I => \N__33102\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__33165\,
            I => \N__33102\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__33162\,
            I => \N__33102\
        );

    \I__6754\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33099\
        );

    \I__6753\ : Span4Mux_v
    port map (
            O => \N__33150\,
            I => \N__33094\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__33147\,
            I => \N__33091\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__33144\,
            I => \N__33088\
        );

    \I__6750\ : Span4Mux_h
    port map (
            O => \N__33135\,
            I => \N__33079\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__33132\,
            I => \N__33079\
        );

    \I__6748\ : Span4Mux_h
    port map (
            O => \N__33127\,
            I => \N__33079\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__33124\,
            I => \N__33079\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__33121\,
            I => \N__33076\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33073\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__33115\,
            I => \N__33068\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__33112\,
            I => \N__33068\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__33109\,
            I => \N__33065\
        );

    \I__6741\ : Span4Mux_v
    port map (
            O => \N__33102\,
            I => \N__33060\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__33099\,
            I => \N__33060\
        );

    \I__6739\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33057\
        );

    \I__6738\ : CascadeMux
    port map (
            O => \N__33097\,
            I => \N__33054\
        );

    \I__6737\ : Span4Mux_h
    port map (
            O => \N__33094\,
            I => \N__33048\
        );

    \I__6736\ : Span4Mux_v
    port map (
            O => \N__33091\,
            I => \N__33048\
        );

    \I__6735\ : Span12Mux_h
    port map (
            O => \N__33088\,
            I => \N__33045\
        );

    \I__6734\ : Span4Mux_v
    port map (
            O => \N__33079\,
            I => \N__33040\
        );

    \I__6733\ : Span4Mux_v
    port map (
            O => \N__33076\,
            I => \N__33040\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__33073\,
            I => \N__33037\
        );

    \I__6731\ : Span4Mux_v
    port map (
            O => \N__33068\,
            I => \N__33030\
        );

    \I__6730\ : Span4Mux_h
    port map (
            O => \N__33065\,
            I => \N__33030\
        );

    \I__6729\ : Span4Mux_h
    port map (
            O => \N__33060\,
            I => \N__33030\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__33057\,
            I => \N__33027\
        );

    \I__6727\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33022\
        );

    \I__6726\ : InMux
    port map (
            O => \N__33053\,
            I => \N__33022\
        );

    \I__6725\ : Odrv4
    port map (
            O => \N__33048\,
            I => n9452
        );

    \I__6724\ : Odrv12
    port map (
            O => \N__33045\,
            I => n9452
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__33040\,
            I => n9452
        );

    \I__6722\ : Odrv4
    port map (
            O => \N__33037\,
            I => n9452
        );

    \I__6721\ : Odrv4
    port map (
            O => \N__33030\,
            I => n9452
        );

    \I__6720\ : Odrv12
    port map (
            O => \N__33027\,
            I => n9452
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__33022\,
            I => n9452
        );

    \I__6718\ : InMux
    port map (
            O => \N__33007\,
            I => \N__32993\
        );

    \I__6717\ : InMux
    port map (
            O => \N__33006\,
            I => \N__32990\
        );

    \I__6716\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32985\
        );

    \I__6715\ : InMux
    port map (
            O => \N__33004\,
            I => \N__32982\
        );

    \I__6714\ : InMux
    port map (
            O => \N__33003\,
            I => \N__32979\
        );

    \I__6713\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32976\
        );

    \I__6712\ : InMux
    port map (
            O => \N__33001\,
            I => \N__32973\
        );

    \I__6711\ : InMux
    port map (
            O => \N__33000\,
            I => \N__32970\
        );

    \I__6710\ : InMux
    port map (
            O => \N__32999\,
            I => \N__32967\
        );

    \I__6709\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32964\
        );

    \I__6708\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32961\
        );

    \I__6707\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32956\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__32993\,
            I => \N__32951\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__32990\,
            I => \N__32951\
        );

    \I__6704\ : InMux
    port map (
            O => \N__32989\,
            I => \N__32948\
        );

    \I__6703\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32943\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__32985\,
            I => \N__32938\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__32982\,
            I => \N__32938\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__32979\,
            I => \N__32935\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__32976\,
            I => \N__32922\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__32973\,
            I => \N__32922\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__32970\,
            I => \N__32922\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__32967\,
            I => \N__32922\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__32964\,
            I => \N__32922\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__32961\,
            I => \N__32922\
        );

    \I__6693\ : InMux
    port map (
            O => \N__32960\,
            I => \N__32919\
        );

    \I__6692\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32915\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__32956\,
            I => \N__32903\
        );

    \I__6690\ : Span4Mux_v
    port map (
            O => \N__32951\,
            I => \N__32903\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__32948\,
            I => \N__32903\
        );

    \I__6688\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32900\
        );

    \I__6687\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32897\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__32943\,
            I => \N__32889\
        );

    \I__6685\ : Span4Mux_v
    port map (
            O => \N__32938\,
            I => \N__32880\
        );

    \I__6684\ : Span4Mux_s1_h
    port map (
            O => \N__32935\,
            I => \N__32880\
        );

    \I__6683\ : Span4Mux_v
    port map (
            O => \N__32922\,
            I => \N__32880\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__32919\,
            I => \N__32880\
        );

    \I__6681\ : InMux
    port map (
            O => \N__32918\,
            I => \N__32877\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__32915\,
            I => \N__32874\
        );

    \I__6679\ : InMux
    port map (
            O => \N__32914\,
            I => \N__32871\
        );

    \I__6678\ : InMux
    port map (
            O => \N__32913\,
            I => \N__32868\
        );

    \I__6677\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32865\
        );

    \I__6676\ : InMux
    port map (
            O => \N__32911\,
            I => \N__32862\
        );

    \I__6675\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32859\
        );

    \I__6674\ : Span4Mux_h
    port map (
            O => \N__32903\,
            I => \N__32852\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__32900\,
            I => \N__32852\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__32897\,
            I => \N__32852\
        );

    \I__6671\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32849\
        );

    \I__6670\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32842\
        );

    \I__6669\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32842\
        );

    \I__6668\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32839\
        );

    \I__6667\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32836\
        );

    \I__6666\ : Span4Mux_v
    port map (
            O => \N__32889\,
            I => \N__32827\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__32880\,
            I => \N__32827\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__32877\,
            I => \N__32827\
        );

    \I__6663\ : Span4Mux_v
    port map (
            O => \N__32874\,
            I => \N__32823\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__32871\,
            I => \N__32816\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__32868\,
            I => \N__32816\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32816\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__32862\,
            I => \N__32807\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__32859\,
            I => \N__32807\
        );

    \I__6657\ : Span4Mux_v
    port map (
            O => \N__32852\,
            I => \N__32807\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__32849\,
            I => \N__32807\
        );

    \I__6655\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32804\
        );

    \I__6654\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32799\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__32842\,
            I => \N__32796\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__32839\,
            I => \N__32791\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__32836\,
            I => \N__32791\
        );

    \I__6650\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32787\
        );

    \I__6649\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32784\
        );

    \I__6648\ : Span4Mux_h
    port map (
            O => \N__32827\,
            I => \N__32780\
        );

    \I__6647\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32777\
        );

    \I__6646\ : Span4Mux_h
    port map (
            O => \N__32823\,
            I => \N__32768\
        );

    \I__6645\ : Span4Mux_v
    port map (
            O => \N__32816\,
            I => \N__32768\
        );

    \I__6644\ : Span4Mux_s3_h
    port map (
            O => \N__32807\,
            I => \N__32768\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__32804\,
            I => \N__32768\
        );

    \I__6642\ : InMux
    port map (
            O => \N__32803\,
            I => \N__32765\
        );

    \I__6641\ : InMux
    port map (
            O => \N__32802\,
            I => \N__32762\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__32799\,
            I => \N__32755\
        );

    \I__6639\ : Span4Mux_v
    port map (
            O => \N__32796\,
            I => \N__32755\
        );

    \I__6638\ : Span4Mux_h
    port map (
            O => \N__32791\,
            I => \N__32755\
        );

    \I__6637\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32752\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__32787\,
            I => \N__32747\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__32784\,
            I => \N__32747\
        );

    \I__6634\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32744\
        );

    \I__6633\ : Odrv4
    port map (
            O => \N__32780\,
            I => n12933
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__32777\,
            I => n12933
        );

    \I__6631\ : Odrv4
    port map (
            O => \N__32768\,
            I => n12933
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__32765\,
            I => n12933
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__32762\,
            I => n12933
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__32755\,
            I => n12933
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__32752\,
            I => n12933
        );

    \I__6626\ : Odrv12
    port map (
            O => \N__32747\,
            I => n12933
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__32744\,
            I => n12933
        );

    \I__6624\ : InMux
    port map (
            O => \N__32725\,
            I => \N__32722\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__32722\,
            I => \N__32719\
        );

    \I__6622\ : Span4Mux_h
    port map (
            O => \N__32719\,
            I => \N__32716\
        );

    \I__6621\ : Span4Mux_h
    port map (
            O => \N__32716\,
            I => \N__32713\
        );

    \I__6620\ : Odrv4
    port map (
            O => \N__32713\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_0\
        );

    \I__6619\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32706\
        );

    \I__6618\ : CascadeMux
    port map (
            O => \N__32709\,
            I => \N__32701\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__32706\,
            I => \N__32698\
        );

    \I__6616\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32695\
        );

    \I__6615\ : InMux
    port map (
            O => \N__32704\,
            I => \N__32692\
        );

    \I__6614\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32687\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__32698\,
            I => \N__32682\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__32695\,
            I => \N__32682\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__32692\,
            I => \N__32679\
        );

    \I__6610\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32676\
        );

    \I__6609\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32673\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__32687\,
            I => \N__32670\
        );

    \I__6607\ : Span4Mux_v
    port map (
            O => \N__32682\,
            I => \N__32666\
        );

    \I__6606\ : Span4Mux_v
    port map (
            O => \N__32679\,
            I => \N__32659\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__32676\,
            I => \N__32659\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__32673\,
            I => \N__32659\
        );

    \I__6603\ : Span4Mux_v
    port map (
            O => \N__32670\,
            I => \N__32656\
        );

    \I__6602\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32653\
        );

    \I__6601\ : Sp12to4
    port map (
            O => \N__32666\,
            I => \N__32650\
        );

    \I__6600\ : Span4Mux_v
    port map (
            O => \N__32659\,
            I => \N__32645\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__32656\,
            I => \N__32645\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__32653\,
            I => \N__32642\
        );

    \I__6597\ : Span12Mux_s10_h
    port map (
            O => \N__32650\,
            I => \N__32639\
        );

    \I__6596\ : Span4Mux_h
    port map (
            O => \N__32645\,
            I => \N__32636\
        );

    \I__6595\ : Span4Mux_h
    port map (
            O => \N__32642\,
            I => \N__32633\
        );

    \I__6594\ : Odrv12
    port map (
            O => \N__32639\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__6593\ : Odrv4
    port map (
            O => \N__32636\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__32633\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__6591\ : SRMux
    port map (
            O => \N__32626\,
            I => \N__32623\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__32623\,
            I => \N__32620\
        );

    \I__6589\ : Span4Mux_v
    port map (
            O => \N__32620\,
            I => \N__32617\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__32617\,
            I => \c0.n3\
        );

    \I__6587\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32611\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__32611\,
            I => \N__32606\
        );

    \I__6585\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32603\
        );

    \I__6584\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32600\
        );

    \I__6583\ : Span4Mux_h
    port map (
            O => \N__32606\,
            I => \N__32597\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__32603\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__32600\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__6580\ : Odrv4
    port map (
            O => \N__32597\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__6579\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32585\
        );

    \I__6578\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32578\
        );

    \I__6577\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32578\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__32585\,
            I => \N__32575\
        );

    \I__6575\ : CascadeMux
    port map (
            O => \N__32584\,
            I => \N__32572\
        );

    \I__6574\ : CascadeMux
    port map (
            O => \N__32583\,
            I => \N__32568\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__32578\,
            I => \N__32563\
        );

    \I__6572\ : Span4Mux_h
    port map (
            O => \N__32575\,
            I => \N__32560\
        );

    \I__6571\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32549\
        );

    \I__6570\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32549\
        );

    \I__6569\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32549\
        );

    \I__6568\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32549\
        );

    \I__6567\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32549\
        );

    \I__6566\ : Odrv12
    port map (
            O => \N__32563\,
            I => \c0.n4_adj_2360\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__32560\,
            I => \c0.n4_adj_2360\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__32549\,
            I => \c0.n4_adj_2360\
        );

    \I__6563\ : SRMux
    port map (
            O => \N__32542\,
            I => \N__32539\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__32539\,
            I => \N__32536\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__32536\,
            I => \N__32533\
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__32533\,
            I => \c0.n16449\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__32530\,
            I => \N__32526\
        );

    \I__6558\ : InMux
    port map (
            O => \N__32529\,
            I => \N__32523\
        );

    \I__6557\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32520\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__32523\,
            I => data_out_frame2_18_2
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__32520\,
            I => data_out_frame2_18_2
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__32515\,
            I => \c0.n18119_cascade_\
        );

    \I__6553\ : CascadeMux
    port map (
            O => \N__32512\,
            I => \c0.n18122_cascade_\
        );

    \I__6552\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32506\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__32506\,
            I => \N__32503\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__32503\,
            I => \N__32500\
        );

    \I__6549\ : Span4Mux_v
    port map (
            O => \N__32500\,
            I => \N__32497\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__32497\,
            I => \c0.tx2.r_Tx_Data_2\
        );

    \I__6547\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32491\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__32491\,
            I => \N__32488\
        );

    \I__6545\ : Odrv4
    port map (
            O => \N__32488\,
            I => \c0.n17340\
        );

    \I__6544\ : InMux
    port map (
            O => \N__32485\,
            I => \N__32482\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__32482\,
            I => \c0.n2_adj_2137\
        );

    \I__6542\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32475\
        );

    \I__6541\ : InMux
    port map (
            O => \N__32478\,
            I => \N__32472\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__32475\,
            I => \c0.data_out_1_4\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__32472\,
            I => \c0.data_out_1_4\
        );

    \I__6538\ : InMux
    port map (
            O => \N__32467\,
            I => \N__32464\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__32464\,
            I => \N__32461\
        );

    \I__6536\ : Odrv12
    port map (
            O => \N__32461\,
            I => n16776
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__32458\,
            I => \N__32455\
        );

    \I__6534\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32451\
        );

    \I__6533\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32448\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__32451\,
            I => \N__32444\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32441\
        );

    \I__6530\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32438\
        );

    \I__6529\ : Span4Mux_v
    port map (
            O => \N__32444\,
            I => \N__32435\
        );

    \I__6528\ : Span4Mux_v
    port map (
            O => \N__32441\,
            I => \N__32432\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__32438\,
            I => \N__32429\
        );

    \I__6526\ : Span4Mux_h
    port map (
            O => \N__32435\,
            I => \N__32424\
        );

    \I__6525\ : Span4Mux_s2_h
    port map (
            O => \N__32432\,
            I => \N__32424\
        );

    \I__6524\ : Odrv4
    port map (
            O => \N__32429\,
            I => n17208
        );

    \I__6523\ : Odrv4
    port map (
            O => \N__32424\,
            I => n17208
        );

    \I__6522\ : InMux
    port map (
            O => \N__32419\,
            I => \N__32416\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__32416\,
            I => \N__32413\
        );

    \I__6520\ : Span4Mux_v
    port map (
            O => \N__32413\,
            I => \N__32410\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__32410\,
            I => \N__32407\
        );

    \I__6518\ : Odrv4
    port map (
            O => \N__32407\,
            I => n8828
        );

    \I__6517\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32398\
        );

    \I__6516\ : InMux
    port map (
            O => \N__32403\,
            I => \N__32398\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__32398\,
            I => \N__32393\
        );

    \I__6514\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32390\
        );

    \I__6513\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32386\
        );

    \I__6512\ : Span4Mux_h
    port map (
            O => \N__32393\,
            I => \N__32383\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__32390\,
            I => \N__32380\
        );

    \I__6510\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32377\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__32386\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__6508\ : Odrv4
    port map (
            O => \N__32383\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__6507\ : Odrv12
    port map (
            O => \N__32380\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__32377\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__6505\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32364\
        );

    \I__6504\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32361\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__32364\,
            I => \N__32358\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__32361\,
            I => \N__32355\
        );

    \I__6501\ : Span4Mux_v
    port map (
            O => \N__32358\,
            I => \N__32352\
        );

    \I__6500\ : Span4Mux_h
    port map (
            O => \N__32355\,
            I => \N__32349\
        );

    \I__6499\ : Span4Mux_h
    port map (
            O => \N__32352\,
            I => \N__32344\
        );

    \I__6498\ : Span4Mux_v
    port map (
            O => \N__32349\,
            I => \N__32344\
        );

    \I__6497\ : Odrv4
    port map (
            O => \N__32344\,
            I => \c0.n47\
        );

    \I__6496\ : CascadeMux
    port map (
            O => \N__32341\,
            I => \N__32338\
        );

    \I__6495\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32335\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__32335\,
            I => \N__32332\
        );

    \I__6493\ : Span12Mux_s10_h
    port map (
            O => \N__32332\,
            I => \N__32329\
        );

    \I__6492\ : Odrv12
    port map (
            O => \N__32329\,
            I => \c0.n6_adj_2140\
        );

    \I__6491\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32319\
        );

    \I__6490\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32319\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__32324\,
            I => \N__32314\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__32319\,
            I => \N__32311\
        );

    \I__6487\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32307\
        );

    \I__6486\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32303\
        );

    \I__6485\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32300\
        );

    \I__6484\ : Span4Mux_v
    port map (
            O => \N__32311\,
            I => \N__32296\
        );

    \I__6483\ : InMux
    port map (
            O => \N__32310\,
            I => \N__32293\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__32307\,
            I => \N__32289\
        );

    \I__6481\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32286\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__32303\,
            I => \N__32283\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__32300\,
            I => \N__32280\
        );

    \I__6478\ : InMux
    port map (
            O => \N__32299\,
            I => \N__32277\
        );

    \I__6477\ : Span4Mux_h
    port map (
            O => \N__32296\,
            I => \N__32272\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__32293\,
            I => \N__32272\
        );

    \I__6475\ : InMux
    port map (
            O => \N__32292\,
            I => \N__32269\
        );

    \I__6474\ : Span4Mux_v
    port map (
            O => \N__32289\,
            I => \N__32265\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__32286\,
            I => \N__32262\
        );

    \I__6472\ : Span4Mux_h
    port map (
            O => \N__32283\,
            I => \N__32253\
        );

    \I__6471\ : Span4Mux_v
    port map (
            O => \N__32280\,
            I => \N__32253\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__32277\,
            I => \N__32253\
        );

    \I__6469\ : Span4Mux_v
    port map (
            O => \N__32272\,
            I => \N__32248\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__32269\,
            I => \N__32248\
        );

    \I__6467\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32245\
        );

    \I__6466\ : Span4Mux_h
    port map (
            O => \N__32265\,
            I => \N__32240\
        );

    \I__6465\ : Span4Mux_v
    port map (
            O => \N__32262\,
            I => \N__32240\
        );

    \I__6464\ : InMux
    port map (
            O => \N__32261\,
            I => \N__32235\
        );

    \I__6463\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32235\
        );

    \I__6462\ : Span4Mux_h
    port map (
            O => \N__32253\,
            I => \N__32232\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__32248\,
            I => \N__32229\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__32245\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__6459\ : Odrv4
    port map (
            O => \N__32240\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__32235\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__6457\ : Odrv4
    port map (
            O => \N__32232\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__6456\ : Odrv4
    port map (
            O => \N__32229\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__6455\ : InMux
    port map (
            O => \N__32218\,
            I => \N__32215\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__32215\,
            I => \N__32212\
        );

    \I__6453\ : Span4Mux_v
    port map (
            O => \N__32212\,
            I => \N__32209\
        );

    \I__6452\ : Odrv4
    port map (
            O => \N__32209\,
            I => \c0.n5_adj_2339\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__32206\,
            I => \c0.n16814_cascade_\
        );

    \I__6450\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32200\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__32200\,
            I => \N__32197\
        );

    \I__6448\ : Odrv4
    port map (
            O => \N__32197\,
            I => \c0.tx2.n89\
        );

    \I__6447\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32187\
        );

    \I__6446\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32182\
        );

    \I__6445\ : InMux
    port map (
            O => \N__32192\,
            I => \N__32182\
        );

    \I__6444\ : InMux
    port map (
            O => \N__32191\,
            I => \N__32177\
        );

    \I__6443\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32177\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__32187\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__32182\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__32177\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__6439\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32166\
        );

    \I__6438\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32163\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__32166\,
            I => \r_Tx_Data_7\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__32163\,
            I => \r_Tx_Data_7\
        );

    \I__6435\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32155\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__32155\,
            I => \c0.n18014\
        );

    \I__6433\ : CascadeMux
    port map (
            O => \N__32152\,
            I => \N__32149\
        );

    \I__6432\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32146\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__32146\,
            I => \N__32143\
        );

    \I__6430\ : Span4Mux_v
    port map (
            O => \N__32143\,
            I => \N__32140\
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__32140\,
            I => \c0.n17585\
        );

    \I__6428\ : InMux
    port map (
            O => \N__32137\,
            I => \N__32134\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__32134\,
            I => n10_adj_2423
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__32131\,
            I => \n18044_cascade_\
        );

    \I__6425\ : InMux
    port map (
            O => \N__32128\,
            I => \N__32125\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__32125\,
            I => n10_adj_2414
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__32122\,
            I => \N__32118\
        );

    \I__6422\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32115\
        );

    \I__6421\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32112\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__32115\,
            I => data_out_0_1
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__32112\,
            I => data_out_0_1
        );

    \I__6418\ : InMux
    port map (
            O => \N__32107\,
            I => \N__32104\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__32104\,
            I => \N__32101\
        );

    \I__6416\ : Odrv4
    port map (
            O => \N__32101\,
            I => \c0.n18080\
        );

    \I__6415\ : InMux
    port map (
            O => \N__32098\,
            I => \N__32094\
        );

    \I__6414\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32091\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__32094\,
            I => data_out_3_7
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__32091\,
            I => data_out_3_7
        );

    \I__6411\ : CascadeMux
    port map (
            O => \N__32086\,
            I => \c0.n29_cascade_\
        );

    \I__6410\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32079\
        );

    \I__6409\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32076\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__32079\,
            I => \N__32073\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__32076\,
            I => \r_Tx_Data_1\
        );

    \I__6406\ : Odrv12
    port map (
            O => \N__32073\,
            I => \r_Tx_Data_1\
        );

    \I__6405\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32062\
        );

    \I__6404\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32062\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__32062\,
            I => \r_Tx_Data_5\
        );

    \I__6402\ : InMux
    port map (
            O => \N__32059\,
            I => \N__32056\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__32056\,
            I => \N__32052\
        );

    \I__6400\ : InMux
    port map (
            O => \N__32055\,
            I => \N__32049\
        );

    \I__6399\ : Span4Mux_h
    port map (
            O => \N__32052\,
            I => \N__32046\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__32049\,
            I => \c0.data_out_0_6\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__32046\,
            I => \c0.data_out_0_6\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__32041\,
            I => \c0.n9_adj_2143_cascade_\
        );

    \I__6395\ : InMux
    port map (
            O => \N__32038\,
            I => \N__32035\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__32035\,
            I => \c0.n23\
        );

    \I__6393\ : InMux
    port map (
            O => \N__32032\,
            I => \N__32029\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__32029\,
            I => \N__32026\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__32026\,
            I => \N__32023\
        );

    \I__6390\ : Odrv4
    port map (
            O => \N__32023\,
            I => \c0.n17547\
        );

    \I__6389\ : CascadeMux
    port map (
            O => \N__32020\,
            I => \c0.n5_adj_2326_cascade_\
        );

    \I__6388\ : InMux
    port map (
            O => \N__32017\,
            I => \N__32014\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__32014\,
            I => \N__32011\
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__32011\,
            I => \c0.n18023\
        );

    \I__6385\ : InMux
    port map (
            O => \N__32008\,
            I => \N__32002\
        );

    \I__6384\ : InMux
    port map (
            O => \N__32007\,
            I => \N__32002\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__32002\,
            I => \N__31985\
        );

    \I__6382\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31976\
        );

    \I__6381\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31976\
        );

    \I__6380\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31976\
        );

    \I__6379\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31976\
        );

    \I__6378\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31967\
        );

    \I__6377\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31967\
        );

    \I__6376\ : InMux
    port map (
            O => \N__31995\,
            I => \N__31967\
        );

    \I__6375\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31967\
        );

    \I__6374\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31964\
        );

    \I__6373\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31961\
        );

    \I__6372\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31956\
        );

    \I__6371\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31956\
        );

    \I__6370\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31951\
        );

    \I__6369\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31951\
        );

    \I__6368\ : Odrv12
    port map (
            O => \N__31985\,
            I => \c0.n16891\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__31976\,
            I => \c0.n16891\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__31967\,
            I => \c0.n16891\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__31964\,
            I => \c0.n16891\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__31961\,
            I => \c0.n16891\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__31956\,
            I => \c0.n16891\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__31951\,
            I => \c0.n16891\
        );

    \I__6361\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31926\
        );

    \I__6360\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31926\
        );

    \I__6359\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31926\
        );

    \I__6358\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31914\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__31926\,
            I => \N__31911\
        );

    \I__6356\ : InMux
    port map (
            O => \N__31925\,
            I => \N__31908\
        );

    \I__6355\ : InMux
    port map (
            O => \N__31924\,
            I => \N__31905\
        );

    \I__6354\ : InMux
    port map (
            O => \N__31923\,
            I => \N__31896\
        );

    \I__6353\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31896\
        );

    \I__6352\ : InMux
    port map (
            O => \N__31921\,
            I => \N__31896\
        );

    \I__6351\ : InMux
    port map (
            O => \N__31920\,
            I => \N__31896\
        );

    \I__6350\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31893\
        );

    \I__6349\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31888\
        );

    \I__6348\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31888\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__31914\,
            I => \N__31885\
        );

    \I__6346\ : Span4Mux_h
    port map (
            O => \N__31911\,
            I => \N__31880\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31880\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__31905\,
            I => \N__31874\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__31896\,
            I => \N__31867\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__31893\,
            I => \N__31867\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__31888\,
            I => \N__31867\
        );

    \I__6340\ : Span4Mux_v
    port map (
            O => \N__31885\,
            I => \N__31864\
        );

    \I__6339\ : Sp12to4
    port map (
            O => \N__31880\,
            I => \N__31861\
        );

    \I__6338\ : InMux
    port map (
            O => \N__31879\,
            I => \N__31856\
        );

    \I__6337\ : InMux
    port map (
            O => \N__31878\,
            I => \N__31856\
        );

    \I__6336\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31853\
        );

    \I__6335\ : Span4Mux_v
    port map (
            O => \N__31874\,
            I => \N__31848\
        );

    \I__6334\ : Span4Mux_v
    port map (
            O => \N__31867\,
            I => \N__31848\
        );

    \I__6333\ : Sp12to4
    port map (
            O => \N__31864\,
            I => \N__31839\
        );

    \I__6332\ : Span12Mux_v
    port map (
            O => \N__31861\,
            I => \N__31839\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__31856\,
            I => \N__31839\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__31853\,
            I => \N__31839\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__31848\,
            I => \c0.n8\
        );

    \I__6328\ : Odrv12
    port map (
            O => \N__31839\,
            I => \c0.n8\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__31834\,
            I => \N__31831\
        );

    \I__6326\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31827\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__31830\,
            I => \N__31823\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__31827\,
            I => \N__31820\
        );

    \I__6323\ : CascadeMux
    port map (
            O => \N__31826\,
            I => \N__31816\
        );

    \I__6322\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31813\
        );

    \I__6321\ : Span4Mux_h
    port map (
            O => \N__31820\,
            I => \N__31809\
        );

    \I__6320\ : InMux
    port map (
            O => \N__31819\,
            I => \N__31804\
        );

    \I__6319\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31804\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__31813\,
            I => \N__31801\
        );

    \I__6317\ : InMux
    port map (
            O => \N__31812\,
            I => \N__31798\
        );

    \I__6316\ : Span4Mux_h
    port map (
            O => \N__31809\,
            I => \N__31789\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__31804\,
            I => \N__31789\
        );

    \I__6314\ : Sp12to4
    port map (
            O => \N__31801\,
            I => \N__31784\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__31798\,
            I => \N__31784\
        );

    \I__6312\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31781\
        );

    \I__6311\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31778\
        );

    \I__6310\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31775\
        );

    \I__6309\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31772\
        );

    \I__6308\ : Odrv4
    port map (
            O => \N__31789\,
            I => rx_data_4
        );

    \I__6307\ : Odrv12
    port map (
            O => \N__31784\,
            I => rx_data_4
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__31781\,
            I => rx_data_4
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__31778\,
            I => rx_data_4
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__31775\,
            I => rx_data_4
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__31772\,
            I => rx_data_4
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__31759\,
            I => \N__31755\
        );

    \I__6301\ : InMux
    port map (
            O => \N__31758\,
            I => \N__31752\
        );

    \I__6300\ : InMux
    port map (
            O => \N__31755\,
            I => \N__31749\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__31752\,
            I => \N__31744\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__31749\,
            I => \N__31744\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__31744\,
            I => \c0.data_in_frame_2_4\
        );

    \I__6296\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31738\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__31738\,
            I => \N__31732\
        );

    \I__6294\ : CascadeMux
    port map (
            O => \N__31737\,
            I => \N__31729\
        );

    \I__6293\ : InMux
    port map (
            O => \N__31736\,
            I => \N__31725\
        );

    \I__6292\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31722\
        );

    \I__6291\ : Span4Mux_v
    port map (
            O => \N__31732\,
            I => \N__31718\
        );

    \I__6290\ : InMux
    port map (
            O => \N__31729\,
            I => \N__31715\
        );

    \I__6289\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31712\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__31725\,
            I => \N__31707\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__31722\,
            I => \N__31707\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__31721\,
            I => \N__31703\
        );

    \I__6285\ : Span4Mux_h
    port map (
            O => \N__31718\,
            I => \N__31698\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__31715\,
            I => \N__31698\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__31712\,
            I => \N__31695\
        );

    \I__6282\ : Span4Mux_h
    port map (
            O => \N__31707\,
            I => \N__31692\
        );

    \I__6281\ : InMux
    port map (
            O => \N__31706\,
            I => \N__31687\
        );

    \I__6280\ : InMux
    port map (
            O => \N__31703\,
            I => \N__31687\
        );

    \I__6279\ : Span4Mux_h
    port map (
            O => \N__31698\,
            I => \N__31684\
        );

    \I__6278\ : Span12Mux_v
    port map (
            O => \N__31695\,
            I => \N__31681\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__31692\,
            I => \c0.r_SM_Main_2_N_2036_0\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__31687\,
            I => \c0.r_SM_Main_2_N_2036_0\
        );

    \I__6275\ : Odrv4
    port map (
            O => \N__31684\,
            I => \c0.r_SM_Main_2_N_2036_0\
        );

    \I__6274\ : Odrv12
    port map (
            O => \N__31681\,
            I => \c0.r_SM_Main_2_N_2036_0\
        );

    \I__6273\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31667\
        );

    \I__6272\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31664\
        );

    \I__6271\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31661\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__31667\,
            I => \N__31657\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__31664\,
            I => \N__31654\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__31661\,
            I => \N__31651\
        );

    \I__6267\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31648\
        );

    \I__6266\ : Span4Mux_v
    port map (
            O => \N__31657\,
            I => \N__31645\
        );

    \I__6265\ : Span4Mux_h
    port map (
            O => \N__31654\,
            I => \N__31639\
        );

    \I__6264\ : Span4Mux_h
    port map (
            O => \N__31651\,
            I => \N__31636\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__31648\,
            I => \N__31633\
        );

    \I__6262\ : Span4Mux_h
    port map (
            O => \N__31645\,
            I => \N__31630\
        );

    \I__6261\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31623\
        );

    \I__6260\ : InMux
    port map (
            O => \N__31643\,
            I => \N__31623\
        );

    \I__6259\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31623\
        );

    \I__6258\ : Odrv4
    port map (
            O => \N__31639\,
            I => tx_active
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__31636\,
            I => tx_active
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__31633\,
            I => tx_active
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__31630\,
            I => tx_active
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__31623\,
            I => tx_active
        );

    \I__6253\ : CascadeMux
    port map (
            O => \N__31612\,
            I => \N__31609\
        );

    \I__6252\ : InMux
    port map (
            O => \N__31609\,
            I => \N__31605\
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__31608\,
            I => \N__31602\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31598\
        );

    \I__6249\ : InMux
    port map (
            O => \N__31602\,
            I => \N__31595\
        );

    \I__6248\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31592\
        );

    \I__6247\ : Span4Mux_s2_v
    port map (
            O => \N__31598\,
            I => \N__31589\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__31595\,
            I => \N__31584\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__31592\,
            I => \N__31584\
        );

    \I__6244\ : Span4Mux_h
    port map (
            O => \N__31589\,
            I => \N__31579\
        );

    \I__6243\ : Span4Mux_s2_v
    port map (
            O => \N__31584\,
            I => \N__31579\
        );

    \I__6242\ : Span4Mux_h
    port map (
            O => \N__31579\,
            I => \N__31576\
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__31576\,
            I => n17230
        );

    \I__6240\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31567\
        );

    \I__6239\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31567\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__31567\,
            I => data_out_1_7
        );

    \I__6237\ : InMux
    port map (
            O => \N__31564\,
            I => \N__31561\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__31561\,
            I => \N__31558\
        );

    \I__6235\ : Span4Mux_h
    port map (
            O => \N__31558\,
            I => \N__31555\
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__31555\,
            I => \c0.n10\
        );

    \I__6233\ : InMux
    port map (
            O => \N__31552\,
            I => \N__31547\
        );

    \I__6232\ : InMux
    port map (
            O => \N__31551\,
            I => \N__31542\
        );

    \I__6231\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31539\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__31547\,
            I => \N__31536\
        );

    \I__6229\ : CascadeMux
    port map (
            O => \N__31546\,
            I => \N__31533\
        );

    \I__6228\ : InMux
    port map (
            O => \N__31545\,
            I => \N__31529\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__31542\,
            I => \N__31526\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__31539\,
            I => \N__31521\
        );

    \I__6225\ : Span4Mux_v
    port map (
            O => \N__31536\,
            I => \N__31518\
        );

    \I__6224\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31515\
        );

    \I__6223\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31510\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31505\
        );

    \I__6221\ : Span4Mux_v
    port map (
            O => \N__31526\,
            I => \N__31505\
        );

    \I__6220\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31500\
        );

    \I__6219\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31500\
        );

    \I__6218\ : Span4Mux_v
    port map (
            O => \N__31521\,
            I => \N__31489\
        );

    \I__6217\ : Span4Mux_h
    port map (
            O => \N__31518\,
            I => \N__31489\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__31515\,
            I => \N__31489\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__31514\,
            I => \N__31482\
        );

    \I__6214\ : InMux
    port map (
            O => \N__31513\,
            I => \N__31478\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__31510\,
            I => \N__31475\
        );

    \I__6212\ : Span4Mux_h
    port map (
            O => \N__31505\,
            I => \N__31470\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__31500\,
            I => \N__31470\
        );

    \I__6210\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31467\
        );

    \I__6209\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31462\
        );

    \I__6208\ : InMux
    port map (
            O => \N__31497\,
            I => \N__31462\
        );

    \I__6207\ : InMux
    port map (
            O => \N__31496\,
            I => \N__31459\
        );

    \I__6206\ : Span4Mux_h
    port map (
            O => \N__31489\,
            I => \N__31456\
        );

    \I__6205\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31449\
        );

    \I__6204\ : InMux
    port map (
            O => \N__31487\,
            I => \N__31449\
        );

    \I__6203\ : InMux
    port map (
            O => \N__31486\,
            I => \N__31449\
        );

    \I__6202\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31442\
        );

    \I__6201\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31442\
        );

    \I__6200\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31442\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__31478\,
            I => \N__31435\
        );

    \I__6198\ : Span4Mux_s1_h
    port map (
            O => \N__31475\,
            I => \N__31435\
        );

    \I__6197\ : Span4Mux_h
    port map (
            O => \N__31470\,
            I => \N__31435\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__31467\,
            I => \r_SM_Main_2_adj_2443\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__31462\,
            I => \r_SM_Main_2_adj_2443\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__31459\,
            I => \r_SM_Main_2_adj_2443\
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__31456\,
            I => \r_SM_Main_2_adj_2443\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__31449\,
            I => \r_SM_Main_2_adj_2443\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__31442\,
            I => \r_SM_Main_2_adj_2443\
        );

    \I__6190\ : Odrv4
    port map (
            O => \N__31435\,
            I => \r_SM_Main_2_adj_2443\
        );

    \I__6189\ : InMux
    port map (
            O => \N__31420\,
            I => \N__31417\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__31417\,
            I => \N__31414\
        );

    \I__6187\ : Span12Mux_h
    port map (
            O => \N__31414\,
            I => \N__31411\
        );

    \I__6186\ : Odrv12
    port map (
            O => \N__31411\,
            I => n17544
        );

    \I__6185\ : CascadeMux
    port map (
            O => \N__31408\,
            I => \N__31404\
        );

    \I__6184\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31400\
        );

    \I__6183\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31397\
        );

    \I__6182\ : InMux
    port map (
            O => \N__31403\,
            I => \N__31394\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__31400\,
            I => \N__31389\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31389\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__31394\,
            I => \r_Clock_Count_0_adj_2454\
        );

    \I__6178\ : Odrv12
    port map (
            O => \N__31389\,
            I => \r_Clock_Count_0_adj_2454\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__31384\,
            I => \N__31380\
        );

    \I__6176\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31374\
        );

    \I__6175\ : InMux
    port map (
            O => \N__31380\,
            I => \N__31371\
        );

    \I__6174\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31368\
        );

    \I__6173\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31365\
        );

    \I__6172\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31362\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__31374\,
            I => \N__31356\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__31371\,
            I => \N__31356\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__31368\,
            I => \N__31353\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__31365\,
            I => \N__31350\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__31362\,
            I => \N__31347\
        );

    \I__6166\ : CascadeMux
    port map (
            O => \N__31361\,
            I => \N__31344\
        );

    \I__6165\ : Span4Mux_v
    port map (
            O => \N__31356\,
            I => \N__31338\
        );

    \I__6164\ : Span4Mux_v
    port map (
            O => \N__31353\,
            I => \N__31338\
        );

    \I__6163\ : Span4Mux_v
    port map (
            O => \N__31350\,
            I => \N__31333\
        );

    \I__6162\ : Span4Mux_v
    port map (
            O => \N__31347\,
            I => \N__31333\
        );

    \I__6161\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31330\
        );

    \I__6160\ : InMux
    port map (
            O => \N__31343\,
            I => \N__31327\
        );

    \I__6159\ : Sp12to4
    port map (
            O => \N__31338\,
            I => \N__31322\
        );

    \I__6158\ : Sp12to4
    port map (
            O => \N__31333\,
            I => \N__31322\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__31330\,
            I => \r_Bit_Index_1\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__31327\,
            I => \r_Bit_Index_1\
        );

    \I__6155\ : Odrv12
    port map (
            O => \N__31322\,
            I => \r_Bit_Index_1\
        );

    \I__6154\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31312\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__31312\,
            I => \N__31309\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__31309\,
            I => \N__31306\
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__31306\,
            I => n17398
        );

    \I__6150\ : CascadeMux
    port map (
            O => \N__31303\,
            I => \c0.n17918_cascade_\
        );

    \I__6149\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31297\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__31297\,
            I => \c0.n17343\
        );

    \I__6147\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31288\
        );

    \I__6146\ : InMux
    port map (
            O => \N__31293\,
            I => \N__31288\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31285\
        );

    \I__6144\ : Span4Mux_h
    port map (
            O => \N__31285\,
            I => \N__31281\
        );

    \I__6143\ : InMux
    port map (
            O => \N__31284\,
            I => \N__31278\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__31281\,
            I => \c0.n17769\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__31278\,
            I => \c0.n17769\
        );

    \I__6140\ : InMux
    port map (
            O => \N__31273\,
            I => \N__31270\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__31270\,
            I => \N__31267\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__31267\,
            I => \N__31264\
        );

    \I__6137\ : Odrv4
    port map (
            O => \N__31264\,
            I => \c0.n18\
        );

    \I__6136\ : InMux
    port map (
            O => \N__31261\,
            I => \N__31258\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__31258\,
            I => \N__31255\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__31255\,
            I => \N__31252\
        );

    \I__6133\ : Odrv4
    port map (
            O => \N__31252\,
            I => \c0.n17\
        );

    \I__6132\ : CascadeMux
    port map (
            O => \N__31249\,
            I => \N__31246\
        );

    \I__6131\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31243\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__31243\,
            I => \c0.n26_adj_2147\
        );

    \I__6129\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31237\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__31237\,
            I => \N__31234\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__31234\,
            I => \c0.n30_adj_2148\
        );

    \I__6126\ : CascadeMux
    port map (
            O => \N__31231\,
            I => \N__31225\
        );

    \I__6125\ : CascadeMux
    port map (
            O => \N__31230\,
            I => \N__31222\
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__31229\,
            I => \N__31218\
        );

    \I__6123\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31213\
        );

    \I__6122\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31209\
        );

    \I__6121\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31206\
        );

    \I__6120\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31203\
        );

    \I__6119\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31199\
        );

    \I__6118\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31194\
        );

    \I__6117\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31194\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__31213\,
            I => \N__31191\
        );

    \I__6115\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31188\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31181\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__31206\,
            I => \N__31181\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__31203\,
            I => \N__31181\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__31202\,
            I => \N__31178\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__31199\,
            I => \N__31175\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31172\
        );

    \I__6108\ : Span4Mux_v
    port map (
            O => \N__31191\,
            I => \N__31169\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__31188\,
            I => \N__31164\
        );

    \I__6106\ : Span4Mux_h
    port map (
            O => \N__31181\,
            I => \N__31164\
        );

    \I__6105\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31161\
        );

    \I__6104\ : Span4Mux_v
    port map (
            O => \N__31175\,
            I => \N__31158\
        );

    \I__6103\ : Span4Mux_h
    port map (
            O => \N__31172\,
            I => \N__31155\
        );

    \I__6102\ : Span4Mux_v
    port map (
            O => \N__31169\,
            I => \N__31150\
        );

    \I__6101\ : Span4Mux_h
    port map (
            O => \N__31164\,
            I => \N__31150\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__31161\,
            I => rx_data_5
        );

    \I__6099\ : Odrv4
    port map (
            O => \N__31158\,
            I => rx_data_5
        );

    \I__6098\ : Odrv4
    port map (
            O => \N__31155\,
            I => rx_data_5
        );

    \I__6097\ : Odrv4
    port map (
            O => \N__31150\,
            I => rx_data_5
        );

    \I__6096\ : InMux
    port map (
            O => \N__31141\,
            I => \N__31138\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__31138\,
            I => \N__31130\
        );

    \I__6094\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31127\
        );

    \I__6093\ : InMux
    port map (
            O => \N__31136\,
            I => \N__31124\
        );

    \I__6092\ : InMux
    port map (
            O => \N__31135\,
            I => \N__31121\
        );

    \I__6091\ : InMux
    port map (
            O => \N__31134\,
            I => \N__31116\
        );

    \I__6090\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31116\
        );

    \I__6089\ : Span4Mux_h
    port map (
            O => \N__31130\,
            I => \N__31104\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__31127\,
            I => \N__31095\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__31124\,
            I => \N__31095\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__31121\,
            I => \N__31095\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__31116\,
            I => \N__31095\
        );

    \I__6084\ : InMux
    port map (
            O => \N__31115\,
            I => \N__31092\
        );

    \I__6083\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31089\
        );

    \I__6082\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31086\
        );

    \I__6081\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31079\
        );

    \I__6080\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31079\
        );

    \I__6079\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31079\
        );

    \I__6078\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31072\
        );

    \I__6077\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31072\
        );

    \I__6076\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31072\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__31104\,
            I => \c0.n16882\
        );

    \I__6074\ : Odrv12
    port map (
            O => \N__31095\,
            I => \c0.n16882\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__31092\,
            I => \c0.n16882\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__31089\,
            I => \c0.n16882\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31086\,
            I => \c0.n16882\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__31079\,
            I => \c0.n16882\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__31072\,
            I => \c0.n16882\
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__31057\,
            I => \N__31054\
        );

    \I__6067\ : InMux
    port map (
            O => \N__31054\,
            I => \N__31050\
        );

    \I__6066\ : InMux
    port map (
            O => \N__31053\,
            I => \N__31047\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__31050\,
            I => \N__31044\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__31047\,
            I => \c0.data_in_frame_10_5\
        );

    \I__6063\ : Odrv4
    port map (
            O => \N__31044\,
            I => \c0.data_in_frame_10_5\
        );

    \I__6062\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31035\
        );

    \I__6061\ : InMux
    port map (
            O => \N__31038\,
            I => \N__31032\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__31035\,
            I => \N__31029\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__31032\,
            I => \N__31023\
        );

    \I__6058\ : Span4Mux_v
    port map (
            O => \N__31029\,
            I => \N__31018\
        );

    \I__6057\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31015\
        );

    \I__6056\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31010\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31026\,
            I => \N__31007\
        );

    \I__6054\ : Span4Mux_v
    port map (
            O => \N__31023\,
            I => \N__31004\
        );

    \I__6053\ : InMux
    port map (
            O => \N__31022\,
            I => \N__31001\
        );

    \I__6052\ : CascadeMux
    port map (
            O => \N__31021\,
            I => \N__30998\
        );

    \I__6051\ : Span4Mux_h
    port map (
            O => \N__31018\,
            I => \N__30989\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__31015\,
            I => \N__30989\
        );

    \I__6049\ : InMux
    port map (
            O => \N__31014\,
            I => \N__30986\
        );

    \I__6048\ : InMux
    port map (
            O => \N__31013\,
            I => \N__30983\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__31010\,
            I => \N__30974\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__31007\,
            I => \N__30974\
        );

    \I__6045\ : Sp12to4
    port map (
            O => \N__31004\,
            I => \N__30974\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__31001\,
            I => \N__30974\
        );

    \I__6043\ : InMux
    port map (
            O => \N__30998\,
            I => \N__30969\
        );

    \I__6042\ : InMux
    port map (
            O => \N__30997\,
            I => \N__30969\
        );

    \I__6041\ : InMux
    port map (
            O => \N__30996\,
            I => \N__30964\
        );

    \I__6040\ : InMux
    port map (
            O => \N__30995\,
            I => \N__30964\
        );

    \I__6039\ : InMux
    port map (
            O => \N__30994\,
            I => \N__30961\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__30989\,
            I => \N__30958\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__30986\,
            I => \r_SM_Main_1_adj_2444\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__30983\,
            I => \r_SM_Main_1_adj_2444\
        );

    \I__6035\ : Odrv12
    port map (
            O => \N__30974\,
            I => \r_SM_Main_1_adj_2444\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__30969\,
            I => \r_SM_Main_1_adj_2444\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__30964\,
            I => \r_SM_Main_1_adj_2444\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__30961\,
            I => \r_SM_Main_1_adj_2444\
        );

    \I__6031\ : Odrv4
    port map (
            O => \N__30958\,
            I => \r_SM_Main_1_adj_2444\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__30943\,
            I => \N__30940\
        );

    \I__6029\ : InMux
    port map (
            O => \N__30940\,
            I => \N__30937\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__30937\,
            I => \N__30934\
        );

    \I__6027\ : Span4Mux_h
    port map (
            O => \N__30934\,
            I => \N__30931\
        );

    \I__6026\ : Span4Mux_h
    port map (
            O => \N__30931\,
            I => \N__30928\
        );

    \I__6025\ : Odrv4
    port map (
            O => \N__30928\,
            I => \c0.tx2.n6480\
        );

    \I__6024\ : InMux
    port map (
            O => \N__30925\,
            I => \N__30922\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__30922\,
            I => \N__30919\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__30919\,
            I => \N__30916\
        );

    \I__6021\ : Span4Mux_h
    port map (
            O => \N__30916\,
            I => \N__30913\
        );

    \I__6020\ : Odrv4
    port map (
            O => \N__30913\,
            I => \c0.tx2.n1\
        );

    \I__6019\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30907\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__30907\,
            I => \N__30904\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__30904\,
            I => \c0.tx2.n10101\
        );

    \I__6016\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30898\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__30898\,
            I => \N__30894\
        );

    \I__6014\ : InMux
    port map (
            O => \N__30897\,
            I => \N__30891\
        );

    \I__6013\ : Span4Mux_h
    port map (
            O => \N__30894\,
            I => \N__30888\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__30891\,
            I => data_out_frame2_18_5
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__30888\,
            I => data_out_frame2_18_5
        );

    \I__6010\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30880\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__30880\,
            I => \N__30877\
        );

    \I__6008\ : Span4Mux_h
    port map (
            O => \N__30877\,
            I => \N__30871\
        );

    \I__6007\ : InMux
    port map (
            O => \N__30876\,
            I => \N__30868\
        );

    \I__6006\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30865\
        );

    \I__6005\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30861\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__30871\,
            I => \N__30854\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__30868\,
            I => \N__30854\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__30865\,
            I => \N__30854\
        );

    \I__6001\ : InMux
    port map (
            O => \N__30864\,
            I => \N__30849\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__30861\,
            I => \N__30845\
        );

    \I__5999\ : Span4Mux_h
    port map (
            O => \N__30854\,
            I => \N__30842\
        );

    \I__5998\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30837\
        );

    \I__5997\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30837\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__30849\,
            I => \N__30834\
        );

    \I__5995\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30831\
        );

    \I__5994\ : Span4Mux_v
    port map (
            O => \N__30845\,
            I => \N__30827\
        );

    \I__5993\ : Span4Mux_v
    port map (
            O => \N__30842\,
            I => \N__30824\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__30837\,
            I => \N__30821\
        );

    \I__5991\ : Span4Mux_h
    port map (
            O => \N__30834\,
            I => \N__30816\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__30831\,
            I => \N__30816\
        );

    \I__5989\ : InMux
    port map (
            O => \N__30830\,
            I => \N__30813\
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__30827\,
            I => \r_SM_Main_2_adj_2439\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__30824\,
            I => \r_SM_Main_2_adj_2439\
        );

    \I__5986\ : Odrv12
    port map (
            O => \N__30821\,
            I => \r_SM_Main_2_adj_2439\
        );

    \I__5985\ : Odrv4
    port map (
            O => \N__30816\,
            I => \r_SM_Main_2_adj_2439\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__30813\,
            I => \r_SM_Main_2_adj_2439\
        );

    \I__5983\ : InMux
    port map (
            O => \N__30802\,
            I => \N__30799\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__30799\,
            I => \N__30796\
        );

    \I__5981\ : Span4Mux_v
    port map (
            O => \N__30796\,
            I => \N__30793\
        );

    \I__5980\ : Span4Mux_h
    port map (
            O => \N__30793\,
            I => \N__30790\
        );

    \I__5979\ : Odrv4
    port map (
            O => \N__30790\,
            I => n13440
        );

    \I__5978\ : CascadeMux
    port map (
            O => \N__30787\,
            I => \N__30784\
        );

    \I__5977\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30781\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__30781\,
            I => \N__30776\
        );

    \I__5975\ : InMux
    port map (
            O => \N__30780\,
            I => \N__30771\
        );

    \I__5974\ : InMux
    port map (
            O => \N__30779\,
            I => \N__30771\
        );

    \I__5973\ : Span4Mux_v
    port map (
            O => \N__30776\,
            I => \N__30765\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__30771\,
            I => \N__30762\
        );

    \I__5971\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30756\
        );

    \I__5970\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30753\
        );

    \I__5969\ : CascadeMux
    port map (
            O => \N__30768\,
            I => \N__30750\
        );

    \I__5968\ : Span4Mux_h
    port map (
            O => \N__30765\,
            I => \N__30744\
        );

    \I__5967\ : Span4Mux_v
    port map (
            O => \N__30762\,
            I => \N__30744\
        );

    \I__5966\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30739\
        );

    \I__5965\ : InMux
    port map (
            O => \N__30760\,
            I => \N__30739\
        );

    \I__5964\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30736\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30730\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__30753\,
            I => \N__30730\
        );

    \I__5961\ : InMux
    port map (
            O => \N__30750\,
            I => \N__30727\
        );

    \I__5960\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30724\
        );

    \I__5959\ : Sp12to4
    port map (
            O => \N__30744\,
            I => \N__30721\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__30739\,
            I => \N__30716\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__30736\,
            I => \N__30716\
        );

    \I__5956\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30713\
        );

    \I__5955\ : Span4Mux_s2_h
    port map (
            O => \N__30730\,
            I => \N__30710\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__30727\,
            I => \r_SM_Main_1_adj_2440\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__30724\,
            I => \r_SM_Main_1_adj_2440\
        );

    \I__5952\ : Odrv12
    port map (
            O => \N__30721\,
            I => \r_SM_Main_1_adj_2440\
        );

    \I__5951\ : Odrv4
    port map (
            O => \N__30716\,
            I => \r_SM_Main_1_adj_2440\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__30713\,
            I => \r_SM_Main_1_adj_2440\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__30710\,
            I => \r_SM_Main_1_adj_2440\
        );

    \I__5948\ : InMux
    port map (
            O => \N__30697\,
            I => \N__30690\
        );

    \I__5947\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30687\
        );

    \I__5946\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30684\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__30694\,
            I => \N__30680\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__30693\,
            I => \N__30676\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30669\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__30687\,
            I => \N__30669\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__30684\,
            I => \N__30669\
        );

    \I__5940\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30666\
        );

    \I__5939\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30662\
        );

    \I__5938\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30659\
        );

    \I__5937\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30656\
        );

    \I__5936\ : Span4Mux_v
    port map (
            O => \N__30669\,
            I => \N__30653\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__30666\,
            I => \N__30650\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__30665\,
            I => \N__30646\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__30662\,
            I => \N__30639\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__30659\,
            I => \N__30639\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__30656\,
            I => \N__30639\
        );

    \I__5930\ : Span4Mux_h
    port map (
            O => \N__30653\,
            I => \N__30636\
        );

    \I__5929\ : Span4Mux_v
    port map (
            O => \N__30650\,
            I => \N__30633\
        );

    \I__5928\ : InMux
    port map (
            O => \N__30649\,
            I => \N__30628\
        );

    \I__5927\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30628\
        );

    \I__5926\ : Odrv12
    port map (
            O => \N__30639\,
            I => rx_data_1
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__30636\,
            I => rx_data_1
        );

    \I__5924\ : Odrv4
    port map (
            O => \N__30633\,
            I => rx_data_1
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__30628\,
            I => rx_data_1
        );

    \I__5922\ : InMux
    port map (
            O => \N__30619\,
            I => \N__30615\
        );

    \I__5921\ : InMux
    port map (
            O => \N__30618\,
            I => \N__30612\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__30615\,
            I => \N__30609\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__30612\,
            I => \c0.data_in_frame_2_1\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__30609\,
            I => \c0.data_in_frame_2_1\
        );

    \I__5917\ : InMux
    port map (
            O => \N__30604\,
            I => \N__30598\
        );

    \I__5916\ : InMux
    port map (
            O => \N__30603\,
            I => \N__30598\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__30598\,
            I => \N__30594\
        );

    \I__5914\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30591\
        );

    \I__5913\ : Sp12to4
    port map (
            O => \N__30594\,
            I => \N__30588\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__30591\,
            I => \c0.tx2.tx2_active\
        );

    \I__5911\ : Odrv12
    port map (
            O => \N__30588\,
            I => \c0.tx2.tx2_active\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__30583\,
            I => \c0.n17334_cascade_\
        );

    \I__5909\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30576\
        );

    \I__5908\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30572\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__30576\,
            I => \N__30569\
        );

    \I__5906\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30566\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__30572\,
            I => \N__30563\
        );

    \I__5904\ : Odrv12
    port map (
            O => \N__30569\,
            I => \c0.n2334\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__30566\,
            I => \c0.n2334\
        );

    \I__5902\ : Odrv4
    port map (
            O => \N__30563\,
            I => \c0.n2334\
        );

    \I__5901\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30552\
        );

    \I__5900\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30549\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__30552\,
            I => \N__30546\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__30549\,
            I => \N__30543\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__30546\,
            I => \c0.n2351\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__30543\,
            I => \c0.n2351\
        );

    \I__5895\ : InMux
    port map (
            O => \N__30538\,
            I => \N__30535\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__30535\,
            I => \c0.n18_adj_2343\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__30532\,
            I => \N__30528\
        );

    \I__5892\ : CascadeMux
    port map (
            O => \N__30531\,
            I => \N__30525\
        );

    \I__5891\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30519\
        );

    \I__5890\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30516\
        );

    \I__5889\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30513\
        );

    \I__5888\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30509\
        );

    \I__5887\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30506\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30500\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30500\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__30513\,
            I => \N__30497\
        );

    \I__5883\ : InMux
    port map (
            O => \N__30512\,
            I => \N__30494\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__30509\,
            I => \N__30489\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__30506\,
            I => \N__30489\
        );

    \I__5880\ : InMux
    port map (
            O => \N__30505\,
            I => \N__30484\
        );

    \I__5879\ : Span4Mux_v
    port map (
            O => \N__30500\,
            I => \N__30479\
        );

    \I__5878\ : Span4Mux_h
    port map (
            O => \N__30497\,
            I => \N__30479\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__30494\,
            I => \N__30476\
        );

    \I__5876\ : Span4Mux_v
    port map (
            O => \N__30489\,
            I => \N__30473\
        );

    \I__5875\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30470\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__30487\,
            I => \N__30467\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__30484\,
            I => \N__30464\
        );

    \I__5872\ : Span4Mux_h
    port map (
            O => \N__30479\,
            I => \N__30461\
        );

    \I__5871\ : Span4Mux_v
    port map (
            O => \N__30476\,
            I => \N__30454\
        );

    \I__5870\ : Span4Mux_s3_h
    port map (
            O => \N__30473\,
            I => \N__30454\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__30470\,
            I => \N__30454\
        );

    \I__5868\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30451\
        );

    \I__5867\ : Odrv12
    port map (
            O => \N__30464\,
            I => rx_data_3
        );

    \I__5866\ : Odrv4
    port map (
            O => \N__30461\,
            I => rx_data_3
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__30454\,
            I => rx_data_3
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__30451\,
            I => rx_data_3
        );

    \I__5863\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30438\
        );

    \I__5862\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30431\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30428\
        );

    \I__5860\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30423\
        );

    \I__5859\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30423\
        );

    \I__5858\ : InMux
    port map (
            O => \N__30435\,
            I => \N__30418\
        );

    \I__5857\ : InMux
    port map (
            O => \N__30434\,
            I => \N__30415\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__30431\,
            I => \N__30412\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__30428\,
            I => \N__30407\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__30423\,
            I => \N__30407\
        );

    \I__5853\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30402\
        );

    \I__5852\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30402\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30397\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__30415\,
            I => \N__30397\
        );

    \I__5849\ : Span4Mux_v
    port map (
            O => \N__30412\,
            I => \N__30390\
        );

    \I__5848\ : Span4Mux_h
    port map (
            O => \N__30407\,
            I => \N__30390\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30390\
        );

    \I__5846\ : Span12Mux_s11_v
    port map (
            O => \N__30397\,
            I => \N__30387\
        );

    \I__5845\ : Span4Mux_v
    port map (
            O => \N__30390\,
            I => \N__30384\
        );

    \I__5844\ : Odrv12
    port map (
            O => \N__30387\,
            I => n16897
        );

    \I__5843\ : Odrv4
    port map (
            O => \N__30384\,
            I => n16897
        );

    \I__5842\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30372\
        );

    \I__5841\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30372\
        );

    \I__5840\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30368\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__30372\,
            I => \N__30365\
        );

    \I__5838\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30362\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__30368\,
            I => \N__30359\
        );

    \I__5836\ : Span4Mux_h
    port map (
            O => \N__30365\,
            I => \N__30356\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__30362\,
            I => data_in_frame_0_3
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__30359\,
            I => data_in_frame_0_3
        );

    \I__5833\ : Odrv4
    port map (
            O => \N__30356\,
            I => data_in_frame_0_3
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__30349\,
            I => \c0.n17337_cascade_\
        );

    \I__5831\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30343\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__30343\,
            I => \N__30340\
        );

    \I__5829\ : Span4Mux_v
    port map (
            O => \N__30340\,
            I => \N__30336\
        );

    \I__5828\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30331\
        );

    \I__5827\ : Span4Mux_h
    port map (
            O => \N__30336\,
            I => \N__30328\
        );

    \I__5826\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30323\
        );

    \I__5825\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30323\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__30331\,
            I => data_in_frame_0_4
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__30328\,
            I => data_in_frame_0_4
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__30323\,
            I => data_in_frame_0_4
        );

    \I__5821\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30312\
        );

    \I__5820\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30309\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__30312\,
            I => \N__30306\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__30309\,
            I => \N__30301\
        );

    \I__5817\ : Span4Mux_h
    port map (
            O => \N__30306\,
            I => \N__30296\
        );

    \I__5816\ : InMux
    port map (
            O => \N__30305\,
            I => \N__30291\
        );

    \I__5815\ : InMux
    port map (
            O => \N__30304\,
            I => \N__30291\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__30301\,
            I => \N__30288\
        );

    \I__5813\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30285\
        );

    \I__5812\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30282\
        );

    \I__5811\ : Odrv4
    port map (
            O => \N__30296\,
            I => data_in_frame_0_5
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__30291\,
            I => data_in_frame_0_5
        );

    \I__5809\ : Odrv4
    port map (
            O => \N__30288\,
            I => data_in_frame_0_5
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__30285\,
            I => data_in_frame_0_5
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__30282\,
            I => data_in_frame_0_5
        );

    \I__5806\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30268\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__30268\,
            I => \N__30264\
        );

    \I__5804\ : InMux
    port map (
            O => \N__30267\,
            I => \N__30261\
        );

    \I__5803\ : Span4Mux_v
    port map (
            O => \N__30264\,
            I => \N__30258\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__30261\,
            I => \N__30255\
        );

    \I__5801\ : Span4Mux_h
    port map (
            O => \N__30258\,
            I => \N__30252\
        );

    \I__5800\ : Span4Mux_v
    port map (
            O => \N__30255\,
            I => \N__30249\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__30252\,
            I => \c0.n2338\
        );

    \I__5798\ : Odrv4
    port map (
            O => \N__30249\,
            I => \c0.n2338\
        );

    \I__5797\ : InMux
    port map (
            O => \N__30244\,
            I => \N__30241\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__30241\,
            I => \N__30238\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__30238\,
            I => \N__30234\
        );

    \I__5794\ : InMux
    port map (
            O => \N__30237\,
            I => \N__30231\
        );

    \I__5793\ : Span4Mux_h
    port map (
            O => \N__30234\,
            I => \N__30228\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__30231\,
            I => \c0.data_in_frame_2_6\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__30228\,
            I => \c0.data_in_frame_2_6\
        );

    \I__5790\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30220\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__30220\,
            I => \N__30216\
        );

    \I__5788\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30213\
        );

    \I__5787\ : Span4Mux_h
    port map (
            O => \N__30216\,
            I => \N__30210\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__30213\,
            I => \N__30207\
        );

    \I__5785\ : Span4Mux_h
    port map (
            O => \N__30210\,
            I => \N__30204\
        );

    \I__5784\ : Odrv4
    port map (
            O => \N__30207\,
            I => \c0.data_in_frame_2_0\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__30204\,
            I => \c0.data_in_frame_2_0\
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__30199\,
            I => \c0.n2338_cascade_\
        );

    \I__5781\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__30193\,
            I => \N__30188\
        );

    \I__5779\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30185\
        );

    \I__5778\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30182\
        );

    \I__5777\ : Span4Mux_v
    port map (
            O => \N__30188\,
            I => \N__30177\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__30185\,
            I => \N__30177\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__30182\,
            I => \c0.n2352\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__30177\,
            I => \c0.n2352\
        );

    \I__5773\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30169\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__30169\,
            I => \N__30166\
        );

    \I__5771\ : Span4Mux_h
    port map (
            O => \N__30166\,
            I => \N__30163\
        );

    \I__5770\ : Odrv4
    port map (
            O => \N__30163\,
            I => \c0.n26_adj_2344\
        );

    \I__5769\ : CascadeMux
    port map (
            O => \N__30160\,
            I => \c0.n17_adj_2346_cascade_\
        );

    \I__5768\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__30154\,
            I => \c0.n30_adj_2345\
        );

    \I__5766\ : CascadeMux
    port map (
            O => \N__30151\,
            I => \n31_cascade_\
        );

    \I__5765\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30145\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__30145\,
            I => \N__30142\
        );

    \I__5763\ : Odrv4
    port map (
            O => \N__30142\,
            I => \c0.n5_adj_2322\
        );

    \I__5762\ : CascadeMux
    port map (
            O => \N__30139\,
            I => \c0.n5_cascade_\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__30136\,
            I => \c0.n17328_cascade_\
        );

    \I__5760\ : InMux
    port map (
            O => \N__30133\,
            I => \N__30130\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__30130\,
            I => \N__30126\
        );

    \I__5758\ : InMux
    port map (
            O => \N__30129\,
            I => \N__30123\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__30126\,
            I => \N__30118\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__30123\,
            I => \N__30118\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__30118\,
            I => \N__30114\
        );

    \I__5754\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30111\
        );

    \I__5753\ : Span4Mux_h
    port map (
            O => \N__30114\,
            I => \N__30104\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__30111\,
            I => \N__30104\
        );

    \I__5751\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30101\
        );

    \I__5750\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30098\
        );

    \I__5749\ : Span4Mux_v
    port map (
            O => \N__30104\,
            I => \N__30095\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__30101\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__30098\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5746\ : Odrv4
    port map (
            O => \N__30095\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5745\ : CascadeMux
    port map (
            O => \N__30088\,
            I => \N__30085\
        );

    \I__5744\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30081\
        );

    \I__5743\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30078\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__30081\,
            I => \N__30073\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__30078\,
            I => \N__30073\
        );

    \I__5740\ : Span4Mux_h
    port map (
            O => \N__30073\,
            I => \N__30070\
        );

    \I__5739\ : Span4Mux_h
    port map (
            O => \N__30070\,
            I => \N__30067\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__30067\,
            I => \c0.n16905\
        );

    \I__5737\ : CascadeMux
    port map (
            O => \N__30064\,
            I => \N__30061\
        );

    \I__5736\ : InMux
    port map (
            O => \N__30061\,
            I => \N__30058\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__30058\,
            I => \N__30052\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30049\
        );

    \I__5733\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30044\
        );

    \I__5732\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30044\
        );

    \I__5731\ : Span4Mux_v
    port map (
            O => \N__30052\,
            I => \N__30041\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__30049\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__30044\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__5728\ : Odrv4
    port map (
            O => \N__30041\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__5727\ : SRMux
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__30031\,
            I => \c0.n16345\
        );

    \I__5725\ : InMux
    port map (
            O => \N__30028\,
            I => \N__30022\
        );

    \I__5724\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30019\
        );

    \I__5723\ : InMux
    port map (
            O => \N__30026\,
            I => \N__30015\
        );

    \I__5722\ : InMux
    port map (
            O => \N__30025\,
            I => \N__30012\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__30022\,
            I => \N__30009\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__30019\,
            I => \N__30006\
        );

    \I__5719\ : InMux
    port map (
            O => \N__30018\,
            I => \N__30003\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__30015\,
            I => \N__30000\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__30012\,
            I => \N__29995\
        );

    \I__5716\ : Span4Mux_h
    port map (
            O => \N__30009\,
            I => \N__29995\
        );

    \I__5715\ : Span4Mux_v
    port map (
            O => \N__30006\,
            I => \N__29992\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__30003\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__5713\ : Odrv12
    port map (
            O => \N__30000\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__5712\ : Odrv4
    port map (
            O => \N__29995\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__29992\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__5710\ : CascadeMux
    port map (
            O => \N__29983\,
            I => \N__29978\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__29982\,
            I => \N__29975\
        );

    \I__5708\ : CascadeMux
    port map (
            O => \N__29981\,
            I => \N__29969\
        );

    \I__5707\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29955\
        );

    \I__5706\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29955\
        );

    \I__5705\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29955\
        );

    \I__5704\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29955\
        );

    \I__5703\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29955\
        );

    \I__5702\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29949\
        );

    \I__5701\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29949\
        );

    \I__5700\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29946\
        );

    \I__5699\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29942\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__29955\,
            I => \N__29938\
        );

    \I__5697\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29935\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__29949\,
            I => \N__29930\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__29946\,
            I => \N__29930\
        );

    \I__5694\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29927\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__29942\,
            I => \N__29924\
        );

    \I__5692\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29921\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__29938\,
            I => \N__29912\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__29935\,
            I => \N__29912\
        );

    \I__5689\ : Span4Mux_v
    port map (
            O => \N__29930\,
            I => \N__29907\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__29927\,
            I => \N__29907\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__29924\,
            I => \N__29904\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__29921\,
            I => \N__29901\
        );

    \I__5685\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29898\
        );

    \I__5684\ : InMux
    port map (
            O => \N__29919\,
            I => \N__29895\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__29918\,
            I => \N__29890\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__29917\,
            I => \N__29886\
        );

    \I__5681\ : Span4Mux_h
    port map (
            O => \N__29912\,
            I => \N__29881\
        );

    \I__5680\ : Span4Mux_v
    port map (
            O => \N__29907\,
            I => \N__29878\
        );

    \I__5679\ : Span4Mux_v
    port map (
            O => \N__29904\,
            I => \N__29873\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__29901\,
            I => \N__29873\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__29898\,
            I => \N__29868\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__29895\,
            I => \N__29868\
        );

    \I__5675\ : InMux
    port map (
            O => \N__29894\,
            I => \N__29865\
        );

    \I__5674\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29862\
        );

    \I__5673\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29851\
        );

    \I__5672\ : InMux
    port map (
            O => \N__29889\,
            I => \N__29851\
        );

    \I__5671\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29851\
        );

    \I__5670\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29851\
        );

    \I__5669\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29851\
        );

    \I__5668\ : Odrv4
    port map (
            O => \N__29881\,
            I => \c0.n4\
        );

    \I__5667\ : Odrv4
    port map (
            O => \N__29878\,
            I => \c0.n4\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__29873\,
            I => \c0.n4\
        );

    \I__5665\ : Odrv12
    port map (
            O => \N__29868\,
            I => \c0.n4\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__29865\,
            I => \c0.n4\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__29862\,
            I => \c0.n4\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__29851\,
            I => \c0.n4\
        );

    \I__5661\ : SRMux
    port map (
            O => \N__29836\,
            I => \N__29833\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__29833\,
            I => \N__29830\
        );

    \I__5659\ : Span4Mux_h
    port map (
            O => \N__29830\,
            I => \N__29827\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__29827\,
            I => \c0.n16339\
        );

    \I__5657\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29820\
        );

    \I__5656\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29817\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29813\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__29817\,
            I => \N__29810\
        );

    \I__5653\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29806\
        );

    \I__5652\ : Span4Mux_v
    port map (
            O => \N__29813\,
            I => \N__29803\
        );

    \I__5651\ : Span4Mux_v
    port map (
            O => \N__29810\,
            I => \N__29800\
        );

    \I__5650\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29797\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__29806\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__29803\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__29800\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__29797\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__29788\,
            I => \N__29785\
        );

    \I__5644\ : InMux
    port map (
            O => \N__29785\,
            I => \N__29782\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__29782\,
            I => \N__29779\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__29779\,
            I => \c0.n16871\
        );

    \I__5641\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29772\
        );

    \I__5640\ : InMux
    port map (
            O => \N__29775\,
            I => \N__29769\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__29772\,
            I => \N__29766\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__29769\,
            I => \N__29763\
        );

    \I__5637\ : Span12Mux_v
    port map (
            O => \N__29766\,
            I => \N__29760\
        );

    \I__5636\ : Span4Mux_h
    port map (
            O => \N__29763\,
            I => \N__29757\
        );

    \I__5635\ : Odrv12
    port map (
            O => \N__29760\,
            I => \c0.n16772\
        );

    \I__5634\ : Odrv4
    port map (
            O => \N__29757\,
            I => \c0.n16772\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__29752\,
            I => \c0.n17349_cascade_\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__29749\,
            I => \N__29746\
        );

    \I__5631\ : InMux
    port map (
            O => \N__29746\,
            I => \N__29736\
        );

    \I__5630\ : InMux
    port map (
            O => \N__29745\,
            I => \N__29736\
        );

    \I__5629\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29736\
        );

    \I__5628\ : InMux
    port map (
            O => \N__29743\,
            I => \N__29729\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__29736\,
            I => \N__29723\
        );

    \I__5626\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29716\
        );

    \I__5625\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29716\
        );

    \I__5624\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29716\
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__29732\,
            I => \N__29713\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__29729\,
            I => \N__29702\
        );

    \I__5621\ : InMux
    port map (
            O => \N__29728\,
            I => \N__29695\
        );

    \I__5620\ : InMux
    port map (
            O => \N__29727\,
            I => \N__29695\
        );

    \I__5619\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29695\
        );

    \I__5618\ : Span4Mux_h
    port map (
            O => \N__29723\,
            I => \N__29690\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__29716\,
            I => \N__29690\
        );

    \I__5616\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29685\
        );

    \I__5615\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29685\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__29711\,
            I => \N__29681\
        );

    \I__5613\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29672\
        );

    \I__5612\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29672\
        );

    \I__5611\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29672\
        );

    \I__5610\ : CascadeMux
    port map (
            O => \N__29707\,
            I => \N__29669\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__29706\,
            I => \N__29666\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__29705\,
            I => \N__29662\
        );

    \I__5607\ : Span4Mux_h
    port map (
            O => \N__29702\,
            I => \N__29653\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__29695\,
            I => \N__29650\
        );

    \I__5605\ : Span4Mux_v
    port map (
            O => \N__29690\,
            I => \N__29645\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__29685\,
            I => \N__29642\
        );

    \I__5603\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29633\
        );

    \I__5602\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29633\
        );

    \I__5601\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29633\
        );

    \I__5600\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29633\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__29672\,
            I => \N__29630\
        );

    \I__5598\ : InMux
    port map (
            O => \N__29669\,
            I => \N__29619\
        );

    \I__5597\ : InMux
    port map (
            O => \N__29666\,
            I => \N__29619\
        );

    \I__5596\ : InMux
    port map (
            O => \N__29665\,
            I => \N__29619\
        );

    \I__5595\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29619\
        );

    \I__5594\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29619\
        );

    \I__5593\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29608\
        );

    \I__5592\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29608\
        );

    \I__5591\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29608\
        );

    \I__5590\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29608\
        );

    \I__5589\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29608\
        );

    \I__5588\ : Span4Mux_h
    port map (
            O => \N__29653\,
            I => \N__29603\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__29650\,
            I => \N__29603\
        );

    \I__5586\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29598\
        );

    \I__5585\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29598\
        );

    \I__5584\ : Odrv4
    port map (
            O => \N__29645\,
            I => \c0.n1439\
        );

    \I__5583\ : Odrv12
    port map (
            O => \N__29642\,
            I => \c0.n1439\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__29633\,
            I => \c0.n1439\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__29630\,
            I => \c0.n1439\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__29619\,
            I => \c0.n1439\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__29608\,
            I => \c0.n1439\
        );

    \I__5578\ : Odrv4
    port map (
            O => \N__29603\,
            I => \c0.n1439\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__29598\,
            I => \c0.n1439\
        );

    \I__5576\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29578\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__29578\,
            I => \N__29575\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__29575\,
            I => \N__29571\
        );

    \I__5573\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29568\
        );

    \I__5572\ : Span4Mux_h
    port map (
            O => \N__29571\,
            I => \N__29565\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__29568\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_0\
        );

    \I__5570\ : Odrv4
    port map (
            O => \N__29565\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_0\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__29560\,
            I => \c0.n17590_cascade_\
        );

    \I__5568\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29554\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__29554\,
            I => n18026
        );

    \I__5566\ : SRMux
    port map (
            O => \N__29551\,
            I => \N__29548\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__29548\,
            I => \N__29545\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__29545\,
            I => \N__29542\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__29542\,
            I => \N__29539\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__29539\,
            I => \c0.n16347\
        );

    \I__5561\ : CascadeMux
    port map (
            O => \N__29536\,
            I => \N__29533\
        );

    \I__5560\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29529\
        );

    \I__5559\ : InMux
    port map (
            O => \N__29532\,
            I => \N__29526\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__29529\,
            I => \N__29523\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29520\
        );

    \I__5556\ : Span4Mux_h
    port map (
            O => \N__29523\,
            I => \N__29517\
        );

    \I__5555\ : Span4Mux_h
    port map (
            O => \N__29520\,
            I => \N__29514\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__29517\,
            I => \c0.n16761\
        );

    \I__5553\ : Odrv4
    port map (
            O => \N__29514\,
            I => \c0.n16761\
        );

    \I__5552\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29506\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29500\
        );

    \I__5550\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29493\
        );

    \I__5549\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29493\
        );

    \I__5548\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29493\
        );

    \I__5547\ : Span4Mux_h
    port map (
            O => \N__29500\,
            I => \N__29490\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__29493\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__29490\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__5544\ : SRMux
    port map (
            O => \N__29485\,
            I => \N__29482\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__29482\,
            I => \N__29479\
        );

    \I__5542\ : Odrv4
    port map (
            O => \N__29479\,
            I => \c0.n16353\
        );

    \I__5541\ : CascadeMux
    port map (
            O => \N__29476\,
            I => \N__29469\
        );

    \I__5540\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29466\
        );

    \I__5539\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29463\
        );

    \I__5538\ : InMux
    port map (
            O => \N__29473\,
            I => \N__29460\
        );

    \I__5537\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29455\
        );

    \I__5536\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29455\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__29466\,
            I => \N__29452\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__29463\,
            I => \N__29449\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__29460\,
            I => \N__29444\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__29455\,
            I => \N__29444\
        );

    \I__5531\ : Span4Mux_h
    port map (
            O => \N__29452\,
            I => \N__29439\
        );

    \I__5530\ : Span4Mux_h
    port map (
            O => \N__29449\,
            I => \N__29439\
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__29444\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__29439\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__5527\ : SRMux
    port map (
            O => \N__29434\,
            I => \N__29431\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__29431\,
            I => \c0.n16361\
        );

    \I__5525\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29422\
        );

    \I__5524\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29422\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__29422\,
            I => \r_Tx_Data_0\
        );

    \I__5522\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29416\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__29416\,
            I => \N__29413\
        );

    \I__5520\ : Span4Mux_h
    port map (
            O => \N__29413\,
            I => \N__29410\
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__29410\,
            I => n17394
        );

    \I__5518\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29404\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__29404\,
            I => \N__29401\
        );

    \I__5516\ : Odrv4
    port map (
            O => \N__29401\,
            I => \c0.n8_adj_2160\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__29398\,
            I => \c0.n15_cascade_\
        );

    \I__5514\ : CascadeMux
    port map (
            O => \N__29395\,
            I => \c0.n12_adj_2150_cascade_\
        );

    \I__5513\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29388\
        );

    \I__5512\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29385\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__29388\,
            I => \r_Tx_Data_2\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__29385\,
            I => \r_Tx_Data_2\
        );

    \I__5509\ : CascadeMux
    port map (
            O => \N__29380\,
            I => \N__29377\
        );

    \I__5508\ : InMux
    port map (
            O => \N__29377\,
            I => \N__29374\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__29374\,
            I => n10_adj_2426
        );

    \I__5506\ : CascadeMux
    port map (
            O => \N__29371\,
            I => \n10_adj_2407_cascade_\
        );

    \I__5505\ : InMux
    port map (
            O => \N__29368\,
            I => \N__29365\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__29365\,
            I => \N__29362\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__29362\,
            I => \N__29358\
        );

    \I__5502\ : InMux
    port map (
            O => \N__29361\,
            I => \N__29355\
        );

    \I__5501\ : Span4Mux_h
    port map (
            O => \N__29358\,
            I => \N__29352\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__29355\,
            I => \r_Tx_Data_4\
        );

    \I__5499\ : Odrv4
    port map (
            O => \N__29352\,
            I => \r_Tx_Data_4\
        );

    \I__5498\ : CascadeMux
    port map (
            O => \N__29347\,
            I => \c0.tx2.o_Tx_Serial_N_2064_cascade_\
        );

    \I__5497\ : CascadeMux
    port map (
            O => \N__29344\,
            I => \N__29337\
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__29343\,
            I => \N__29334\
        );

    \I__5495\ : InMux
    port map (
            O => \N__29342\,
            I => \N__29331\
        );

    \I__5494\ : InMux
    port map (
            O => \N__29341\,
            I => \N__29328\
        );

    \I__5493\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29322\
        );

    \I__5492\ : InMux
    port map (
            O => \N__29337\,
            I => \N__29315\
        );

    \I__5491\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29315\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__29331\,
            I => \N__29310\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__29328\,
            I => \N__29310\
        );

    \I__5488\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29307\
        );

    \I__5487\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29302\
        );

    \I__5486\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29302\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__29322\,
            I => \N__29299\
        );

    \I__5484\ : InMux
    port map (
            O => \N__29321\,
            I => \N__29296\
        );

    \I__5483\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29293\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__29315\,
            I => \N__29288\
        );

    \I__5481\ : Span4Mux_h
    port map (
            O => \N__29310\,
            I => \N__29288\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__29307\,
            I => \r_SM_Main_0_adj_2445\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__29302\,
            I => \r_SM_Main_0_adj_2445\
        );

    \I__5478\ : Odrv12
    port map (
            O => \N__29299\,
            I => \r_SM_Main_0_adj_2445\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__29296\,
            I => \r_SM_Main_0_adj_2445\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__29293\,
            I => \r_SM_Main_0_adj_2445\
        );

    \I__5475\ : Odrv4
    port map (
            O => \N__29288\,
            I => \r_SM_Main_0_adj_2445\
        );

    \I__5474\ : InMux
    port map (
            O => \N__29275\,
            I => \N__29272\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__29272\,
            I => \N__29269\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__29269\,
            I => n3
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__29266\,
            I => \N__29263\
        );

    \I__5470\ : InMux
    port map (
            O => \N__29263\,
            I => \N__29260\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__29260\,
            I => n5029
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__29257\,
            I => \N__29252\
        );

    \I__5467\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29249\
        );

    \I__5466\ : InMux
    port map (
            O => \N__29255\,
            I => \N__29244\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29244\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__29249\,
            I => \r_Bit_Index_2_adj_2455\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__29244\,
            I => \r_Bit_Index_2_adj_2455\
        );

    \I__5462\ : CascadeMux
    port map (
            O => \N__29239\,
            I => \N__29236\
        );

    \I__5461\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29233\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29229\
        );

    \I__5459\ : InMux
    port map (
            O => \N__29232\,
            I => \N__29226\
        );

    \I__5458\ : Odrv12
    port map (
            O => \N__29229\,
            I => \c0.tx2.n13281\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__29226\,
            I => \c0.tx2.n13281\
        );

    \I__5456\ : CascadeMux
    port map (
            O => \N__29221\,
            I => \c0.n2_adj_2266_cascade_\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__29218\,
            I => \c0.n18098_cascade_\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__29215\,
            I => \c0.n10_adj_2139_cascade_\
        );

    \I__5453\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29209\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__29209\,
            I => \N__29206\
        );

    \I__5451\ : Span4Mux_h
    port map (
            O => \N__29206\,
            I => \N__29203\
        );

    \I__5450\ : IoSpan4Mux
    port map (
            O => \N__29203\,
            I => \N__29200\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__29200\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__5448\ : CascadeMux
    port map (
            O => \N__29197\,
            I => \c0.tx2.n18113_cascade_\
        );

    \I__5447\ : InMux
    port map (
            O => \N__29194\,
            I => \N__29188\
        );

    \I__5446\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29188\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__29188\,
            I => n10398
        );

    \I__5444\ : InMux
    port map (
            O => \N__29185\,
            I => \N__29177\
        );

    \I__5443\ : InMux
    port map (
            O => \N__29184\,
            I => \N__29177\
        );

    \I__5442\ : InMux
    port map (
            O => \N__29183\,
            I => \N__29172\
        );

    \I__5441\ : InMux
    port map (
            O => \N__29182\,
            I => \N__29172\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29169\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__29172\,
            I => \N__29166\
        );

    \I__5438\ : Span12Mux_h
    port map (
            O => \N__29169\,
            I => \N__29163\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__29166\,
            I => \N__29160\
        );

    \I__5436\ : Odrv12
    port map (
            O => \N__29163\,
            I => n17194
        );

    \I__5435\ : Odrv4
    port map (
            O => \N__29160\,
            I => n17194
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__29155\,
            I => \n10398_cascade_\
        );

    \I__5433\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29149\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__29149\,
            I => \c0.tx2.n17906\
        );

    \I__5431\ : InMux
    port map (
            O => \N__29146\,
            I => \N__29143\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__29143\,
            I => \N__29140\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__29140\,
            I => \c0.tx2.n18116\
        );

    \I__5428\ : InMux
    port map (
            O => \N__29137\,
            I => \N__29134\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__29134\,
            I => \N__29129\
        );

    \I__5426\ : InMux
    port map (
            O => \N__29133\,
            I => \N__29126\
        );

    \I__5425\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29123\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__29129\,
            I => \N__29116\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__29126\,
            I => \N__29116\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__29123\,
            I => \N__29116\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__29116\,
            I => \N__29111\
        );

    \I__5420\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29106\
        );

    \I__5419\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29106\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__29111\,
            I => \c0.data_in_frame_1_1\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__29106\,
            I => \c0.data_in_frame_1_1\
        );

    \I__5416\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29098\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29095\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__29095\,
            I => \N__29092\
        );

    \I__5413\ : Odrv4
    port map (
            O => \N__29092\,
            I => \c0.n17014\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__29089\,
            I => \c0.n23_adj_2156_cascade_\
        );

    \I__5411\ : InMux
    port map (
            O => \N__29086\,
            I => \N__29082\
        );

    \I__5410\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29079\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__29082\,
            I => \N__29076\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__29079\,
            I => \N__29073\
        );

    \I__5407\ : Span4Mux_h
    port map (
            O => \N__29076\,
            I => \N__29070\
        );

    \I__5406\ : Span4Mux_h
    port map (
            O => \N__29073\,
            I => \N__29067\
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__29070\,
            I => \c0.n17001\
        );

    \I__5404\ : Odrv4
    port map (
            O => \N__29067\,
            I => \c0.n17001\
        );

    \I__5403\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29059\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__29059\,
            I => \c0.n28_adj_2183\
        );

    \I__5401\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29052\
        );

    \I__5400\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29046\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__29052\,
            I => \N__29042\
        );

    \I__5398\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29037\
        );

    \I__5397\ : InMux
    port map (
            O => \N__29050\,
            I => \N__29037\
        );

    \I__5396\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29033\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__29046\,
            I => \N__29030\
        );

    \I__5394\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29027\
        );

    \I__5393\ : Span4Mux_h
    port map (
            O => \N__29042\,
            I => \N__29022\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__29037\,
            I => \N__29022\
        );

    \I__5391\ : InMux
    port map (
            O => \N__29036\,
            I => \N__29019\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__29033\,
            I => \N__29014\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__29030\,
            I => \N__29014\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__29027\,
            I => data_in_frame_0_6
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__29022\,
            I => data_in_frame_0_6
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__29019\,
            I => data_in_frame_0_6
        );

    \I__5385\ : Odrv4
    port map (
            O => \N__29014\,
            I => data_in_frame_0_6
        );

    \I__5384\ : InMux
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__28999\,
            I => \c0.n2340\
        );

    \I__5381\ : CascadeMux
    port map (
            O => \N__28996\,
            I => \N__28993\
        );

    \I__5380\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28989\
        );

    \I__5379\ : InMux
    port map (
            O => \N__28992\,
            I => \N__28986\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__28989\,
            I => \N__28983\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__28986\,
            I => \c0.data_in_frame_9_0\
        );

    \I__5376\ : Odrv12
    port map (
            O => \N__28983\,
            I => \c0.data_in_frame_9_0\
        );

    \I__5375\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28974\
        );

    \I__5374\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28971\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__28974\,
            I => \N__28968\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__28971\,
            I => \N__28965\
        );

    \I__5371\ : Odrv12
    port map (
            O => \N__28968\,
            I => \c0.n17004\
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__28965\,
            I => \c0.n17004\
        );

    \I__5369\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28957\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__28957\,
            I => \c0.n19\
        );

    \I__5367\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28950\
        );

    \I__5366\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28947\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__28950\,
            I => \N__28944\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__28947\,
            I => data_in_frame_7_3
        );

    \I__5363\ : Odrv12
    port map (
            O => \N__28944\,
            I => data_in_frame_7_3
        );

    \I__5362\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28935\
        );

    \I__5361\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28932\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__28935\,
            I => \N__28929\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__28932\,
            I => \N__28926\
        );

    \I__5358\ : Span4Mux_v
    port map (
            O => \N__28929\,
            I => \N__28923\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__28926\,
            I => \c0.n2336\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__28923\,
            I => \c0.n2336\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__28918\,
            I => \N__28915\
        );

    \I__5354\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28912\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__28912\,
            I => \N__28909\
        );

    \I__5352\ : Span4Mux_h
    port map (
            O => \N__28909\,
            I => \N__28905\
        );

    \I__5351\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28902\
        );

    \I__5350\ : Span4Mux_h
    port map (
            O => \N__28905\,
            I => \N__28899\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__28902\,
            I => data_in_frame_7_5
        );

    \I__5348\ : Odrv4
    port map (
            O => \N__28899\,
            I => data_in_frame_7_5
        );

    \I__5347\ : InMux
    port map (
            O => \N__28894\,
            I => \N__28891\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__28891\,
            I => \N__28888\
        );

    \I__5345\ : Span4Mux_h
    port map (
            O => \N__28888\,
            I => \N__28884\
        );

    \I__5344\ : InMux
    port map (
            O => \N__28887\,
            I => \N__28881\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__28884\,
            I => \c0.n9541\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__28881\,
            I => \c0.n9541\
        );

    \I__5341\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28873\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__28873\,
            I => \N__28869\
        );

    \I__5339\ : InMux
    port map (
            O => \N__28872\,
            I => \N__28866\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__28869\,
            I => \N__28863\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__28866\,
            I => data_in_frame_6_0
        );

    \I__5336\ : Odrv4
    port map (
            O => \N__28863\,
            I => data_in_frame_6_0
        );

    \I__5335\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28855\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__28855\,
            I => \N__28852\
        );

    \I__5333\ : Span4Mux_h
    port map (
            O => \N__28852\,
            I => \N__28848\
        );

    \I__5332\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28845\
        );

    \I__5331\ : Span4Mux_h
    port map (
            O => \N__28848\,
            I => \N__28842\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__28845\,
            I => data_in_frame_6_5
        );

    \I__5329\ : Odrv4
    port map (
            O => \N__28842\,
            I => data_in_frame_6_5
        );

    \I__5328\ : CascadeMux
    port map (
            O => \N__28837\,
            I => \c0.n20_cascade_\
        );

    \I__5327\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28828\
        );

    \I__5326\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28828\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__28828\,
            I => \N__28824\
        );

    \I__5324\ : InMux
    port map (
            O => \N__28827\,
            I => \N__28821\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__28824\,
            I => \c0.n2342\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__28821\,
            I => \c0.n2342\
        );

    \I__5321\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28812\
        );

    \I__5320\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28809\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__28812\,
            I => \c0.data_in_frame_9_1\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__28809\,
            I => \c0.data_in_frame_9_1\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__28804\,
            I => \N__28792\
        );

    \I__5316\ : InMux
    port map (
            O => \N__28803\,
            I => \N__28789\
        );

    \I__5315\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28786\
        );

    \I__5314\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28782\
        );

    \I__5313\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28779\
        );

    \I__5312\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28770\
        );

    \I__5311\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28770\
        );

    \I__5310\ : InMux
    port map (
            O => \N__28797\,
            I => \N__28770\
        );

    \I__5309\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28770\
        );

    \I__5308\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28765\
        );

    \I__5307\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28765\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__28789\,
            I => \N__28755\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__28786\,
            I => \N__28755\
        );

    \I__5304\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28752\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__28782\,
            I => \N__28747\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__28779\,
            I => \N__28747\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__28770\,
            I => \N__28742\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__28765\,
            I => \N__28742\
        );

    \I__5299\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28739\
        );

    \I__5298\ : InMux
    port map (
            O => \N__28763\,
            I => \N__28736\
        );

    \I__5297\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28729\
        );

    \I__5296\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28729\
        );

    \I__5295\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28729\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__28755\,
            I => \N__28726\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28723\
        );

    \I__5292\ : Span4Mux_v
    port map (
            O => \N__28747\,
            I => \N__28718\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__28742\,
            I => \N__28718\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__28739\,
            I => \c0.n8_adj_2310\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__28736\,
            I => \c0.n8_adj_2310\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__28729\,
            I => \c0.n8_adj_2310\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__28726\,
            I => \c0.n8_adj_2310\
        );

    \I__5286\ : Odrv12
    port map (
            O => \N__28723\,
            I => \c0.n8_adj_2310\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__28718\,
            I => \c0.n8_adj_2310\
        );

    \I__5284\ : InMux
    port map (
            O => \N__28705\,
            I => \N__28699\
        );

    \I__5283\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28699\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__28699\,
            I => \c0.data_in_frame_9_5\
        );

    \I__5281\ : IoInMux
    port map (
            O => \N__28696\,
            I => \N__28693\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__5279\ : IoSpan4Mux
    port map (
            O => \N__28690\,
            I => \N__28686\
        );

    \I__5278\ : InMux
    port map (
            O => \N__28689\,
            I => \N__28683\
        );

    \I__5277\ : Sp12to4
    port map (
            O => \N__28686\,
            I => \N__28678\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__28683\,
            I => \N__28678\
        );

    \I__5275\ : Span12Mux_s6_h
    port map (
            O => \N__28678\,
            I => \N__28674\
        );

    \I__5274\ : InMux
    port map (
            O => \N__28677\,
            I => \N__28671\
        );

    \I__5273\ : Odrv12
    port map (
            O => \N__28674\,
            I => tx2_o
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__28671\,
            I => tx2_o
        );

    \I__5271\ : SRMux
    port map (
            O => \N__28666\,
            I => \N__28663\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28660\
        );

    \I__5269\ : Span4Mux_h
    port map (
            O => \N__28660\,
            I => \N__28657\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__28657\,
            I => \c0.n3_adj_2240\
        );

    \I__5267\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28651\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28646\
        );

    \I__5265\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28638\
        );

    \I__5264\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28638\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__28646\,
            I => \N__28635\
        );

    \I__5262\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28632\
        );

    \I__5261\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28627\
        );

    \I__5260\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28627\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__28638\,
            I => \N__28624\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__28635\,
            I => data_in_frame_0_7
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__28632\,
            I => data_in_frame_0_7
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__28627\,
            I => data_in_frame_0_7
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__28624\,
            I => data_in_frame_0_7
        );

    \I__5254\ : CascadeMux
    port map (
            O => \N__28615\,
            I => \N__28612\
        );

    \I__5253\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28607\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__28611\,
            I => \N__28604\
        );

    \I__5251\ : InMux
    port map (
            O => \N__28610\,
            I => \N__28600\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__28607\,
            I => \N__28597\
        );

    \I__5249\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28594\
        );

    \I__5248\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28591\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__28600\,
            I => \N__28586\
        );

    \I__5246\ : Span4Mux_v
    port map (
            O => \N__28597\,
            I => \N__28586\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__28594\,
            I => \c0.data_in_frame_1_7\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__28591\,
            I => \c0.data_in_frame_1_7\
        );

    \I__5243\ : Odrv4
    port map (
            O => \N__28586\,
            I => \c0.data_in_frame_1_7\
        );

    \I__5242\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28576\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__28576\,
            I => \N__28572\
        );

    \I__5240\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28569\
        );

    \I__5239\ : Span4Mux_v
    port map (
            O => \N__28572\,
            I => \N__28565\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__28569\,
            I => \N__28562\
        );

    \I__5237\ : InMux
    port map (
            O => \N__28568\,
            I => \N__28558\
        );

    \I__5236\ : Span4Mux_h
    port map (
            O => \N__28565\,
            I => \N__28555\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__28562\,
            I => \N__28552\
        );

    \I__5234\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28549\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__28558\,
            I => \c0.data_in_frame_1_4\
        );

    \I__5232\ : Odrv4
    port map (
            O => \N__28555\,
            I => \c0.data_in_frame_1_4\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__28552\,
            I => \c0.data_in_frame_1_4\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__28549\,
            I => \c0.data_in_frame_1_4\
        );

    \I__5229\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28537\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__28537\,
            I => \N__28534\
        );

    \I__5227\ : Span4Mux_v
    port map (
            O => \N__28534\,
            I => \N__28531\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__28531\,
            I => \c0.n27_adj_2342\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__28528\,
            I => \c0.n23_adj_2341_cascade_\
        );

    \I__5224\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28521\
        );

    \I__5223\ : CascadeMux
    port map (
            O => \N__28524\,
            I => \N__28518\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__28521\,
            I => \N__28515\
        );

    \I__5221\ : InMux
    port map (
            O => \N__28518\,
            I => \N__28510\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__28515\,
            I => \N__28507\
        );

    \I__5219\ : InMux
    port map (
            O => \N__28514\,
            I => \N__28502\
        );

    \I__5218\ : InMux
    port map (
            O => \N__28513\,
            I => \N__28502\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__28510\,
            I => \c0.data_in_frame_1_3\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__28507\,
            I => \c0.data_in_frame_1_3\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__28502\,
            I => \c0.data_in_frame_1_3\
        );

    \I__5214\ : InMux
    port map (
            O => \N__28495\,
            I => \N__28492\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__28492\,
            I => \N__28489\
        );

    \I__5212\ : Odrv12
    port map (
            O => \N__28489\,
            I => \c0.n21_adj_2171\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__28486\,
            I => \N__28483\
        );

    \I__5210\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28480\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__28480\,
            I => \N__28477\
        );

    \I__5208\ : Span4Mux_h
    port map (
            O => \N__28477\,
            I => \N__28474\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__28474\,
            I => \c0.n15930\
        );

    \I__5206\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28468\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__28468\,
            I => \N__28464\
        );

    \I__5204\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28461\
        );

    \I__5203\ : Span4Mux_h
    port map (
            O => \N__28464\,
            I => \N__28458\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__28461\,
            I => \c0.data_in_frame_10_7\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__28458\,
            I => \c0.data_in_frame_10_7\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__28453\,
            I => \c0.n17352_cascade_\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__28450\,
            I => \N__28447\
        );

    \I__5198\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28444\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__28444\,
            I => \c0.n27_adj_2196\
        );

    \I__5196\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28438\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__28438\,
            I => \N__28435\
        );

    \I__5194\ : Odrv12
    port map (
            O => \N__28435\,
            I => \c0.n25\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__28432\,
            I => \c0.n15846_cascade_\
        );

    \I__5192\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28426\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__28426\,
            I => \N__28423\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__28423\,
            I => \c0.n15929\
        );

    \I__5189\ : InMux
    port map (
            O => \N__28420\,
            I => \N__28417\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__28417\,
            I => \c0.n26_adj_2184\
        );

    \I__5187\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28411\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__28411\,
            I => \N__28408\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__28408\,
            I => \N__28405\
        );

    \I__5184\ : Odrv4
    port map (
            O => \N__28405\,
            I => \c0.n15938\
        );

    \I__5183\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28399\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__28399\,
            I => \N__28394\
        );

    \I__5181\ : InMux
    port map (
            O => \N__28398\,
            I => \N__28389\
        );

    \I__5180\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28386\
        );

    \I__5179\ : Span4Mux_v
    port map (
            O => \N__28394\,
            I => \N__28383\
        );

    \I__5178\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28380\
        );

    \I__5177\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28377\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__28389\,
            I => \N__28374\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__28386\,
            I => \c0.data_in_frame_1_2\
        );

    \I__5174\ : Odrv4
    port map (
            O => \N__28383\,
            I => \c0.data_in_frame_1_2\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__28380\,
            I => \c0.data_in_frame_1_2\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__28377\,
            I => \c0.data_in_frame_1_2\
        );

    \I__5171\ : Odrv4
    port map (
            O => \N__28374\,
            I => \c0.data_in_frame_1_2\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__28363\,
            I => \N__28360\
        );

    \I__5169\ : InMux
    port map (
            O => \N__28360\,
            I => \N__28357\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__28357\,
            I => \N__28353\
        );

    \I__5167\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28350\
        );

    \I__5166\ : Span4Mux_v
    port map (
            O => \N__28353\,
            I => \N__28347\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__28350\,
            I => \c0.data_in_frame_9_3\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__28347\,
            I => \c0.data_in_frame_9_3\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__28342\,
            I => \N__28339\
        );

    \I__5162\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28336\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__28336\,
            I => \N__28333\
        );

    \I__5160\ : Span4Mux_v
    port map (
            O => \N__28333\,
            I => \N__28330\
        );

    \I__5159\ : Span4Mux_h
    port map (
            O => \N__28330\,
            I => \N__28327\
        );

    \I__5158\ : Odrv4
    port map (
            O => \N__28327\,
            I => \c0.n8603\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__28324\,
            I => \N__28318\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__28323\,
            I => \N__28315\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__28322\,
            I => \N__28312\
        );

    \I__5154\ : InMux
    port map (
            O => \N__28321\,
            I => \N__28309\
        );

    \I__5153\ : InMux
    port map (
            O => \N__28318\,
            I => \N__28304\
        );

    \I__5152\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28304\
        );

    \I__5151\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28301\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__28309\,
            I => \N__28298\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__28304\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__28301\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__5147\ : Odrv12
    port map (
            O => \N__28298\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__5146\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28287\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__28290\,
            I => \N__28284\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__28287\,
            I => \N__28279\
        );

    \I__5143\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28274\
        );

    \I__5142\ : InMux
    port map (
            O => \N__28283\,
            I => \N__28274\
        );

    \I__5141\ : InMux
    port map (
            O => \N__28282\,
            I => \N__28271\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__28279\,
            I => \N__28268\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__28274\,
            I => \N__28261\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__28271\,
            I => \N__28261\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__28268\,
            I => \N__28261\
        );

    \I__5136\ : Odrv4
    port map (
            O => \N__28261\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__28258\,
            I => \N__28255\
        );

    \I__5134\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28251\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__28254\,
            I => \N__28246\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__28251\,
            I => \N__28243\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__28250\,
            I => \N__28240\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__28249\,
            I => \N__28237\
        );

    \I__5129\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28234\
        );

    \I__5128\ : Span4Mux_v
    port map (
            O => \N__28243\,
            I => \N__28231\
        );

    \I__5127\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28226\
        );

    \I__5126\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28226\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__28234\,
            I => \N__28223\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__28231\,
            I => \N__28220\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__28226\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__28223\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__28220\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__5120\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28210\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__28210\,
            I => \N__28207\
        );

    \I__5118\ : Odrv4
    port map (
            O => \N__28207\,
            I => \c0.n48\
        );

    \I__5117\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28201\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__28201\,
            I => \N__28198\
        );

    \I__5115\ : Span4Mux_h
    port map (
            O => \N__28198\,
            I => \N__28195\
        );

    \I__5114\ : Span4Mux_h
    port map (
            O => \N__28195\,
            I => \N__28192\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__28192\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_10\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__28189\,
            I => \N__28186\
        );

    \I__5111\ : InMux
    port map (
            O => \N__28186\,
            I => \N__28179\
        );

    \I__5110\ : InMux
    port map (
            O => \N__28185\,
            I => \N__28179\
        );

    \I__5109\ : InMux
    port map (
            O => \N__28184\,
            I => \N__28176\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__28179\,
            I => \N__28173\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__28176\,
            I => \N__28170\
        );

    \I__5106\ : Sp12to4
    port map (
            O => \N__28173\,
            I => \N__28164\
        );

    \I__5105\ : Span12Mux_s10_v
    port map (
            O => \N__28170\,
            I => \N__28164\
        );

    \I__5104\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28161\
        );

    \I__5103\ : Odrv12
    port map (
            O => \N__28164\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__28161\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__5101\ : SRMux
    port map (
            O => \N__28156\,
            I => \N__28153\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__28153\,
            I => \N__28150\
        );

    \I__5099\ : Span4Mux_h
    port map (
            O => \N__28150\,
            I => \N__28147\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__28147\,
            I => \c0.n3_adj_2247\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__28144\,
            I => \c0.n9819_cascade_\
        );

    \I__5096\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28136\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28133\
        );

    \I__5094\ : InMux
    port map (
            O => \N__28139\,
            I => \N__28129\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__28136\,
            I => \N__28126\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28123\
        );

    \I__5091\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28120\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__28129\,
            I => \N__28117\
        );

    \I__5089\ : Span4Mux_h
    port map (
            O => \N__28126\,
            I => \N__28114\
        );

    \I__5088\ : Span4Mux_h
    port map (
            O => \N__28123\,
            I => \N__28111\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__28120\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__5086\ : Odrv4
    port map (
            O => \N__28117\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__28114\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__28111\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__5083\ : SRMux
    port map (
            O => \N__28102\,
            I => \N__28099\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__28099\,
            I => \N__28096\
        );

    \I__5081\ : Odrv12
    port map (
            O => \N__28096\,
            I => \c0.n16359\
        );

    \I__5080\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28090\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__28090\,
            I => \N__28087\
        );

    \I__5078\ : Odrv12
    port map (
            O => \N__28087\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_17\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__28084\,
            I => \N__28078\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__28083\,
            I => \N__28075\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__28082\,
            I => \N__28072\
        );

    \I__5074\ : InMux
    port map (
            O => \N__28081\,
            I => \N__28069\
        );

    \I__5073\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28066\
        );

    \I__5072\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28063\
        );

    \I__5071\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28060\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28057\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__28066\,
            I => \N__28054\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__28063\,
            I => \N__28049\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__28060\,
            I => \N__28049\
        );

    \I__5066\ : Span4Mux_h
    port map (
            O => \N__28057\,
            I => \N__28046\
        );

    \I__5065\ : Span4Mux_h
    port map (
            O => \N__28054\,
            I => \N__28043\
        );

    \I__5064\ : Odrv12
    port map (
            O => \N__28049\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__5063\ : Odrv4
    port map (
            O => \N__28046\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__28043\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__5061\ : InMux
    port map (
            O => \N__28036\,
            I => \N__28033\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__28033\,
            I => \N__28030\
        );

    \I__5059\ : Span4Mux_h
    port map (
            O => \N__28030\,
            I => \N__28026\
        );

    \I__5058\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28023\
        );

    \I__5057\ : Span4Mux_h
    port map (
            O => \N__28026\,
            I => \N__28020\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__28023\,
            I => \N__28017\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__28020\,
            I => n17
        );

    \I__5054\ : Odrv4
    port map (
            O => \N__28017\,
            I => n17
        );

    \I__5053\ : SRMux
    port map (
            O => \N__28012\,
            I => \N__28009\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__28009\,
            I => \N__28006\
        );

    \I__5051\ : Span4Mux_h
    port map (
            O => \N__28006\,
            I => \N__28003\
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__28003\,
            I => \c0.n16369\
        );

    \I__5049\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27997\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__27997\,
            I => \N__27994\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__27994\,
            I => \c0.n12_adj_2189\
        );

    \I__5046\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27987\
        );

    \I__5045\ : InMux
    port map (
            O => \N__27990\,
            I => \N__27984\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__27987\,
            I => \N__27978\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27975\
        );

    \I__5042\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27972\
        );

    \I__5041\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27969\
        );

    \I__5040\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27966\
        );

    \I__5039\ : Span4Mux_v
    port map (
            O => \N__27978\,
            I => \N__27963\
        );

    \I__5038\ : Span4Mux_h
    port map (
            O => \N__27975\,
            I => \N__27958\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__27972\,
            I => \N__27958\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__27969\,
            I => \N__27955\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__27966\,
            I => \N__27948\
        );

    \I__5034\ : Span4Mux_h
    port map (
            O => \N__27963\,
            I => \N__27948\
        );

    \I__5033\ : Span4Mux_v
    port map (
            O => \N__27958\,
            I => \N__27948\
        );

    \I__5032\ : Odrv12
    port map (
            O => \N__27955\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__27948\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__5030\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27940\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__27940\,
            I => \N__27934\
        );

    \I__5028\ : InMux
    port map (
            O => \N__27939\,
            I => \N__27931\
        );

    \I__5027\ : InMux
    port map (
            O => \N__27938\,
            I => \N__27926\
        );

    \I__5026\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27926\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__27934\,
            I => \N__27923\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27920\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27917\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__27923\,
            I => n9460
        );

    \I__5021\ : Odrv12
    port map (
            O => \N__27920\,
            I => n9460
        );

    \I__5020\ : Odrv12
    port map (
            O => \N__27917\,
            I => n9460
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__27910\,
            I => \n9460_cascade_\
        );

    \I__5018\ : InMux
    port map (
            O => \N__27907\,
            I => \N__27903\
        );

    \I__5017\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27900\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__27903\,
            I => \N__27897\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__27900\,
            I => \N__27894\
        );

    \I__5014\ : Span4Mux_h
    port map (
            O => \N__27897\,
            I => \N__27891\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__27894\,
            I => \N__27888\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__27891\,
            I => \N__27885\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__27888\,
            I => n9462
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__27885\,
            I => n9462
        );

    \I__5009\ : InMux
    port map (
            O => \N__27880\,
            I => \N__27875\
        );

    \I__5008\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27872\
        );

    \I__5007\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27869\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__27875\,
            I => \N__27866\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__27872\,
            I => \N__27861\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__27869\,
            I => \N__27856\
        );

    \I__5003\ : Span4Mux_v
    port map (
            O => \N__27866\,
            I => \N__27856\
        );

    \I__5002\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27851\
        );

    \I__5001\ : InMux
    port map (
            O => \N__27864\,
            I => \N__27851\
        );

    \I__5000\ : Span4Mux_h
    port map (
            O => \N__27861\,
            I => \N__27848\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__27856\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__27851\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__27848\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__4996\ : SRMux
    port map (
            O => \N__27841\,
            I => \N__27838\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__27838\,
            I => \c0.n16343\
        );

    \I__4994\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27832\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__4992\ : Span4Mux_v
    port map (
            O => \N__27829\,
            I => \N__27825\
        );

    \I__4991\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27821\
        );

    \I__4990\ : Span4Mux_h
    port map (
            O => \N__27825\,
            I => \N__27818\
        );

    \I__4989\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27815\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__27821\,
            I => data_in_2_6
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__27818\,
            I => data_in_2_6
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__27815\,
            I => data_in_2_6
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__4984\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27791\
        );

    \I__4983\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27791\
        );

    \I__4982\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27791\
        );

    \I__4981\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27791\
        );

    \I__4980\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27787\
        );

    \I__4979\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27784\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__27791\,
            I => \N__27779\
        );

    \I__4977\ : InMux
    port map (
            O => \N__27790\,
            I => \N__27776\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__27787\,
            I => \N__27771\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__27784\,
            I => \N__27771\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__27783\,
            I => \N__27765\
        );

    \I__4973\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27758\
        );

    \I__4972\ : Span4Mux_v
    port map (
            O => \N__27779\,
            I => \N__27753\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__27776\,
            I => \N__27753\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__27771\,
            I => \N__27750\
        );

    \I__4969\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27747\
        );

    \I__4968\ : InMux
    port map (
            O => \N__27769\,
            I => \N__27736\
        );

    \I__4967\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27736\
        );

    \I__4966\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27731\
        );

    \I__4965\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27731\
        );

    \I__4964\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27724\
        );

    \I__4963\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27724\
        );

    \I__4962\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27724\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__27758\,
            I => \N__27721\
        );

    \I__4960\ : Span4Mux_h
    port map (
            O => \N__27753\,
            I => \N__27714\
        );

    \I__4959\ : Span4Mux_v
    port map (
            O => \N__27750\,
            I => \N__27714\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__27747\,
            I => \N__27714\
        );

    \I__4957\ : InMux
    port map (
            O => \N__27746\,
            I => \N__27695\
        );

    \I__4956\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27695\
        );

    \I__4955\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27695\
        );

    \I__4954\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27695\
        );

    \I__4953\ : InMux
    port map (
            O => \N__27742\,
            I => \N__27690\
        );

    \I__4952\ : InMux
    port map (
            O => \N__27741\,
            I => \N__27690\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__27736\,
            I => \N__27687\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__27731\,
            I => \N__27680\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__27724\,
            I => \N__27680\
        );

    \I__4948\ : Span4Mux_v
    port map (
            O => \N__27721\,
            I => \N__27680\
        );

    \I__4947\ : Span4Mux_h
    port map (
            O => \N__27714\,
            I => \N__27677\
        );

    \I__4946\ : CascadeMux
    port map (
            O => \N__27713\,
            I => \N__27674\
        );

    \I__4945\ : InMux
    port map (
            O => \N__27712\,
            I => \N__27666\
        );

    \I__4944\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27666\
        );

    \I__4943\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27657\
        );

    \I__4942\ : InMux
    port map (
            O => \N__27709\,
            I => \N__27657\
        );

    \I__4941\ : InMux
    port map (
            O => \N__27708\,
            I => \N__27657\
        );

    \I__4940\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27657\
        );

    \I__4939\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27650\
        );

    \I__4938\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27650\
        );

    \I__4937\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27650\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__27695\,
            I => \N__27647\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__27690\,
            I => \N__27644\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__27687\,
            I => \N__27641\
        );

    \I__4933\ : Span4Mux_h
    port map (
            O => \N__27680\,
            I => \N__27636\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__27677\,
            I => \N__27636\
        );

    \I__4931\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27627\
        );

    \I__4930\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27627\
        );

    \I__4929\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27627\
        );

    \I__4928\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27627\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__27666\,
            I => rx_data_ready
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__27657\,
            I => rx_data_ready
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__27650\,
            I => rx_data_ready
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__27647\,
            I => rx_data_ready
        );

    \I__4923\ : Odrv12
    port map (
            O => \N__27644\,
            I => rx_data_ready
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__27641\,
            I => rx_data_ready
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__27636\,
            I => rx_data_ready
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__27627\,
            I => rx_data_ready
        );

    \I__4919\ : InMux
    port map (
            O => \N__27610\,
            I => \N__27605\
        );

    \I__4918\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27600\
        );

    \I__4917\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27600\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__27605\,
            I => \N__27597\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__27600\,
            I => \N__27593\
        );

    \I__4914\ : Span12Mux_s8_h
    port map (
            O => \N__27597\,
            I => \N__27590\
        );

    \I__4913\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27587\
        );

    \I__4912\ : Span4Mux_h
    port map (
            O => \N__27593\,
            I => \N__27584\
        );

    \I__4911\ : Odrv12
    port map (
            O => \N__27590\,
            I => data_in_1_6
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__27587\,
            I => data_in_1_6
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__27584\,
            I => data_in_1_6
        );

    \I__4908\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27570\
        );

    \I__4907\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27565\
        );

    \I__4906\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27560\
        );

    \I__4905\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27560\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__27573\,
            I => \N__27553\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__27570\,
            I => \N__27545\
        );

    \I__4902\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27540\
        );

    \I__4901\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27540\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N__27535\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__27560\,
            I => \N__27535\
        );

    \I__4898\ : InMux
    port map (
            O => \N__27559\,
            I => \N__27529\
        );

    \I__4897\ : InMux
    port map (
            O => \N__27558\,
            I => \N__27520\
        );

    \I__4896\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27520\
        );

    \I__4895\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27520\
        );

    \I__4894\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27520\
        );

    \I__4893\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27515\
        );

    \I__4892\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27515\
        );

    \I__4891\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27510\
        );

    \I__4890\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27510\
        );

    \I__4889\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27507\
        );

    \I__4888\ : Span4Mux_v
    port map (
            O => \N__27545\,
            I => \N__27500\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__27540\,
            I => \N__27500\
        );

    \I__4886\ : Span4Mux_s1_v
    port map (
            O => \N__27535\,
            I => \N__27500\
        );

    \I__4885\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27495\
        );

    \I__4884\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27495\
        );

    \I__4883\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27492\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__27529\,
            I => n29
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__27520\,
            I => n29
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__27515\,
            I => n29
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__27510\,
            I => n29
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__27507\,
            I => n29
        );

    \I__4877\ : Odrv4
    port map (
            O => \N__27500\,
            I => n29
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__27495\,
            I => n29
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__27492\,
            I => n29
        );

    \I__4874\ : CascadeMux
    port map (
            O => \N__27475\,
            I => \N__27472\
        );

    \I__4873\ : InMux
    port map (
            O => \N__27472\,
            I => \N__27468\
        );

    \I__4872\ : InMux
    port map (
            O => \N__27471\,
            I => \N__27465\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__27468\,
            I => \N__27461\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__27465\,
            I => \N__27458\
        );

    \I__4869\ : CascadeMux
    port map (
            O => \N__27464\,
            I => \N__27455\
        );

    \I__4868\ : Span4Mux_s3_v
    port map (
            O => \N__27461\,
            I => \N__27452\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__27458\,
            I => \N__27449\
        );

    \I__4866\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27446\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__27452\,
            I => \N__27443\
        );

    \I__4864\ : Sp12to4
    port map (
            O => \N__27449\,
            I => \N__27438\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27438\
        );

    \I__4862\ : Span4Mux_v
    port map (
            O => \N__27443\,
            I => \N__27435\
        );

    \I__4861\ : Span12Mux_s10_v
    port map (
            O => \N__27438\,
            I => \N__27432\
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__27435\,
            I => n445
        );

    \I__4859\ : Odrv12
    port map (
            O => \N__27432\,
            I => n445
        );

    \I__4858\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27422\
        );

    \I__4857\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27417\
        );

    \I__4856\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27417\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__27422\,
            I => n10031
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__27417\,
            I => n10031
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__27412\,
            I => \n17479_cascade_\
        );

    \I__4852\ : InMux
    port map (
            O => \N__27409\,
            I => \N__27406\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__27406\,
            I => \N__27403\
        );

    \I__4850\ : Span4Mux_h
    port map (
            O => \N__27403\,
            I => \N__27399\
        );

    \I__4849\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27396\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__27399\,
            I => n16886
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__27396\,
            I => n16886
        );

    \I__4846\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27388\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__27388\,
            I => n38
        );

    \I__4844\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27382\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__27382\,
            I => \c0.n44_adj_2163\
        );

    \I__4842\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27366\
        );

    \I__4841\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27366\
        );

    \I__4840\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27366\
        );

    \I__4839\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27366\
        );

    \I__4838\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27363\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__27366\,
            I => n9357
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__27363\,
            I => n9357
        );

    \I__4835\ : CascadeMux
    port map (
            O => \N__27358\,
            I => \N__27354\
        );

    \I__4834\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27349\
        );

    \I__4833\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27344\
        );

    \I__4832\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27339\
        );

    \I__4831\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27339\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__27349\,
            I => \N__27335\
        );

    \I__4829\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27330\
        );

    \I__4828\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27330\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__27344\,
            I => \N__27325\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__27339\,
            I => \N__27325\
        );

    \I__4825\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27322\
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__27335\,
            I => \c0.tx_transmit_N_1949_2\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__27330\,
            I => \c0.tx_transmit_N_1949_2\
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__27325\,
            I => \c0.tx_transmit_N_1949_2\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__27322\,
            I => \c0.tx_transmit_N_1949_2\
        );

    \I__4820\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27303\
        );

    \I__4819\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27303\
        );

    \I__4818\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27300\
        );

    \I__4817\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27297\
        );

    \I__4816\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27294\
        );

    \I__4815\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27291\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__27303\,
            I => \c0.n4_adj_2311\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__27300\,
            I => \c0.n4_adj_2311\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__27297\,
            I => \c0.n4_adj_2311\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__27294\,
            I => \c0.n4_adj_2311\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__27291\,
            I => \c0.n4_adj_2311\
        );

    \I__4809\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27277\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__27277\,
            I => \N__27274\
        );

    \I__4807\ : Odrv12
    port map (
            O => \N__27274\,
            I => \c0.n17475\
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__27271\,
            I => \c0.tx2_transmit_N_1997_cascade_\
        );

    \I__4805\ : InMux
    port map (
            O => \N__27268\,
            I => \N__27265\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__27265\,
            I => \c0.tx2.n113\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__27262\,
            I => \c0.tx2.n113_cascade_\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__27259\,
            I => \N__27256\
        );

    \I__4801\ : InMux
    port map (
            O => \N__27256\,
            I => \N__27253\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__27253\,
            I => \N__27250\
        );

    \I__4799\ : Span4Mux_v
    port map (
            O => \N__27250\,
            I => \N__27245\
        );

    \I__4798\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27242\
        );

    \I__4797\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27239\
        );

    \I__4796\ : Span4Mux_h
    port map (
            O => \N__27245\,
            I => \N__27236\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__27242\,
            I => \N__27231\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__27239\,
            I => \N__27231\
        );

    \I__4793\ : Span4Mux_h
    port map (
            O => \N__27236\,
            I => \N__27226\
        );

    \I__4792\ : Span12Mux_v
    port map (
            O => \N__27231\,
            I => \N__27223\
        );

    \I__4791\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27218\
        );

    \I__4790\ : InMux
    port map (
            O => \N__27229\,
            I => \N__27218\
        );

    \I__4789\ : Span4Mux_v
    port map (
            O => \N__27226\,
            I => \N__27215\
        );

    \I__4788\ : Odrv12
    port map (
            O => \N__27223\,
            I => \c0.r_SM_Main_2_N_2036_0_adj_2261\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__27218\,
            I => \c0.r_SM_Main_2_N_2036_0_adj_2261\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__27215\,
            I => \c0.r_SM_Main_2_N_2036_0_adj_2261\
        );

    \I__4785\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27205\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__27205\,
            I => \N__27202\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__27202\,
            I => \N__27199\
        );

    \I__4782\ : Odrv4
    port map (
            O => \N__27199\,
            I => n491
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__27196\,
            I => \n491_cascade_\
        );

    \I__4780\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27190\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__27190\,
            I => \N__27185\
        );

    \I__4778\ : InMux
    port map (
            O => \N__27189\,
            I => \N__27182\
        );

    \I__4777\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27179\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__27185\,
            I => \c0.n8938\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__27182\,
            I => \c0.n8938\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__27179\,
            I => \c0.n8938\
        );

    \I__4773\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27165\
        );

    \I__4772\ : InMux
    port map (
            O => \N__27171\,
            I => \N__27160\
        );

    \I__4771\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27160\
        );

    \I__4770\ : InMux
    port map (
            O => \N__27169\,
            I => \N__27155\
        );

    \I__4769\ : InMux
    port map (
            O => \N__27168\,
            I => \N__27155\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__27165\,
            I => \c0.tx_transmit_N_1949_3\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__27160\,
            I => \c0.tx_transmit_N_1949_3\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__27155\,
            I => \c0.tx_transmit_N_1949_3\
        );

    \I__4765\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27135\
        );

    \I__4764\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27135\
        );

    \I__4763\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27135\
        );

    \I__4762\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27132\
        );

    \I__4761\ : InMux
    port map (
            O => \N__27144\,
            I => \N__27125\
        );

    \I__4760\ : InMux
    port map (
            O => \N__27143\,
            I => \N__27125\
        );

    \I__4759\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27125\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__27135\,
            I => \c0.n16839\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__27132\,
            I => \c0.n16839\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__27125\,
            I => \c0.n16839\
        );

    \I__4755\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27114\
        );

    \I__4754\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27111\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__27114\,
            I => \c0.tx_transmit_N_1949_7\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__27111\,
            I => \c0.tx_transmit_N_1949_7\
        );

    \I__4751\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27102\
        );

    \I__4750\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27099\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__27102\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__27099\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__27094\,
            I => \n17834_cascade_\
        );

    \I__4746\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27088\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__27088\,
            I => n17162
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__27085\,
            I => \n9358_cascade_\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__27082\,
            I => \n41_cascade_\
        );

    \I__4742\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27076\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__27076\,
            I => n35
        );

    \I__4740\ : InMux
    port map (
            O => \N__27073\,
            I => \N__27070\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__27070\,
            I => \c0.n17254\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__27067\,
            I => \c0.n17254_cascade_\
        );

    \I__4737\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27061\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__27061\,
            I => \N__27058\
        );

    \I__4735\ : Span4Mux_s2_v
    port map (
            O => \N__27058\,
            I => \N__27055\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__27055\,
            I => \c0.n17290\
        );

    \I__4733\ : CascadeMux
    port map (
            O => \N__27052\,
            I => \N__27049\
        );

    \I__4732\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27043\
        );

    \I__4731\ : InMux
    port map (
            O => \N__27048\,
            I => \N__27043\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__27043\,
            I => \c0.tx_transmit_N_1949_5\
        );

    \I__4729\ : InMux
    port map (
            O => \N__27040\,
            I => \N__27036\
        );

    \I__4728\ : InMux
    port map (
            O => \N__27039\,
            I => \N__27033\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__27036\,
            I => \c0.n5_adj_2319\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__27033\,
            I => \c0.n5_adj_2319\
        );

    \I__4725\ : InMux
    port map (
            O => \N__27028\,
            I => \N__27021\
        );

    \I__4724\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27021\
        );

    \I__4723\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27018\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__27021\,
            I => \c0.tx_transmit_N_1949_6\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__27018\,
            I => \c0.tx_transmit_N_1949_6\
        );

    \I__4720\ : InMux
    port map (
            O => \N__27013\,
            I => \N__27009\
        );

    \I__4719\ : InMux
    port map (
            O => \N__27012\,
            I => \N__27006\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__27009\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__27006\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__4716\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26998\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__26998\,
            I => \c0.n23_adj_2309\
        );

    \I__4714\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26992\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__26992\,
            I => \N__26989\
        );

    \I__4712\ : Odrv12
    port map (
            O => \N__26989\,
            I => \c0.n17278\
        );

    \I__4711\ : InMux
    port map (
            O => \N__26986\,
            I => \N__26983\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__26983\,
            I => \N__26980\
        );

    \I__4709\ : Span4Mux_s2_v
    port map (
            O => \N__26980\,
            I => \N__26977\
        );

    \I__4708\ : Odrv4
    port map (
            O => \N__26977\,
            I => \c0.n17276\
        );

    \I__4707\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26970\
        );

    \I__4706\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26967\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__26970\,
            I => \c0.tx_transmit_N_1949_0\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__26967\,
            I => \c0.tx_transmit_N_1949_0\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__26962\,
            I => \c0.n16839_cascade_\
        );

    \I__4702\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26954\
        );

    \I__4701\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26951\
        );

    \I__4700\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26948\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__26954\,
            I => \c0.tx_transmit_N_1949_4\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__26951\,
            I => \c0.tx_transmit_N_1949_4\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__26948\,
            I => \c0.tx_transmit_N_1949_4\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__26941\,
            I => \N__26937\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__26940\,
            I => \N__26933\
        );

    \I__4694\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26929\
        );

    \I__4693\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26926\
        );

    \I__4692\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26923\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__26932\,
            I => \N__26920\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__26929\,
            I => \N__26915\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__26926\,
            I => \N__26912\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__26923\,
            I => \N__26907\
        );

    \I__4687\ : InMux
    port map (
            O => \N__26920\,
            I => \N__26902\
        );

    \I__4686\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26902\
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__26918\,
            I => \N__26898\
        );

    \I__4684\ : Span4Mux_v
    port map (
            O => \N__26915\,
            I => \N__26895\
        );

    \I__4683\ : Span4Mux_h
    port map (
            O => \N__26912\,
            I => \N__26892\
        );

    \I__4682\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26889\
        );

    \I__4681\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26886\
        );

    \I__4680\ : Span4Mux_h
    port map (
            O => \N__26907\,
            I => \N__26881\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__26902\,
            I => \N__26881\
        );

    \I__4678\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26878\
        );

    \I__4677\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26875\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__26895\,
            I => rx_data_2
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__26892\,
            I => rx_data_2
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__26889\,
            I => rx_data_2
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__26886\,
            I => rx_data_2
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__26881\,
            I => rx_data_2
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__26878\,
            I => rx_data_2
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__26875\,
            I => rx_data_2
        );

    \I__4669\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26853\
        );

    \I__4668\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26853\
        );

    \I__4667\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26848\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__26853\,
            I => \N__26845\
        );

    \I__4665\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26840\
        );

    \I__4664\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26840\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__26848\,
            I => data_in_frame_0_0
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__26845\,
            I => data_in_frame_0_0
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__26840\,
            I => data_in_frame_0_0
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__26833\,
            I => \N__26828\
        );

    \I__4659\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26825\
        );

    \I__4658\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26821\
        );

    \I__4657\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26817\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__26825\,
            I => \N__26814\
        );

    \I__4655\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26811\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__26821\,
            I => \N__26808\
        );

    \I__4653\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26805\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__26817\,
            I => \c0.data_in_frame_1_6\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__26814\,
            I => \c0.data_in_frame_1_6\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__26811\,
            I => \c0.data_in_frame_1_6\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__26808\,
            I => \c0.data_in_frame_1_6\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__26805\,
            I => \c0.data_in_frame_1_6\
        );

    \I__4647\ : CascadeMux
    port map (
            O => \N__26794\,
            I => \N__26790\
        );

    \I__4646\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26785\
        );

    \I__4645\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26785\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__26785\,
            I => \c0.data_in_frame_10_2\
        );

    \I__4643\ : InMux
    port map (
            O => \N__26782\,
            I => \N__26775\
        );

    \I__4642\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26775\
        );

    \I__4641\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26770\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__26775\,
            I => \N__26767\
        );

    \I__4639\ : InMux
    port map (
            O => \N__26774\,
            I => \N__26762\
        );

    \I__4638\ : InMux
    port map (
            O => \N__26773\,
            I => \N__26762\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__26770\,
            I => data_in_frame_0_1
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__26767\,
            I => data_in_frame_0_1
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__26762\,
            I => data_in_frame_0_1
        );

    \I__4634\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26752\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__26752\,
            I => \c0.n17460\
        );

    \I__4632\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26746\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26742\
        );

    \I__4630\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26739\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__26742\,
            I => \r_Tx_Data_3\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__26739\,
            I => \r_Tx_Data_3\
        );

    \I__4627\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26729\
        );

    \I__4626\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26726\
        );

    \I__4625\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26722\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__26729\,
            I => \N__26719\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__26726\,
            I => \N__26716\
        );

    \I__4622\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26713\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__26722\,
            I => \c0.delay_counter_13\
        );

    \I__4620\ : Odrv12
    port map (
            O => \N__26719\,
            I => \c0.delay_counter_13\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__26716\,
            I => \c0.delay_counter_13\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__26713\,
            I => \c0.delay_counter_13\
        );

    \I__4617\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26700\
        );

    \I__4616\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26695\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__26700\,
            I => \N__26692\
        );

    \I__4614\ : InMux
    port map (
            O => \N__26699\,
            I => \N__26689\
        );

    \I__4613\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26686\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__26695\,
            I => \N__26679\
        );

    \I__4611\ : Span4Mux_h
    port map (
            O => \N__26692\,
            I => \N__26679\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__26689\,
            I => \N__26679\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__26686\,
            I => \c0.delay_counter_8\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__26679\,
            I => \c0.delay_counter_8\
        );

    \I__4607\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26671\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__26671\,
            I => \N__26665\
        );

    \I__4605\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26662\
        );

    \I__4604\ : InMux
    port map (
            O => \N__26669\,
            I => \N__26657\
        );

    \I__4603\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26657\
        );

    \I__4602\ : Odrv12
    port map (
            O => \N__26665\,
            I => \c0.delay_counter_4\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__26662\,
            I => \c0.delay_counter_4\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__26657\,
            I => \c0.delay_counter_4\
        );

    \I__4599\ : CascadeMux
    port map (
            O => \N__26650\,
            I => \N__26646\
        );

    \I__4598\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26642\
        );

    \I__4597\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26639\
        );

    \I__4596\ : InMux
    port map (
            O => \N__26645\,
            I => \N__26636\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__26642\,
            I => \N__26632\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__26639\,
            I => \N__26627\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__26636\,
            I => \N__26627\
        );

    \I__4592\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26624\
        );

    \I__4591\ : Span4Mux_s1_v
    port map (
            O => \N__26632\,
            I => \N__26621\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__26627\,
            I => \c0.delay_counter_2\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__26624\,
            I => \c0.delay_counter_2\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__26621\,
            I => \c0.delay_counter_2\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__26614\,
            I => \N__26611\
        );

    \I__4586\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26608\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__26608\,
            I => \N__26605\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__26605\,
            I => \c0.n17236\
        );

    \I__4583\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26599\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__26599\,
            I => \c0.n42_adj_2165\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__26596\,
            I => \N__26592\
        );

    \I__4580\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26589\
        );

    \I__4579\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26586\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__26589\,
            I => \c0.byte_transmit_counter_5\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__26586\,
            I => \c0.byte_transmit_counter_5\
        );

    \I__4576\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26574\
        );

    \I__4574\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26571\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__26574\,
            I => \N__26568\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__26571\,
            I => data_in_frame_7_2
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__26568\,
            I => data_in_frame_7_2
        );

    \I__4570\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26559\
        );

    \I__4569\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26556\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__26559\,
            I => \N__26553\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__26556\,
            I => data_in_frame_6_2
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__26553\,
            I => data_in_frame_6_2
        );

    \I__4565\ : CascadeMux
    port map (
            O => \N__26548\,
            I => \c0.n22_cascade_\
        );

    \I__4564\ : InMux
    port map (
            O => \N__26545\,
            I => \N__26542\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__26542\,
            I => \c0.n27\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__26539\,
            I => \N__26533\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__26538\,
            I => \N__26529\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__26537\,
            I => \N__26526\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__26536\,
            I => \N__26522\
        );

    \I__4558\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26517\
        );

    \I__4557\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26514\
        );

    \I__4556\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26511\
        );

    \I__4555\ : InMux
    port map (
            O => \N__26526\,
            I => \N__26508\
        );

    \I__4554\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26505\
        );

    \I__4553\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26502\
        );

    \I__4552\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26499\
        );

    \I__4551\ : InMux
    port map (
            O => \N__26520\,
            I => \N__26496\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__26517\,
            I => \N__26491\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__26514\,
            I => \N__26491\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__26511\,
            I => \N__26485\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__26508\,
            I => \N__26485\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__26505\,
            I => \N__26482\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__26502\,
            I => \N__26477\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__26499\,
            I => \N__26477\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__26496\,
            I => \N__26474\
        );

    \I__4542\ : Span4Mux_v
    port map (
            O => \N__26491\,
            I => \N__26471\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__26490\,
            I => \N__26468\
        );

    \I__4540\ : Span4Mux_v
    port map (
            O => \N__26485\,
            I => \N__26465\
        );

    \I__4539\ : Span4Mux_h
    port map (
            O => \N__26482\,
            I => \N__26462\
        );

    \I__4538\ : Span12Mux_h
    port map (
            O => \N__26477\,
            I => \N__26459\
        );

    \I__4537\ : Span4Mux_v
    port map (
            O => \N__26474\,
            I => \N__26456\
        );

    \I__4536\ : Span4Mux_s3_h
    port map (
            O => \N__26471\,
            I => \N__26453\
        );

    \I__4535\ : InMux
    port map (
            O => \N__26468\,
            I => \N__26450\
        );

    \I__4534\ : Odrv4
    port map (
            O => \N__26465\,
            I => rx_data_7
        );

    \I__4533\ : Odrv4
    port map (
            O => \N__26462\,
            I => rx_data_7
        );

    \I__4532\ : Odrv12
    port map (
            O => \N__26459\,
            I => rx_data_7
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__26456\,
            I => rx_data_7
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__26453\,
            I => rx_data_7
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__26450\,
            I => rx_data_7
        );

    \I__4528\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26432\
        );

    \I__4527\ : CascadeMux
    port map (
            O => \N__26436\,
            I => \N__26429\
        );

    \I__4526\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26425\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__26432\,
            I => \N__26422\
        );

    \I__4524\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26419\
        );

    \I__4523\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26416\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__26425\,
            I => \N__26413\
        );

    \I__4521\ : Span4Mux_h
    port map (
            O => \N__26422\,
            I => \N__26410\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__26419\,
            I => \c0.data_in_frame_1_0\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__26416\,
            I => \c0.data_in_frame_1_0\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__26413\,
            I => \c0.data_in_frame_1_0\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__26410\,
            I => \c0.data_in_frame_1_0\
        );

    \I__4516\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26398\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__26398\,
            I => \N__26395\
        );

    \I__4514\ : Odrv12
    port map (
            O => \N__26395\,
            I => n17634
        );

    \I__4513\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26383\
        );

    \I__4512\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26383\
        );

    \I__4511\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26383\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__26383\,
            I => \N__26379\
        );

    \I__4509\ : InMux
    port map (
            O => \N__26382\,
            I => \N__26375\
        );

    \I__4508\ : Span4Mux_s3_h
    port map (
            O => \N__26379\,
            I => \N__26372\
        );

    \I__4507\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26369\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__26375\,
            I => \N__26366\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__26372\,
            I => \N__26363\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__26369\,
            I => \r_Clock_Count_6_adj_2448\
        );

    \I__4503\ : Odrv12
    port map (
            O => \N__26366\,
            I => \r_Clock_Count_6_adj_2448\
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__26363\,
            I => \r_Clock_Count_6_adj_2448\
        );

    \I__4501\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26353\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__26353\,
            I => \c0.n9585\
        );

    \I__4499\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26346\
        );

    \I__4498\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26343\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26340\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__26343\,
            I => \c0.data_in_frame_2_2\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__26340\,
            I => \c0.data_in_frame_2_2\
        );

    \I__4494\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26332\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__26332\,
            I => \c0.n22_adj_2301\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__26329\,
            I => \c0.n9585_cascade_\
        );

    \I__4491\ : InMux
    port map (
            O => \N__26326\,
            I => \N__26323\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__26323\,
            I => \N__26319\
        );

    \I__4489\ : InMux
    port map (
            O => \N__26322\,
            I => \N__26316\
        );

    \I__4488\ : Sp12to4
    port map (
            O => \N__26319\,
            I => \N__26313\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__26316\,
            I => data_in_frame_7_1
        );

    \I__4486\ : Odrv12
    port map (
            O => \N__26313\,
            I => data_in_frame_7_1
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__26308\,
            I => \N__26305\
        );

    \I__4484\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26301\
        );

    \I__4483\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26298\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__26301\,
            I => \N__26295\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__26298\,
            I => \N__26290\
        );

    \I__4480\ : Span4Mux_v
    port map (
            O => \N__26295\,
            I => \N__26290\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__26290\,
            I => data_in_frame_7_4
        );

    \I__4478\ : InMux
    port map (
            O => \N__26287\,
            I => \N__26283\
        );

    \I__4477\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26280\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__26283\,
            I => \N__26277\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__26280\,
            I => \c0.data_in_frame_2_5\
        );

    \I__4474\ : Odrv12
    port map (
            O => \N__26277\,
            I => \c0.data_in_frame_2_5\
        );

    \I__4473\ : InMux
    port map (
            O => \N__26272\,
            I => \N__26268\
        );

    \I__4472\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26265\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__26268\,
            I => \N__26262\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__26265\,
            I => \c0.data_in_frame_2_3\
        );

    \I__4469\ : Odrv4
    port map (
            O => \N__26262\,
            I => \c0.data_in_frame_2_3\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__26257\,
            I => \c0.n2336_cascade_\
        );

    \I__4467\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26250\
        );

    \I__4466\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26246\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__26250\,
            I => \N__26243\
        );

    \I__4464\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26238\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__26246\,
            I => \N__26235\
        );

    \I__4462\ : Span4Mux_h
    port map (
            O => \N__26243\,
            I => \N__26232\
        );

    \I__4461\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26229\
        );

    \I__4460\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26226\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__26238\,
            I => \c0.data_in_frame_1_5\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__26235\,
            I => \c0.data_in_frame_1_5\
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__26232\,
            I => \c0.data_in_frame_1_5\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__26229\,
            I => \c0.data_in_frame_1_5\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__26226\,
            I => \c0.data_in_frame_1_5\
        );

    \I__4454\ : CascadeMux
    port map (
            O => \N__26215\,
            I => \c0.n20_adj_2340_cascade_\
        );

    \I__4453\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26209\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__26209\,
            I => \N__26204\
        );

    \I__4451\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26200\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__26207\,
            I => \N__26197\
        );

    \I__4449\ : Span4Mux_h
    port map (
            O => \N__26204\,
            I => \N__26194\
        );

    \I__4448\ : InMux
    port map (
            O => \N__26203\,
            I => \N__26191\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__26200\,
            I => \N__26188\
        );

    \I__4446\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26185\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__26194\,
            I => data_in_3_2
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__26191\,
            I => data_in_3_2
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__26188\,
            I => data_in_3_2
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__26185\,
            I => data_in_3_2
        );

    \I__4441\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26170\
        );

    \I__4440\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26165\
        );

    \I__4439\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26165\
        );

    \I__4438\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26162\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__26170\,
            I => \N__26159\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__26165\,
            I => data_in_2_2
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__26162\,
            I => data_in_2_2
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__26159\,
            I => data_in_2_2
        );

    \I__4433\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26145\
        );

    \I__4432\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26145\
        );

    \I__4431\ : InMux
    port map (
            O => \N__26150\,
            I => \N__26141\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__26145\,
            I => \N__26138\
        );

    \I__4429\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26135\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__26141\,
            I => \N__26132\
        );

    \I__4427\ : Span4Mux_h
    port map (
            O => \N__26138\,
            I => \N__26126\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__26135\,
            I => \N__26126\
        );

    \I__4425\ : Span4Mux_h
    port map (
            O => \N__26132\,
            I => \N__26123\
        );

    \I__4424\ : InMux
    port map (
            O => \N__26131\,
            I => \N__26120\
        );

    \I__4423\ : Sp12to4
    port map (
            O => \N__26126\,
            I => \N__26117\
        );

    \I__4422\ : Odrv4
    port map (
            O => \N__26123\,
            I => data_in_1_2
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__26120\,
            I => data_in_1_2
        );

    \I__4420\ : Odrv12
    port map (
            O => \N__26117\,
            I => data_in_1_2
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__26110\,
            I => \N__26106\
        );

    \I__4418\ : CascadeMux
    port map (
            O => \N__26109\,
            I => \N__26103\
        );

    \I__4417\ : InMux
    port map (
            O => \N__26106\,
            I => \N__26100\
        );

    \I__4416\ : InMux
    port map (
            O => \N__26103\,
            I => \N__26097\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__26100\,
            I => \c0.data_in_frame_10_3\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__26097\,
            I => \c0.data_in_frame_10_3\
        );

    \I__4413\ : InMux
    port map (
            O => \N__26092\,
            I => \N__26088\
        );

    \I__4412\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26085\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__26088\,
            I => \N__26082\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__26085\,
            I => data_in_frame_6_6
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__26082\,
            I => data_in_frame_6_6
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__26077\,
            I => \N__26074\
        );

    \I__4407\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26071\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__26071\,
            I => \N__26067\
        );

    \I__4405\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26064\
        );

    \I__4404\ : Span4Mux_h
    port map (
            O => \N__26067\,
            I => \N__26061\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__26064\,
            I => data_in_frame_7_7
        );

    \I__4402\ : Odrv4
    port map (
            O => \N__26061\,
            I => data_in_frame_7_7
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__26056\,
            I => \c0.n2351_cascade_\
        );

    \I__4400\ : InMux
    port map (
            O => \N__26053\,
            I => \N__26050\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__26050\,
            I => \N__26046\
        );

    \I__4398\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26043\
        );

    \I__4397\ : Span4Mux_v
    port map (
            O => \N__26046\,
            I => \N__26040\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__26043\,
            I => data_in_frame_6_7
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__26040\,
            I => data_in_frame_6_7
        );

    \I__4394\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26031\
        );

    \I__4393\ : InMux
    port map (
            O => \N__26034\,
            I => \N__26028\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__26031\,
            I => data_in_frame_6_1
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__26028\,
            I => data_in_frame_6_1
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__26023\,
            I => \c0.n2352_cascade_\
        );

    \I__4389\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26017\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__26017\,
            I => \N__26013\
        );

    \I__4387\ : InMux
    port map (
            O => \N__26016\,
            I => \N__26010\
        );

    \I__4386\ : Span4Mux_h
    port map (
            O => \N__26013\,
            I => \N__26007\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__26010\,
            I => data_in_frame_6_3
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__26007\,
            I => data_in_frame_6_3
        );

    \I__4383\ : CascadeMux
    port map (
            O => \N__26002\,
            I => \N__25999\
        );

    \I__4382\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25996\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__25996\,
            I => \N__25993\
        );

    \I__4380\ : Span4Mux_v
    port map (
            O => \N__25993\,
            I => \N__25989\
        );

    \I__4379\ : InMux
    port map (
            O => \N__25992\,
            I => \N__25986\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__25989\,
            I => \N__25983\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__25986\,
            I => data_in_frame_6_4
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__25983\,
            I => data_in_frame_6_4
        );

    \I__4375\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25975\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__25975\,
            I => \c0.n23_adj_2145\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__25972\,
            I => \c0.n9541_cascade_\
        );

    \I__4372\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25966\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__25966\,
            I => \N__25963\
        );

    \I__4370\ : Span4Mux_h
    port map (
            O => \N__25963\,
            I => \N__25959\
        );

    \I__4369\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25956\
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__25959\,
            I => \c0.n16943\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__25956\,
            I => \c0.n16943\
        );

    \I__4366\ : InMux
    port map (
            O => \N__25951\,
            I => \N__25945\
        );

    \I__4365\ : InMux
    port map (
            O => \N__25950\,
            I => \N__25942\
        );

    \I__4364\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25937\
        );

    \I__4363\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25937\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__25945\,
            I => data_in_frame_0_2
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__25942\,
            I => data_in_frame_0_2
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__25937\,
            I => data_in_frame_0_2
        );

    \I__4359\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25926\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__25929\,
            I => \N__25922\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__25926\,
            I => \N__25919\
        );

    \I__4356\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25914\
        );

    \I__4355\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25914\
        );

    \I__4354\ : Span4Mux_v
    port map (
            O => \N__25919\,
            I => \N__25909\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__25914\,
            I => \N__25909\
        );

    \I__4352\ : Span4Mux_h
    port map (
            O => \N__25909\,
            I => \N__25905\
        );

    \I__4351\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25902\
        );

    \I__4350\ : Span4Mux_v
    port map (
            O => \N__25905\,
            I => \N__25899\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__25902\,
            I => data_in_3_5
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__25899\,
            I => data_in_3_5
        );

    \I__4347\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25891\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__25891\,
            I => \N__25888\
        );

    \I__4345\ : Span4Mux_v
    port map (
            O => \N__25888\,
            I => \N__25883\
        );

    \I__4344\ : InMux
    port map (
            O => \N__25887\,
            I => \N__25880\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__25886\,
            I => \N__25876\
        );

    \I__4342\ : Span4Mux_h
    port map (
            O => \N__25883\,
            I => \N__25871\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__25880\,
            I => \N__25871\
        );

    \I__4340\ : InMux
    port map (
            O => \N__25879\,
            I => \N__25866\
        );

    \I__4339\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25866\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__25871\,
            I => data_in_2_5
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__25866\,
            I => data_in_2_5
        );

    \I__4336\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25855\
        );

    \I__4335\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25855\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25852\
        );

    \I__4333\ : Span4Mux_v
    port map (
            O => \N__25852\,
            I => \N__25847\
        );

    \I__4332\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25842\
        );

    \I__4331\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25842\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__25847\,
            I => data_in_2_7
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__25842\,
            I => data_in_2_7
        );

    \I__4328\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25834\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__25834\,
            I => \N__25831\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__25831\,
            I => \c0.n8_adj_2157\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__25828\,
            I => \N__25825\
        );

    \I__4324\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25819\
        );

    \I__4323\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25819\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__25819\,
            I => \N__25814\
        );

    \I__4321\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25809\
        );

    \I__4320\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25809\
        );

    \I__4319\ : Span4Mux_h
    port map (
            O => \N__25814\,
            I => \N__25806\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__25809\,
            I => data_in_3_7
        );

    \I__4317\ : Odrv4
    port map (
            O => \N__25806\,
            I => data_in_3_7
        );

    \I__4316\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25798\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__25798\,
            I => \N__25795\
        );

    \I__4314\ : Span4Mux_h
    port map (
            O => \N__25795\,
            I => \N__25791\
        );

    \I__4313\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25787\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__25791\,
            I => \N__25784\
        );

    \I__4311\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25781\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__25787\,
            I => data_in_3_3
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__25784\,
            I => data_in_3_3
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__25781\,
            I => data_in_3_3
        );

    \I__4307\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25771\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__25771\,
            I => \N__25767\
        );

    \I__4305\ : InMux
    port map (
            O => \N__25770\,
            I => \N__25764\
        );

    \I__4304\ : Span4Mux_v
    port map (
            O => \N__25767\,
            I => \N__25761\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__25764\,
            I => data_in_frame_7_0
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__25761\,
            I => data_in_frame_7_0
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__25756\,
            I => \N__25753\
        );

    \I__4300\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25750\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__25750\,
            I => \N__25746\
        );

    \I__4298\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25743\
        );

    \I__4297\ : Span4Mux_h
    port map (
            O => \N__25746\,
            I => \N__25740\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__25743\,
            I => data_in_frame_7_6
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__25740\,
            I => data_in_frame_7_6
        );

    \I__4294\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25732\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__25732\,
            I => \N__25728\
        );

    \I__4292\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25725\
        );

    \I__4291\ : Span4Mux_h
    port map (
            O => \N__25728\,
            I => \N__25719\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__25725\,
            I => \N__25719\
        );

    \I__4289\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25716\
        );

    \I__4288\ : Span4Mux_v
    port map (
            O => \N__25719\,
            I => \N__25706\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__25716\,
            I => \N__25706\
        );

    \I__4286\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25703\
        );

    \I__4285\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25700\
        );

    \I__4284\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25695\
        );

    \I__4283\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25695\
        );

    \I__4282\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25692\
        );

    \I__4281\ : Span4Mux_h
    port map (
            O => \N__25706\,
            I => \N__25689\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__25703\,
            I => \N__25680\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__25700\,
            I => \N__25680\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__25695\,
            I => \N__25680\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__25692\,
            I => \N__25680\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__25689\,
            I => n16896
        );

    \I__4275\ : Odrv12
    port map (
            O => \N__25680\,
            I => n16896
        );

    \I__4274\ : CascadeMux
    port map (
            O => \N__25675\,
            I => \N__25669\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__25674\,
            I => \N__25666\
        );

    \I__4272\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25661\
        );

    \I__4271\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25658\
        );

    \I__4270\ : InMux
    port map (
            O => \N__25669\,
            I => \N__25653\
        );

    \I__4269\ : InMux
    port map (
            O => \N__25666\,
            I => \N__25653\
        );

    \I__4268\ : CascadeMux
    port map (
            O => \N__25665\,
            I => \N__25650\
        );

    \I__4267\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25646\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__25661\,
            I => \N__25643\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__25658\,
            I => \N__25640\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__25653\,
            I => \N__25635\
        );

    \I__4263\ : InMux
    port map (
            O => \N__25650\,
            I => \N__25630\
        );

    \I__4262\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25630\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__25646\,
            I => \N__25627\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__25643\,
            I => \N__25622\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__25640\,
            I => \N__25622\
        );

    \I__4258\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25619\
        );

    \I__4257\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25616\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__25635\,
            I => rx_data_6
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__25630\,
            I => rx_data_6
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__25627\,
            I => rx_data_6
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__25622\,
            I => rx_data_6
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__25619\,
            I => rx_data_6
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__25616\,
            I => rx_data_6
        );

    \I__4250\ : InMux
    port map (
            O => \N__25603\,
            I => \N__25599\
        );

    \I__4249\ : InMux
    port map (
            O => \N__25602\,
            I => \N__25596\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__25599\,
            I => \N__25590\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__25596\,
            I => \N__25586\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__25595\,
            I => \N__25582\
        );

    \I__4245\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25579\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__25593\,
            I => \N__25576\
        );

    \I__4243\ : Sp12to4
    port map (
            O => \N__25590\,
            I => \N__25573\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__25589\,
            I => \N__25570\
        );

    \I__4241\ : Span4Mux_v
    port map (
            O => \N__25586\,
            I => \N__25567\
        );

    \I__4240\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25564\
        );

    \I__4239\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25559\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__25579\,
            I => \N__25556\
        );

    \I__4237\ : InMux
    port map (
            O => \N__25576\,
            I => \N__25553\
        );

    \I__4236\ : Span12Mux_v
    port map (
            O => \N__25573\,
            I => \N__25550\
        );

    \I__4235\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25547\
        );

    \I__4234\ : Span4Mux_s1_h
    port map (
            O => \N__25567\,
            I => \N__25542\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__25564\,
            I => \N__25542\
        );

    \I__4232\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25539\
        );

    \I__4231\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25536\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__25559\,
            I => rx_data_0
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__25556\,
            I => rx_data_0
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__25553\,
            I => rx_data_0
        );

    \I__4227\ : Odrv12
    port map (
            O => \N__25550\,
            I => rx_data_0
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__25547\,
            I => rx_data_0
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__25542\,
            I => rx_data_0
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__25539\,
            I => rx_data_0
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__25536\,
            I => rx_data_0
        );

    \I__4222\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25516\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__25516\,
            I => \N__25510\
        );

    \I__4220\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25503\
        );

    \I__4219\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25503\
        );

    \I__4218\ : InMux
    port map (
            O => \N__25513\,
            I => \N__25503\
        );

    \I__4217\ : Odrv12
    port map (
            O => \N__25510\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__25503\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__4215\ : SRMux
    port map (
            O => \N__25498\,
            I => \N__25495\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25492\
        );

    \I__4213\ : Span4Mux_v
    port map (
            O => \N__25492\,
            I => \N__25489\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__25489\,
            I => \c0.n16365\
        );

    \I__4211\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25483\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__25483\,
            I => \N__25480\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__25480\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_12\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__25477\,
            I => \N__25474\
        );

    \I__4207\ : InMux
    port map (
            O => \N__25474\,
            I => \N__25471\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__25471\,
            I => \N__25466\
        );

    \I__4205\ : InMux
    port map (
            O => \N__25470\,
            I => \N__25463\
        );

    \I__4204\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25460\
        );

    \I__4203\ : Span4Mux_v
    port map (
            O => \N__25466\,
            I => \N__25455\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__25463\,
            I => \N__25455\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__25460\,
            I => \N__25452\
        );

    \I__4200\ : Span4Mux_h
    port map (
            O => \N__25455\,
            I => \N__25446\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__25452\,
            I => \N__25446\
        );

    \I__4198\ : InMux
    port map (
            O => \N__25451\,
            I => \N__25443\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__25446\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__25443\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__4195\ : SRMux
    port map (
            O => \N__25438\,
            I => \N__25435\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__25435\,
            I => \N__25432\
        );

    \I__4193\ : Span4Mux_h
    port map (
            O => \N__25432\,
            I => \N__25429\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__25429\,
            I => \c0.n3_adj_2245\
        );

    \I__4191\ : SRMux
    port map (
            O => \N__25426\,
            I => \N__25423\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__25423\,
            I => \N__25420\
        );

    \I__4189\ : Span4Mux_v
    port map (
            O => \N__25420\,
            I => \N__25417\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__25417\,
            I => \c0.n16351\
        );

    \I__4187\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25409\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__25413\,
            I => \N__25405\
        );

    \I__4185\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25402\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__25409\,
            I => \N__25399\
        );

    \I__4183\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25394\
        );

    \I__4182\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25394\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__25402\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__4180\ : Odrv12
    port map (
            O => \N__25399\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__25394\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__4178\ : SRMux
    port map (
            O => \N__25387\,
            I => \N__25384\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__25384\,
            I => \N__25381\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__25381\,
            I => \N__25378\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__25378\,
            I => \c0.n16367\
        );

    \I__4174\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25370\
        );

    \I__4173\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25367\
        );

    \I__4172\ : InMux
    port map (
            O => \N__25373\,
            I => \N__25363\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__25370\,
            I => \N__25360\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__25367\,
            I => \N__25357\
        );

    \I__4169\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25354\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__25363\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__4167\ : Odrv12
    port map (
            O => \N__25360\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__25357\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__25354\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__4164\ : SRMux
    port map (
            O => \N__25345\,
            I => \N__25342\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25339\
        );

    \I__4162\ : Span4Mux_v
    port map (
            O => \N__25339\,
            I => \N__25336\
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__25336\,
            I => \c0.n16357\
        );

    \I__4160\ : InMux
    port map (
            O => \N__25333\,
            I => \N__25330\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__25330\,
            I => \N__25325\
        );

    \I__4158\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25322\
        );

    \I__4157\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25319\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__25325\,
            I => \N__25314\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25314\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__25319\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__25314\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__4152\ : SRMux
    port map (
            O => \N__25309\,
            I => \N__25306\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__25306\,
            I => \N__25303\
        );

    \I__4150\ : Span4Mux_s3_h
    port map (
            O => \N__25303\,
            I => \N__25300\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__25300\,
            I => \N__25297\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__25297\,
            I => \c0.n16355\
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__25294\,
            I => \N__25289\
        );

    \I__4146\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25286\
        );

    \I__4145\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25283\
        );

    \I__4144\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25280\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25277\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__25283\,
            I => data_in_0_1
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__25280\,
            I => data_in_0_1
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__25277\,
            I => data_in_0_1
        );

    \I__4139\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25267\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__25267\,
            I => \N__25264\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__25264\,
            I => \c0.n17266\
        );

    \I__4136\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25256\
        );

    \I__4135\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25253\
        );

    \I__4134\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25250\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__25256\,
            I => \N__25247\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__25253\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__25250\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__4130\ : Odrv12
    port map (
            O => \N__25247\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__4129\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25237\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__25237\,
            I => \N__25234\
        );

    \I__4127\ : Odrv4
    port map (
            O => \N__25234\,
            I => \c0.n6_adj_2213\
        );

    \I__4126\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25228\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__25228\,
            I => \c0.n16869\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__25225\,
            I => \c0.n16869_cascade_\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__25222\,
            I => \c0.n16871_cascade_\
        );

    \I__4122\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25216\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__25216\,
            I => \c0.n16876\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__25213\,
            I => \N__25210\
        );

    \I__4119\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25207\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__25207\,
            I => \c0.n50\
        );

    \I__4117\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25201\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25198\
        );

    \I__4115\ : Span4Mux_h
    port map (
            O => \N__25198\,
            I => \N__25195\
        );

    \I__4114\ : Span4Mux_v
    port map (
            O => \N__25195\,
            I => \N__25192\
        );

    \I__4113\ : Odrv4
    port map (
            O => \N__25192\,
            I => \c0.n46\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__25189\,
            I => \c0.n56_adj_2146_cascade_\
        );

    \I__4111\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25183\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__25183\,
            I => \c0.n51\
        );

    \I__4109\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25176\
        );

    \I__4108\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25172\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__25176\,
            I => \N__25169\
        );

    \I__4106\ : InMux
    port map (
            O => \N__25175\,
            I => \N__25165\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__25172\,
            I => \N__25160\
        );

    \I__4104\ : Span4Mux_v
    port map (
            O => \N__25169\,
            I => \N__25160\
        );

    \I__4103\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25157\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__25165\,
            I => \N__25154\
        );

    \I__4101\ : Span4Mux_v
    port map (
            O => \N__25160\,
            I => \N__25151\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__25157\,
            I => \c0.n9346\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__25154\,
            I => \c0.n9346\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__25151\,
            I => \c0.n9346\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__25144\,
            I => \N__25141\
        );

    \I__4096\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25137\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__25140\,
            I => \N__25134\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__25137\,
            I => \N__25131\
        );

    \I__4093\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25128\
        );

    \I__4092\ : Span4Mux_v
    port map (
            O => \N__25131\,
            I => \N__25123\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__25128\,
            I => \N__25123\
        );

    \I__4090\ : Span4Mux_h
    port map (
            O => \N__25123\,
            I => \N__25117\
        );

    \I__4089\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25113\
        );

    \I__4088\ : InMux
    port map (
            O => \N__25121\,
            I => \N__25110\
        );

    \I__4087\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25107\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__25117\,
            I => \N__25104\
        );

    \I__4085\ : InMux
    port map (
            O => \N__25116\,
            I => \N__25101\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__25113\,
            I => \N__25096\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__25110\,
            I => \N__25096\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__25107\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__25104\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__25101\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__4079\ : Odrv12
    port map (
            O => \N__25096\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__4078\ : InMux
    port map (
            O => \N__25087\,
            I => \N__25081\
        );

    \I__4077\ : InMux
    port map (
            O => \N__25086\,
            I => \N__25077\
        );

    \I__4076\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25074\
        );

    \I__4075\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25070\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25067\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__25080\,
            I => \N__25063\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__25077\,
            I => \N__25057\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__25074\,
            I => \N__25057\
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__25073\,
            I => \N__25054\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__25070\,
            I => \N__25051\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__25067\,
            I => \N__25048\
        );

    \I__4067\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25045\
        );

    \I__4066\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25040\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25040\
        );

    \I__4064\ : Span4Mux_v
    port map (
            O => \N__25057\,
            I => \N__25037\
        );

    \I__4063\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25034\
        );

    \I__4062\ : Span4Mux_v
    port map (
            O => \N__25051\,
            I => \N__25029\
        );

    \I__4061\ : Span4Mux_h
    port map (
            O => \N__25048\,
            I => \N__25029\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__25045\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__25040\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__25037\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__25034\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__25029\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__4055\ : CascadeMux
    port map (
            O => \N__25018\,
            I => \N__25013\
        );

    \I__4054\ : InMux
    port map (
            O => \N__25017\,
            I => \N__25010\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__25016\,
            I => \N__25007\
        );

    \I__4052\ : InMux
    port map (
            O => \N__25013\,
            I => \N__25004\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__25010\,
            I => \N__25001\
        );

    \I__4050\ : InMux
    port map (
            O => \N__25007\,
            I => \N__24998\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__25004\,
            I => \N__24994\
        );

    \I__4048\ : Span4Mux_v
    port map (
            O => \N__25001\,
            I => \N__24989\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__24998\,
            I => \N__24989\
        );

    \I__4046\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24986\
        );

    \I__4045\ : Span4Mux_v
    port map (
            O => \N__24994\,
            I => \N__24983\
        );

    \I__4044\ : Span4Mux_h
    port map (
            O => \N__24989\,
            I => \N__24980\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__24986\,
            I => \N__24975\
        );

    \I__4042\ : Span4Mux_v
    port map (
            O => \N__24983\,
            I => \N__24975\
        );

    \I__4041\ : Span4Mux_v
    port map (
            O => \N__24980\,
            I => \N__24972\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__24975\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__24972\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__4038\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__24964\,
            I => \c0.n45\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__24961\,
            I => \N__24957\
        );

    \I__4035\ : InMux
    port map (
            O => \N__24960\,
            I => \N__24952\
        );

    \I__4034\ : InMux
    port map (
            O => \N__24957\,
            I => \N__24949\
        );

    \I__4033\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24946\
        );

    \I__4032\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24943\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__24952\,
            I => \N__24940\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__24949\,
            I => \N__24937\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24934\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__24943\,
            I => \N__24931\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__24940\,
            I => \N__24924\
        );

    \I__4026\ : Span4Mux_v
    port map (
            O => \N__24937\,
            I => \N__24924\
        );

    \I__4025\ : Span4Mux_h
    port map (
            O => \N__24934\,
            I => \N__24924\
        );

    \I__4024\ : Span4Mux_v
    port map (
            O => \N__24931\,
            I => \N__24921\
        );

    \I__4023\ : Span4Mux_h
    port map (
            O => \N__24924\,
            I => \N__24918\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__24921\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__24918\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__24913\,
            I => \N__24910\
        );

    \I__4019\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24904\
        );

    \I__4018\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24901\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__24908\,
            I => \N__24898\
        );

    \I__4016\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24895\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__24904\,
            I => \N__24892\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__24901\,
            I => \N__24889\
        );

    \I__4013\ : InMux
    port map (
            O => \N__24898\,
            I => \N__24886\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__24895\,
            I => \N__24883\
        );

    \I__4011\ : Span4Mux_v
    port map (
            O => \N__24892\,
            I => \N__24880\
        );

    \I__4010\ : Span4Mux_v
    port map (
            O => \N__24889\,
            I => \N__24877\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__24886\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__4008\ : Odrv12
    port map (
            O => \N__24883\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__24880\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__24877\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__24868\,
            I => \N__24865\
        );

    \I__4004\ : InMux
    port map (
            O => \N__24865\,
            I => \N__24861\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__24864\,
            I => \N__24857\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__24861\,
            I => \N__24854\
        );

    \I__4001\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24851\
        );

    \I__4000\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24848\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__24854\,
            I => \N__24840\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__24851\,
            I => \N__24840\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__24848\,
            I => \N__24840\
        );

    \I__3996\ : InMux
    port map (
            O => \N__24847\,
            I => \N__24837\
        );

    \I__3995\ : Span4Mux_h
    port map (
            O => \N__24840\,
            I => \N__24834\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__24837\,
            I => \N__24831\
        );

    \I__3993\ : Span4Mux_h
    port map (
            O => \N__24834\,
            I => \N__24828\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__24831\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__24828\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__24823\,
            I => \N__24819\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__24822\,
            I => \N__24815\
        );

    \I__3988\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24812\
        );

    \I__3987\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24809\
        );

    \I__3986\ : InMux
    port map (
            O => \N__24815\,
            I => \N__24805\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__24812\,
            I => \N__24800\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24800\
        );

    \I__3983\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24797\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__24805\,
            I => \N__24794\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__24800\,
            I => \N__24789\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__24797\,
            I => \N__24789\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__24794\,
            I => \N__24784\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__24789\,
            I => \N__24784\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__24784\,
            I => \N__24781\
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__24781\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__3975\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24775\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__24775\,
            I => \c0.n47_adj_2144\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__24772\,
            I => \N__24769\
        );

    \I__3972\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24765\
        );

    \I__3971\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24762\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__24765\,
            I => \N__24758\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24755\
        );

    \I__3968\ : InMux
    port map (
            O => \N__24761\,
            I => \N__24752\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__24758\,
            I => \N__24748\
        );

    \I__3966\ : Span4Mux_h
    port map (
            O => \N__24755\,
            I => \N__24743\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__24752\,
            I => \N__24743\
        );

    \I__3964\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24740\
        );

    \I__3963\ : Span4Mux_h
    port map (
            O => \N__24748\,
            I => \N__24735\
        );

    \I__3962\ : Span4Mux_h
    port map (
            O => \N__24743\,
            I => \N__24735\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__24740\,
            I => \N__24732\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__24735\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__3959\ : Odrv12
    port map (
            O => \N__24732\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__24727\,
            I => \N__24723\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__24726\,
            I => \N__24719\
        );

    \I__3956\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24716\
        );

    \I__3955\ : InMux
    port map (
            O => \N__24722\,
            I => \N__24713\
        );

    \I__3954\ : InMux
    port map (
            O => \N__24719\,
            I => \N__24709\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__24716\,
            I => \N__24704\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__24713\,
            I => \N__24704\
        );

    \I__3951\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24701\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__24709\,
            I => \N__24698\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__24704\,
            I => \N__24693\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__24701\,
            I => \N__24693\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__24698\,
            I => \N__24688\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__24693\,
            I => \N__24688\
        );

    \I__3945\ : Span4Mux_h
    port map (
            O => \N__24688\,
            I => \N__24685\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__24685\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__3943\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24677\
        );

    \I__3942\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24674\
        );

    \I__3941\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24671\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__24677\,
            I => \N__24668\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__24674\,
            I => \N__24664\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24661\
        );

    \I__3937\ : Span4Mux_h
    port map (
            O => \N__24668\,
            I => \N__24658\
        );

    \I__3936\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24655\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__24664\,
            I => \N__24652\
        );

    \I__3934\ : Odrv4
    port map (
            O => \N__24661\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__3933\ : Odrv4
    port map (
            O => \N__24658\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__24655\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__3931\ : Odrv4
    port map (
            O => \N__24652\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__3930\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24640\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__24640\,
            I => \c0.n49\
        );

    \I__3928\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24634\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__24634\,
            I => \N__24631\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__24631\,
            I => \c0.n59\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__24628\,
            I => \c0.n61_cascade_\
        );

    \I__3924\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24622\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__24622\,
            I => \c0.n10_adj_2336\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__24619\,
            I => \c0.n16133_cascade_\
        );

    \I__3921\ : InMux
    port map (
            O => \N__24616\,
            I => \N__24612\
        );

    \I__3920\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24609\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__24612\,
            I => \c0.n16898\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__24609\,
            I => \c0.n16898\
        );

    \I__3917\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24596\
        );

    \I__3916\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24596\
        );

    \I__3915\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24593\
        );

    \I__3914\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24590\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__24596\,
            I => \N__24587\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__24593\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__24590\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__3910\ : Odrv12
    port map (
            O => \N__24587\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__3909\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24577\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__24577\,
            I => \c0.n52\
        );

    \I__3907\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24571\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__24571\,
            I => \N__24568\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__24568\,
            I => \N__24565\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__24565\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_4\
        );

    \I__3903\ : SRMux
    port map (
            O => \N__24562\,
            I => \N__24559\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__24559\,
            I => \N__24556\
        );

    \I__3901\ : Span4Mux_h
    port map (
            O => \N__24556\,
            I => \N__24553\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__24553\,
            I => \c0.n3_adj_2257\
        );

    \I__3899\ : CascadeMux
    port map (
            O => \N__24550\,
            I => \N__24547\
        );

    \I__3898\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24542\
        );

    \I__3897\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24539\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__24545\,
            I => \N__24536\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__24542\,
            I => \N__24530\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__24539\,
            I => \N__24530\
        );

    \I__3893\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24527\
        );

    \I__3892\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24524\
        );

    \I__3891\ : Span4Mux_v
    port map (
            O => \N__24530\,
            I => \N__24521\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__24527\,
            I => \N__24516\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__24524\,
            I => \N__24516\
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__24521\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__3887\ : Odrv12
    port map (
            O => \N__24516\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__24511\,
            I => \N__24506\
        );

    \I__3885\ : InMux
    port map (
            O => \N__24510\,
            I => \N__24503\
        );

    \I__3884\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24500\
        );

    \I__3883\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24497\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__24503\,
            I => \N__24492\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__24500\,
            I => \N__24492\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__24497\,
            I => \N__24487\
        );

    \I__3879\ : Span4Mux_h
    port map (
            O => \N__24492\,
            I => \N__24484\
        );

    \I__3878\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24479\
        );

    \I__3877\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24479\
        );

    \I__3876\ : Span4Mux_h
    port map (
            O => \N__24487\,
            I => \N__24476\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__24484\,
            I => \N__24472\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24469\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__24476\,
            I => \N__24466\
        );

    \I__3872\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24463\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__24472\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__3870\ : Odrv12
    port map (
            O => \N__24469\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__24466\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__24463\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__3867\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24450\
        );

    \I__3866\ : InMux
    port map (
            O => \N__24453\,
            I => \N__24447\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__24450\,
            I => \N__24441\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__24447\,
            I => \N__24441\
        );

    \I__3863\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24437\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__24441\,
            I => \N__24434\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__24440\,
            I => \N__24430\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__24437\,
            I => \N__24426\
        );

    \I__3859\ : Sp12to4
    port map (
            O => \N__24434\,
            I => \N__24423\
        );

    \I__3858\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24420\
        );

    \I__3857\ : InMux
    port map (
            O => \N__24430\,
            I => \N__24415\
        );

    \I__3856\ : InMux
    port map (
            O => \N__24429\,
            I => \N__24415\
        );

    \I__3855\ : Span4Mux_h
    port map (
            O => \N__24426\,
            I => \N__24412\
        );

    \I__3854\ : Odrv12
    port map (
            O => \N__24423\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__24420\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__24415\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__24412\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__3850\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24399\
        );

    \I__3849\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24395\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__24399\,
            I => \N__24392\
        );

    \I__3847\ : InMux
    port map (
            O => \N__24398\,
            I => \N__24389\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__24395\,
            I => \N__24385\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__24392\,
            I => \N__24382\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__24389\,
            I => \N__24379\
        );

    \I__3843\ : CascadeMux
    port map (
            O => \N__24388\,
            I => \N__24376\
        );

    \I__3842\ : Span4Mux_v
    port map (
            O => \N__24385\,
            I => \N__24373\
        );

    \I__3841\ : Span4Mux_s3_h
    port map (
            O => \N__24382\,
            I => \N__24368\
        );

    \I__3840\ : Span4Mux_h
    port map (
            O => \N__24379\,
            I => \N__24368\
        );

    \I__3839\ : InMux
    port map (
            O => \N__24376\,
            I => \N__24365\
        );

    \I__3838\ : Span4Mux_v
    port map (
            O => \N__24373\,
            I => \N__24362\
        );

    \I__3837\ : Span4Mux_v
    port map (
            O => \N__24368\,
            I => \N__24359\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__24365\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__24362\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__24359\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__24352\,
            I => \c0.n30_cascade_\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__24349\,
            I => \N__24344\
        );

    \I__3831\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24341\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__24347\,
            I => \N__24338\
        );

    \I__3829\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24334\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__24341\,
            I => \N__24331\
        );

    \I__3827\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24326\
        );

    \I__3826\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24326\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__24334\,
            I => \N__24323\
        );

    \I__3824\ : Span4Mux_v
    port map (
            O => \N__24331\,
            I => \N__24320\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__24326\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__3822\ : Odrv4
    port map (
            O => \N__24323\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__24320\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__3820\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24309\
        );

    \I__3819\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24306\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__24309\,
            I => \c0.n56\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__24306\,
            I => \c0.n56\
        );

    \I__3816\ : InMux
    port map (
            O => \N__24301\,
            I => \N__24297\
        );

    \I__3815\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24294\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__24297\,
            I => \N__24291\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__24294\,
            I => \c0.n446\
        );

    \I__3812\ : Odrv12
    port map (
            O => \N__24291\,
            I => \c0.n446\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__24286\,
            I => \c0.n446_cascade_\
        );

    \I__3810\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24277\
        );

    \I__3809\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24277\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__24277\,
            I => \c0.n456\
        );

    \I__3807\ : SRMux
    port map (
            O => \N__24274\,
            I => \N__24271\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__24271\,
            I => \N__24268\
        );

    \I__3805\ : Span4Mux_h
    port map (
            O => \N__24268\,
            I => \N__24265\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__24265\,
            I => \c0.n16371\
        );

    \I__3803\ : SRMux
    port map (
            O => \N__24262\,
            I => \N__24259\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__24259\,
            I => \N__24256\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__24256\,
            I => \c0.n16453\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__24253\,
            I => \c0.n8938_cascade_\
        );

    \I__3799\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24247\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__24247\,
            I => \N__24244\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__24244\,
            I => \c0.n22_adj_2164\
        );

    \I__3796\ : CascadeMux
    port map (
            O => \N__24241\,
            I => \c0.n22_adj_2164_cascade_\
        );

    \I__3795\ : InMux
    port map (
            O => \N__24238\,
            I => \N__24232\
        );

    \I__3794\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24232\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__24232\,
            I => \c0.tx_transmit_N_1949_1\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__24229\,
            I => \c0.n15868_cascade_\
        );

    \I__3791\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24223\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__24223\,
            I => \c0.n8631\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__24220\,
            I => \n10141_cascade_\
        );

    \I__3788\ : InMux
    port map (
            O => \N__24217\,
            I => \c0.n15653\
        );

    \I__3787\ : InMux
    port map (
            O => \N__24214\,
            I => \c0.n15654\
        );

    \I__3786\ : InMux
    port map (
            O => \N__24211\,
            I => \c0.n15655\
        );

    \I__3785\ : InMux
    port map (
            O => \N__24208\,
            I => \c0.n15656\
        );

    \I__3784\ : InMux
    port map (
            O => \N__24205\,
            I => \c0.n15657\
        );

    \I__3783\ : InMux
    port map (
            O => \N__24202\,
            I => \c0.n15658\
        );

    \I__3782\ : InMux
    port map (
            O => \N__24199\,
            I => \c0.n15659\
        );

    \I__3781\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24193\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__24193\,
            I => \c0.n25_adj_2324\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__24190\,
            I => \n4_adj_2458_cascade_\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__24187\,
            I => \N__24184\
        );

    \I__3777\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24179\
        );

    \I__3776\ : InMux
    port map (
            O => \N__24183\,
            I => \N__24174\
        );

    \I__3775\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24174\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__24179\,
            I => \N__24166\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__24174\,
            I => \N__24163\
        );

    \I__3772\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24160\
        );

    \I__3771\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24157\
        );

    \I__3770\ : CascadeMux
    port map (
            O => \N__24171\,
            I => \N__24153\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__24170\,
            I => \N__24150\
        );

    \I__3768\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24147\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__24166\,
            I => \N__24144\
        );

    \I__3766\ : Span4Mux_h
    port map (
            O => \N__24163\,
            I => \N__24139\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__24160\,
            I => \N__24139\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__24157\,
            I => \N__24136\
        );

    \I__3763\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24131\
        );

    \I__3762\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24131\
        );

    \I__3761\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24128\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__24147\,
            I => \r_SM_Main_0\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__24144\,
            I => \r_SM_Main_0\
        );

    \I__3758\ : Odrv4
    port map (
            O => \N__24139\,
            I => \r_SM_Main_0\
        );

    \I__3757\ : Odrv12
    port map (
            O => \N__24136\,
            I => \r_SM_Main_0\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__24131\,
            I => \r_SM_Main_0\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__24128\,
            I => \r_SM_Main_0\
        );

    \I__3754\ : InMux
    port map (
            O => \N__24115\,
            I => \N__24110\
        );

    \I__3753\ : InMux
    port map (
            O => \N__24114\,
            I => \N__24105\
        );

    \I__3752\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24105\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24100\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24097\
        );

    \I__3749\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24094\
        );

    \I__3748\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24091\
        );

    \I__3747\ : Span4Mux_s1_v
    port map (
            O => \N__24100\,
            I => \N__24088\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__24097\,
            I => \N__24083\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__24094\,
            I => \N__24083\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__24091\,
            I => n14060
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__24088\,
            I => n14060
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__24083\,
            I => n14060
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__24076\,
            I => \N__24071\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__24075\,
            I => \N__24068\
        );

    \I__3739\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24056\
        );

    \I__3738\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24056\
        );

    \I__3737\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24056\
        );

    \I__3736\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24053\
        );

    \I__3735\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24050\
        );

    \I__3734\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24046\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__24064\,
            I => \N__24040\
        );

    \I__3732\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24035\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__24056\,
            I => \N__24030\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__24053\,
            I => \N__24030\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__24050\,
            I => \N__24027\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__24049\,
            I => \N__24024\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__24046\,
            I => \N__24020\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24015\
        );

    \I__3725\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24015\
        );

    \I__3724\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24012\
        );

    \I__3723\ : InMux
    port map (
            O => \N__24040\,
            I => \N__24007\
        );

    \I__3722\ : InMux
    port map (
            O => \N__24039\,
            I => \N__24007\
        );

    \I__3721\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24004\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__24035\,
            I => \N__24001\
        );

    \I__3719\ : Span4Mux_v
    port map (
            O => \N__24030\,
            I => \N__23996\
        );

    \I__3718\ : Span4Mux_v
    port map (
            O => \N__24027\,
            I => \N__23996\
        );

    \I__3717\ : InMux
    port map (
            O => \N__24024\,
            I => \N__23991\
        );

    \I__3716\ : InMux
    port map (
            O => \N__24023\,
            I => \N__23991\
        );

    \I__3715\ : Span4Mux_s3_h
    port map (
            O => \N__24020\,
            I => \N__23982\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__24015\,
            I => \N__23982\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__24012\,
            I => \N__23982\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__24007\,
            I => \N__23982\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__24004\,
            I => \r_SM_Main_1\
        );

    \I__3710\ : Odrv12
    port map (
            O => \N__24001\,
            I => \r_SM_Main_1\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__23996\,
            I => \r_SM_Main_1\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__23991\,
            I => \r_SM_Main_1\
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__23982\,
            I => \r_SM_Main_1\
        );

    \I__3706\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23965\
        );

    \I__3705\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23950\
        );

    \I__3704\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23945\
        );

    \I__3703\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23945\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__23965\,
            I => \N__23942\
        );

    \I__3701\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23937\
        );

    \I__3700\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23937\
        );

    \I__3699\ : InMux
    port map (
            O => \N__23962\,
            I => \N__23934\
        );

    \I__3698\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23930\
        );

    \I__3697\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23925\
        );

    \I__3696\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23925\
        );

    \I__3695\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23922\
        );

    \I__3694\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23919\
        );

    \I__3693\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23914\
        );

    \I__3692\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23914\
        );

    \I__3691\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23909\
        );

    \I__3690\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23909\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__23950\,
            I => \N__23906\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__23945\,
            I => \N__23903\
        );

    \I__3687\ : Span4Mux_v
    port map (
            O => \N__23942\,
            I => \N__23896\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__23937\,
            I => \N__23896\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__23934\,
            I => \N__23896\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__23933\,
            I => \N__23893\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__23930\,
            I => \N__23879\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__23925\,
            I => \N__23879\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__23922\,
            I => \N__23879\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__23919\,
            I => \N__23879\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__23914\,
            I => \N__23879\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23879\
        );

    \I__3677\ : Span4Mux_v
    port map (
            O => \N__23906\,
            I => \N__23872\
        );

    \I__3676\ : Span4Mux_s1_h
    port map (
            O => \N__23903\,
            I => \N__23872\
        );

    \I__3675\ : Span4Mux_s3_v
    port map (
            O => \N__23896\,
            I => \N__23869\
        );

    \I__3674\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23864\
        );

    \I__3673\ : InMux
    port map (
            O => \N__23892\,
            I => \N__23864\
        );

    \I__3672\ : Span4Mux_s3_v
    port map (
            O => \N__23879\,
            I => \N__23861\
        );

    \I__3671\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23858\
        );

    \I__3670\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23855\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__23872\,
            I => \N__23852\
        );

    \I__3668\ : Span4Mux_s3_h
    port map (
            O => \N__23869\,
            I => \N__23849\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__23864\,
            I => \N__23844\
        );

    \I__3666\ : Span4Mux_s2_h
    port map (
            O => \N__23861\,
            I => \N__23844\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__23858\,
            I => \r_SM_Main_2\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__23855\,
            I => \r_SM_Main_2\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__23852\,
            I => \r_SM_Main_2\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__23849\,
            I => \r_SM_Main_2\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__23844\,
            I => \r_SM_Main_2\
        );

    \I__3660\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23830\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23827\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__23827\,
            I => n17395
        );

    \I__3657\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23821\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__23821\,
            I => \c0.tx_active_prev\
        );

    \I__3655\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23815\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__23815\,
            I => \c0.n65\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__23812\,
            I => \N__23808\
        );

    \I__3652\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23805\
        );

    \I__3651\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23802\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__23805\,
            I => \c0.data_in_frame_2_7\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__23802\,
            I => \c0.data_in_frame_2_7\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__23797\,
            I => \N__23793\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__23796\,
            I => \N__23790\
        );

    \I__3646\ : InMux
    port map (
            O => \N__23793\,
            I => \N__23785\
        );

    \I__3645\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23785\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__23785\,
            I => \c0.data_in_frame_10_1\
        );

    \I__3643\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23775\
        );

    \I__3642\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23775\
        );

    \I__3641\ : InMux
    port map (
            O => \N__23780\,
            I => \N__23772\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__23775\,
            I => \c0.n9743\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__23772\,
            I => \c0.n9743\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__23767\,
            I => \c0.n16954_cascade_\
        );

    \I__3637\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23758\
        );

    \I__3636\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23758\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__23758\,
            I => \c0.data_in_frame_10_6\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__23755\,
            I => \c0.n18_adj_2174_cascade_\
        );

    \I__3633\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23749\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__23749\,
            I => \c0.n17015\
        );

    \I__3631\ : InMux
    port map (
            O => \N__23746\,
            I => \N__23742\
        );

    \I__3630\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23739\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__23742\,
            I => \c0.data_in_frame_9_4\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__23739\,
            I => \c0.data_in_frame_9_4\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__23734\,
            I => \N__23731\
        );

    \I__3626\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23728\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__23728\,
            I => \N__23725\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__23725\,
            I => \c0.n6_adj_2152\
        );

    \I__3623\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23718\
        );

    \I__3622\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23715\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__23718\,
            I => \N__23709\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23709\
        );

    \I__3619\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23706\
        );

    \I__3618\ : Span4Mux_v
    port map (
            O => \N__23709\,
            I => \N__23703\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__23706\,
            I => \N__23700\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__23703\,
            I => \c0.n13272\
        );

    \I__3615\ : Odrv12
    port map (
            O => \N__23700\,
            I => \c0.n13272\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__23695\,
            I => \c0.n16882_cascade_\
        );

    \I__3613\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23688\
        );

    \I__3612\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23685\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__23688\,
            I => \c0.data_in_frame_10_4\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__23685\,
            I => \c0.data_in_frame_10_4\
        );

    \I__3609\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23676\
        );

    \I__3608\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23673\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__23676\,
            I => \c0.data_in_frame_9_6\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__23673\,
            I => \c0.data_in_frame_9_6\
        );

    \I__3605\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23665\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__23665\,
            I => \N__23661\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__23664\,
            I => \N__23658\
        );

    \I__3602\ : Span4Mux_h
    port map (
            O => \N__23661\,
            I => \N__23655\
        );

    \I__3601\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23652\
        );

    \I__3600\ : Span4Mux_h
    port map (
            O => \N__23655\,
            I => \N__23649\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__23652\,
            I => \c0.data_in_frame_10_0\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__23649\,
            I => \c0.data_in_frame_10_0\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__23644\,
            I => \c0.n17013_cascade_\
        );

    \I__3596\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23638\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23635\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__23635\,
            I => \c0.n17013\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__23632\,
            I => \N__23629\
        );

    \I__3592\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__23626\,
            I => \N__23622\
        );

    \I__3590\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23619\
        );

    \I__3589\ : Span4Mux_h
    port map (
            O => \N__23622\,
            I => \N__23616\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__23619\,
            I => \c0.data_in_frame_9_7\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__23616\,
            I => \c0.data_in_frame_9_7\
        );

    \I__3586\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23608\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__23608\,
            I => \N__23601\
        );

    \I__3584\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23596\
        );

    \I__3583\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23596\
        );

    \I__3582\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23591\
        );

    \I__3581\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23591\
        );

    \I__3580\ : Span4Mux_h
    port map (
            O => \N__23601\,
            I => \N__23588\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__23596\,
            I => data_in_3_6
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__23591\,
            I => data_in_3_6
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__23588\,
            I => data_in_3_6
        );

    \I__3576\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23577\
        );

    \I__3575\ : InMux
    port map (
            O => \N__23580\,
            I => \N__23574\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__23577\,
            I => \N__23569\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__23574\,
            I => \N__23566\
        );

    \I__3572\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23561\
        );

    \I__3571\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23561\
        );

    \I__3570\ : Span4Mux_h
    port map (
            O => \N__23569\,
            I => \N__23558\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__23566\,
            I => \N__23555\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__23561\,
            I => data_in_2_0
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__23558\,
            I => data_in_2_0
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__23555\,
            I => data_in_2_0
        );

    \I__3565\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23545\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__23545\,
            I => \N__23542\
        );

    \I__3563\ : Odrv12
    port map (
            O => \N__23542\,
            I => \c0.n17268\
        );

    \I__3562\ : InMux
    port map (
            O => \N__23539\,
            I => \N__23536\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__23536\,
            I => \N__23532\
        );

    \I__3560\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23527\
        );

    \I__3559\ : Span4Mux_h
    port map (
            O => \N__23532\,
            I => \N__23524\
        );

    \I__3558\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23519\
        );

    \I__3557\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23519\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__23527\,
            I => data_in_1_7
        );

    \I__3555\ : Odrv4
    port map (
            O => \N__23524\,
            I => data_in_1_7
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__23519\,
            I => data_in_1_7
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__23512\,
            I => \N__23508\
        );

    \I__3552\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23504\
        );

    \I__3551\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23499\
        );

    \I__3550\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23499\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__23504\,
            I => data_in_0_3
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__23499\,
            I => data_in_0_3
        );

    \I__3547\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23491\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23488\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__23488\,
            I => \c0.n19_adj_2199\
        );

    \I__3544\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23480\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__23484\,
            I => \N__23476\
        );

    \I__3542\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23473\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__23480\,
            I => \N__23470\
        );

    \I__3540\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23467\
        );

    \I__3539\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23464\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__23473\,
            I => \N__23461\
        );

    \I__3537\ : Span4Mux_v
    port map (
            O => \N__23470\,
            I => \N__23458\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__23467\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__23464\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__23461\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__23458\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__3532\ : SRMux
    port map (
            O => \N__23449\,
            I => \N__23446\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__23446\,
            I => \N__23443\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__23443\,
            I => \c0.n3_adj_2239\
        );

    \I__3529\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23437\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__23437\,
            I => \N__23434\
        );

    \I__3527\ : Odrv12
    port map (
            O => \N__23434\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_17\
        );

    \I__3526\ : InMux
    port map (
            O => \N__23431\,
            I => \N__23423\
        );

    \I__3525\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23410\
        );

    \I__3524\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23410\
        );

    \I__3523\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23403\
        );

    \I__3522\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23403\
        );

    \I__3521\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23403\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__23423\,
            I => \N__23399\
        );

    \I__3519\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23394\
        );

    \I__3518\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23394\
        );

    \I__3517\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23391\
        );

    \I__3516\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23388\
        );

    \I__3515\ : InMux
    port map (
            O => \N__23418\,
            I => \N__23379\
        );

    \I__3514\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23379\
        );

    \I__3513\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23379\
        );

    \I__3512\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23379\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__23410\,
            I => \N__23359\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23359\
        );

    \I__3509\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23348\
        );

    \I__3508\ : Span4Mux_v
    port map (
            O => \N__23399\,
            I => \N__23339\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23339\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__23391\,
            I => \N__23339\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__23388\,
            I => \N__23339\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__23379\,
            I => \N__23336\
        );

    \I__3503\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23327\
        );

    \I__3502\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23327\
        );

    \I__3501\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23327\
        );

    \I__3500\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23327\
        );

    \I__3499\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23312\
        );

    \I__3498\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23312\
        );

    \I__3497\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23312\
        );

    \I__3496\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23312\
        );

    \I__3495\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23312\
        );

    \I__3494\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23312\
        );

    \I__3493\ : InMux
    port map (
            O => \N__23368\,
            I => \N__23312\
        );

    \I__3492\ : InMux
    port map (
            O => \N__23367\,
            I => \N__23303\
        );

    \I__3491\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23303\
        );

    \I__3490\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23303\
        );

    \I__3489\ : InMux
    port map (
            O => \N__23364\,
            I => \N__23303\
        );

    \I__3488\ : Span4Mux_v
    port map (
            O => \N__23359\,
            I => \N__23300\
        );

    \I__3487\ : InMux
    port map (
            O => \N__23358\,
            I => \N__23291\
        );

    \I__3486\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23291\
        );

    \I__3485\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23291\
        );

    \I__3484\ : InMux
    port map (
            O => \N__23355\,
            I => \N__23291\
        );

    \I__3483\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23282\
        );

    \I__3482\ : InMux
    port map (
            O => \N__23353\,
            I => \N__23282\
        );

    \I__3481\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23282\
        );

    \I__3480\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23282\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__23348\,
            I => \N__23277\
        );

    \I__3478\ : Span4Mux_v
    port map (
            O => \N__23339\,
            I => \N__23277\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__23336\,
            I => \c0.n127_adj_2136\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__23327\,
            I => \c0.n127_adj_2136\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__23312\,
            I => \c0.n127_adj_2136\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__23303\,
            I => \c0.n127_adj_2136\
        );

    \I__3473\ : Odrv4
    port map (
            O => \N__23300\,
            I => \c0.n127_adj_2136\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__23291\,
            I => \c0.n127_adj_2136\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__23282\,
            I => \c0.n127_adj_2136\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__23277\,
            I => \c0.n127_adj_2136\
        );

    \I__3469\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23246\
        );

    \I__3468\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23246\
        );

    \I__3467\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23246\
        );

    \I__3466\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23241\
        );

    \I__3465\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23241\
        );

    \I__3464\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23226\
        );

    \I__3463\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23226\
        );

    \I__3462\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23226\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__23246\,
            I => \N__23218\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__23241\,
            I => \N__23218\
        );

    \I__3459\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23215\
        );

    \I__3458\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23206\
        );

    \I__3457\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23206\
        );

    \I__3456\ : InMux
    port map (
            O => \N__23237\,
            I => \N__23206\
        );

    \I__3455\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23206\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__23235\,
            I => \N__23192\
        );

    \I__3453\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23177\
        );

    \I__3452\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23177\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__23226\,
            I => \N__23174\
        );

    \I__3450\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23171\
        );

    \I__3449\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23166\
        );

    \I__3448\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23166\
        );

    \I__3447\ : Span4Mux_h
    port map (
            O => \N__23218\,
            I => \N__23163\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__23215\,
            I => \N__23160\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__23206\,
            I => \N__23157\
        );

    \I__3444\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23148\
        );

    \I__3443\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23148\
        );

    \I__3442\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23148\
        );

    \I__3441\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23148\
        );

    \I__3440\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23133\
        );

    \I__3439\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23133\
        );

    \I__3438\ : InMux
    port map (
            O => \N__23199\,
            I => \N__23133\
        );

    \I__3437\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23133\
        );

    \I__3436\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23133\
        );

    \I__3435\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23133\
        );

    \I__3434\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23133\
        );

    \I__3433\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23124\
        );

    \I__3432\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23124\
        );

    \I__3431\ : InMux
    port map (
            O => \N__23190\,
            I => \N__23124\
        );

    \I__3430\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23124\
        );

    \I__3429\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23113\
        );

    \I__3428\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23113\
        );

    \I__3427\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23113\
        );

    \I__3426\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23113\
        );

    \I__3425\ : InMux
    port map (
            O => \N__23184\,
            I => \N__23113\
        );

    \I__3424\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23108\
        );

    \I__3423\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23108\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__23177\,
            I => \N__23103\
        );

    \I__3421\ : Span4Mux_h
    port map (
            O => \N__23174\,
            I => \N__23103\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__23171\,
            I => \N__23098\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__23166\,
            I => \N__23098\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__23163\,
            I => n127
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__23160\,
            I => n127
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__23157\,
            I => n127
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__23148\,
            I => n127
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__23133\,
            I => n127
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__23124\,
            I => n127
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__23113\,
            I => n127
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__23108\,
            I => n127
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__23103\,
            I => n127
        );

    \I__3409\ : Odrv12
    port map (
            O => \N__23098\,
            I => n127
        );

    \I__3408\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__3406\ : Span4Mux_h
    port map (
            O => \N__23071\,
            I => \N__23068\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__23068\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_16\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__23065\,
            I => \N__23053\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__23064\,
            I => \N__23050\
        );

    \I__3402\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23022\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23022\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23022\
        );

    \I__3399\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23022\
        );

    \I__3398\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23022\
        );

    \I__3397\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23022\
        );

    \I__3396\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23017\
        );

    \I__3395\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23017\
        );

    \I__3394\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23009\
        );

    \I__3393\ : InMux
    port map (
            O => \N__23050\,
            I => \N__23009\
        );

    \I__3392\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23009\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__23048\,
            I => \N__23003\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__23047\,
            I => \N__23000\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__23046\,
            I => \N__22997\
        );

    \I__3388\ : InMux
    port map (
            O => \N__23045\,
            I => \N__22983\
        );

    \I__3387\ : InMux
    port map (
            O => \N__23044\,
            I => \N__22983\
        );

    \I__3386\ : InMux
    port map (
            O => \N__23043\,
            I => \N__22980\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__23042\,
            I => \N__22972\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23041\,
            I => \N__22966\
        );

    \I__3383\ : InMux
    port map (
            O => \N__23040\,
            I => \N__22966\
        );

    \I__3382\ : InMux
    port map (
            O => \N__23039\,
            I => \N__22955\
        );

    \I__3381\ : InMux
    port map (
            O => \N__23038\,
            I => \N__22955\
        );

    \I__3380\ : InMux
    port map (
            O => \N__23037\,
            I => \N__22955\
        );

    \I__3379\ : InMux
    port map (
            O => \N__23036\,
            I => \N__22955\
        );

    \I__3378\ : InMux
    port map (
            O => \N__23035\,
            I => \N__22955\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__23022\,
            I => \N__22949\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__22949\
        );

    \I__3375\ : InMux
    port map (
            O => \N__23016\,
            I => \N__22946\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__22943\
        );

    \I__3373\ : InMux
    port map (
            O => \N__23008\,
            I => \N__22928\
        );

    \I__3372\ : InMux
    port map (
            O => \N__23007\,
            I => \N__22928\
        );

    \I__3371\ : InMux
    port map (
            O => \N__23006\,
            I => \N__22928\
        );

    \I__3370\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22928\
        );

    \I__3369\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22928\
        );

    \I__3368\ : InMux
    port map (
            O => \N__22997\,
            I => \N__22928\
        );

    \I__3367\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22928\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__22995\,
            I => \N__22922\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \N__22919\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__22993\,
            I => \N__22916\
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__22992\,
            I => \N__22912\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__22991\,
            I => \N__22909\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__22990\,
            I => \N__22906\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__22989\,
            I => \N__22892\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__22988\,
            I => \N__22888\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__22983\,
            I => \N__22881\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__22980\,
            I => \N__22881\
        );

    \I__3356\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22866\
        );

    \I__3355\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22866\
        );

    \I__3354\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22866\
        );

    \I__3353\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22866\
        );

    \I__3352\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22866\
        );

    \I__3351\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22866\
        );

    \I__3350\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22866\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22863\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__22955\,
            I => \N__22860\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__22954\,
            I => \N__22857\
        );

    \I__3346\ : Span4Mux_v
    port map (
            O => \N__22949\,
            I => \N__22852\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__22946\,
            I => \N__22849\
        );

    \I__3344\ : Span4Mux_v
    port map (
            O => \N__22943\,
            I => \N__22844\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__22928\,
            I => \N__22844\
        );

    \I__3342\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22829\
        );

    \I__3341\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22829\
        );

    \I__3340\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22829\
        );

    \I__3339\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22829\
        );

    \I__3338\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22829\
        );

    \I__3337\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22829\
        );

    \I__3336\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22829\
        );

    \I__3335\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22814\
        );

    \I__3334\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22814\
        );

    \I__3333\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22814\
        );

    \I__3332\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22814\
        );

    \I__3331\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22814\
        );

    \I__3330\ : InMux
    port map (
            O => \N__22903\,
            I => \N__22814\
        );

    \I__3329\ : InMux
    port map (
            O => \N__22902\,
            I => \N__22814\
        );

    \I__3328\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22799\
        );

    \I__3327\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22799\
        );

    \I__3326\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22799\
        );

    \I__3325\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22799\
        );

    \I__3324\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22799\
        );

    \I__3323\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22799\
        );

    \I__3322\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22799\
        );

    \I__3321\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22788\
        );

    \I__3320\ : InMux
    port map (
            O => \N__22891\,
            I => \N__22788\
        );

    \I__3319\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22788\
        );

    \I__3318\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22788\
        );

    \I__3317\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22788\
        );

    \I__3316\ : Span4Mux_v
    port map (
            O => \N__22881\,
            I => \N__22779\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22779\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__22863\,
            I => \N__22779\
        );

    \I__3313\ : Span4Mux_h
    port map (
            O => \N__22860\,
            I => \N__22779\
        );

    \I__3312\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22772\
        );

    \I__3311\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22772\
        );

    \I__3310\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22772\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__22852\,
            I => n127_adj_2418
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__22849\,
            I => n127_adj_2418
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__22844\,
            I => n127_adj_2418
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__22829\,
            I => n127_adj_2418
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__22814\,
            I => n127_adj_2418
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__22799\,
            I => n127_adj_2418
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__22788\,
            I => n127_adj_2418
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__22779\,
            I => n127_adj_2418
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__22772\,
            I => n127_adj_2418
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__22753\,
            I => \N__22748\
        );

    \I__3299\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22745\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__22751\,
            I => \N__22742\
        );

    \I__3297\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22739\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__22745\,
            I => \N__22736\
        );

    \I__3295\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22733\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__22739\,
            I => \N__22730\
        );

    \I__3293\ : Span4Mux_v
    port map (
            O => \N__22736\,
            I => \N__22727\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__22733\,
            I => \N__22721\
        );

    \I__3291\ : Sp12to4
    port map (
            O => \N__22730\,
            I => \N__22721\
        );

    \I__3290\ : Span4Mux_v
    port map (
            O => \N__22727\,
            I => \N__22718\
        );

    \I__3289\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22715\
        );

    \I__3288\ : Odrv12
    port map (
            O => \N__22721\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__22718\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__22715\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__3285\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22683\
        );

    \I__3284\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22683\
        );

    \I__3283\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22683\
        );

    \I__3282\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22676\
        );

    \I__3281\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22676\
        );

    \I__3280\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22676\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__22702\,
            I => \N__22669\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__22701\,
            I => \N__22662\
        );

    \I__3277\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \N__22659\
        );

    \I__3276\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22652\
        );

    \I__3275\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22652\
        );

    \I__3274\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22652\
        );

    \I__3273\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22641\
        );

    \I__3272\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22641\
        );

    \I__3271\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22641\
        );

    \I__3270\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22641\
        );

    \I__3269\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22641\
        );

    \I__3268\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22636\
        );

    \I__3267\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22636\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22633\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__22676\,
            I => \N__22630\
        );

    \I__3264\ : InMux
    port map (
            O => \N__22675\,
            I => \N__22621\
        );

    \I__3263\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22621\
        );

    \I__3262\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22621\
        );

    \I__3261\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22621\
        );

    \I__3260\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22618\
        );

    \I__3259\ : InMux
    port map (
            O => \N__22668\,
            I => \N__22615\
        );

    \I__3258\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22604\
        );

    \I__3257\ : InMux
    port map (
            O => \N__22666\,
            I => \N__22604\
        );

    \I__3256\ : InMux
    port map (
            O => \N__22665\,
            I => \N__22604\
        );

    \I__3255\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22604\
        );

    \I__3254\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22604\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__22652\,
            I => \N__22599\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__22641\,
            I => \N__22599\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__22636\,
            I => \N__22594\
        );

    \I__3250\ : Span4Mux_v
    port map (
            O => \N__22633\,
            I => \N__22594\
        );

    \I__3249\ : Span4Mux_v
    port map (
            O => \N__22630\,
            I => \N__22587\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__22621\,
            I => \N__22587\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__22618\,
            I => \N__22587\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__22615\,
            I => \c0.n7212\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__22604\,
            I => \c0.n7212\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__22599\,
            I => \c0.n7212\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__22594\,
            I => \c0.n7212\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__22587\,
            I => \c0.n7212\
        );

    \I__3241\ : SRMux
    port map (
            O => \N__22576\,
            I => \N__22573\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__22573\,
            I => \N__22570\
        );

    \I__3239\ : Span12Mux_v
    port map (
            O => \N__22570\,
            I => \N__22567\
        );

    \I__3238\ : Odrv12
    port map (
            O => \N__22567\,
            I => \c0.n3_adj_2241\
        );

    \I__3237\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22560\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__22563\,
            I => \N__22557\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__22560\,
            I => \N__22554\
        );

    \I__3234\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22551\
        );

    \I__3233\ : Span4Mux_h
    port map (
            O => \N__22554\,
            I => \N__22548\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__22551\,
            I => \c0.data_in_frame_9_2\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__22548\,
            I => \c0.data_in_frame_9_2\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__22543\,
            I => \N__22540\
        );

    \I__3229\ : InMux
    port map (
            O => \N__22540\,
            I => \N__22537\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__22534\,
            I => \c0.n15939\
        );

    \I__3226\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22528\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__22528\,
            I => \N__22525\
        );

    \I__3224\ : Span4Mux_v
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__22522\,
            I => \c0.n17264\
        );

    \I__3222\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22516\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__22516\,
            I => \N__22513\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__22513\,
            I => \N__22510\
        );

    \I__3219\ : Sp12to4
    port map (
            O => \N__22510\,
            I => \N__22507\
        );

    \I__3218\ : Odrv12
    port map (
            O => \N__22507\,
            I => \c0.n9493\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__22504\,
            I => \c0.n12_cascade_\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__22501\,
            I => \N__22497\
        );

    \I__3215\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22489\
        );

    \I__3214\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22486\
        );

    \I__3213\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22483\
        );

    \I__3212\ : InMux
    port map (
            O => \N__22495\,
            I => \N__22480\
        );

    \I__3211\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22477\
        );

    \I__3210\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22474\
        );

    \I__3209\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22471\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__22489\,
            I => \N__22466\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22466\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22463\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__22480\,
            I => \N__22460\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__22477\,
            I => \N__22453\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__22474\,
            I => \N__22453\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__22471\,
            I => \N__22453\
        );

    \I__3201\ : Span4Mux_v
    port map (
            O => \N__22466\,
            I => \N__22450\
        );

    \I__3200\ : Span4Mux_h
    port map (
            O => \N__22463\,
            I => \N__22447\
        );

    \I__3199\ : Span4Mux_h
    port map (
            O => \N__22460\,
            I => \N__22442\
        );

    \I__3198\ : Span4Mux_h
    port map (
            O => \N__22453\,
            I => \N__22442\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__22450\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__22447\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__3195\ : Odrv4
    port map (
            O => \N__22442\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__3194\ : CascadeMux
    port map (
            O => \N__22435\,
            I => \n127_adj_2418_cascade_\
        );

    \I__3193\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__22429\,
            I => \c0.n17240\
        );

    \I__3191\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22422\
        );

    \I__3190\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22419\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__22422\,
            I => \N__22413\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__22419\,
            I => \N__22413\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__22418\,
            I => \N__22410\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__22413\,
            I => \N__22405\
        );

    \I__3185\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22400\
        );

    \I__3184\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22400\
        );

    \I__3183\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22397\
        );

    \I__3182\ : Sp12to4
    port map (
            O => \N__22405\,
            I => \N__22392\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__22400\,
            I => \N__22392\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__22397\,
            I => data_in_1_1
        );

    \I__3179\ : Odrv12
    port map (
            O => \N__22392\,
            I => data_in_1_1
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__22387\,
            I => \N__22384\
        );

    \I__3177\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22378\
        );

    \I__3176\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22378\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__22378\,
            I => \c0.n9482\
        );

    \I__3174\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22372\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__22372\,
            I => \N__22368\
        );

    \I__3172\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22365\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__22368\,
            I => \N__22362\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__22365\,
            I => \N__22359\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__22362\,
            I => \c0.n9490\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__22359\,
            I => \c0.n9490\
        );

    \I__3167\ : InMux
    port map (
            O => \N__22354\,
            I => \N__22350\
        );

    \I__3166\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22346\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__22350\,
            I => \N__22343\
        );

    \I__3164\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22340\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__22346\,
            I => \N__22337\
        );

    \I__3162\ : Span4Mux_h
    port map (
            O => \N__22343\,
            I => \N__22332\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__22340\,
            I => \N__22332\
        );

    \I__3160\ : Odrv12
    port map (
            O => \N__22337\,
            I => n16795
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__22332\,
            I => n16795
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__22327\,
            I => \n127_cascade_\
        );

    \I__3157\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22321\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__22321\,
            I => \N__22318\
        );

    \I__3155\ : Span4Mux_h
    port map (
            O => \N__22318\,
            I => \N__22315\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__22315\,
            I => \c0.n2\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__22312\,
            I => \c0.n2_cascade_\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__22309\,
            I => \N__22306\
        );

    \I__3151\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22303\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__22303\,
            I => \N__22300\
        );

    \I__3149\ : Span4Mux_h
    port map (
            O => \N__22300\,
            I => \N__22296\
        );

    \I__3148\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22293\
        );

    \I__3147\ : Odrv4
    port map (
            O => \N__22296\,
            I => n9435
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__22293\,
            I => n9435
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__22288\,
            I => \N__22284\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__22287\,
            I => \N__22281\
        );

    \I__3143\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22270\
        );

    \I__3142\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22270\
        );

    \I__3141\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22270\
        );

    \I__3140\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22270\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22267\
        );

    \I__3138\ : Span4Mux_s3_h
    port map (
            O => \N__22267\,
            I => \N__22264\
        );

    \I__3137\ : Span4Mux_v
    port map (
            O => \N__22264\,
            I => \N__22261\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__22261\,
            I => n7198
        );

    \I__3135\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22255\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__22255\,
            I => \N__22252\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__22252\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_18\
        );

    \I__3132\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22246\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__22246\,
            I => \N__22243\
        );

    \I__3130\ : Odrv4
    port map (
            O => \N__22243\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_18\
        );

    \I__3129\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22234\
        );

    \I__3127\ : Span4Mux_h
    port map (
            O => \N__22234\,
            I => \N__22231\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__22231\,
            I => \c0.n12_adj_2158\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__22228\,
            I => \c0.n9488_cascade_\
        );

    \I__3124\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22222\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__22222\,
            I => \N__22219\
        );

    \I__3122\ : Span4Mux_h
    port map (
            O => \N__22219\,
            I => \N__22216\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__22216\,
            I => \c0.n17262\
        );

    \I__3120\ : InMux
    port map (
            O => \N__22213\,
            I => \N__22210\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__22210\,
            I => \c0.n17256\
        );

    \I__3118\ : InMux
    port map (
            O => \N__22207\,
            I => \N__22200\
        );

    \I__3117\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22200\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__22205\,
            I => \N__22197\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__22200\,
            I => \N__22194\
        );

    \I__3114\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22191\
        );

    \I__3113\ : Span4Mux_v
    port map (
            O => \N__22194\,
            I => \N__22188\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__22191\,
            I => data_in_0_0
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__22188\,
            I => data_in_0_0
        );

    \I__3110\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22179\
        );

    \I__3109\ : InMux
    port map (
            O => \N__22182\,
            I => \N__22176\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__22179\,
            I => \c0.n9485\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__22176\,
            I => \c0.n9485\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__22171\,
            I => \c0.n10_adj_2149_cascade_\
        );

    \I__3105\ : InMux
    port map (
            O => \N__22168\,
            I => \N__22165\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__22165\,
            I => \N__22159\
        );

    \I__3103\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22156\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__22163\,
            I => \N__22153\
        );

    \I__3101\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22150\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__22159\,
            I => \N__22147\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__22156\,
            I => \N__22144\
        );

    \I__3098\ : InMux
    port map (
            O => \N__22153\,
            I => \N__22141\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__22150\,
            I => \N__22138\
        );

    \I__3096\ : Span4Mux_v
    port map (
            O => \N__22147\,
            I => \N__22135\
        );

    \I__3095\ : Span4Mux_h
    port map (
            O => \N__22144\,
            I => \N__22132\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__22141\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__3093\ : Odrv12
    port map (
            O => \N__22138\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__22135\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__22132\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__3090\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22120\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__22120\,
            I => \N__22117\
        );

    \I__3088\ : Span4Mux_h
    port map (
            O => \N__22117\,
            I => \N__22114\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__22114\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_29\
        );

    \I__3086\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22107\
        );

    \I__3085\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22103\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__22107\,
            I => \N__22100\
        );

    \I__3083\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22096\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__22103\,
            I => \N__22091\
        );

    \I__3081\ : Span4Mux_h
    port map (
            O => \N__22100\,
            I => \N__22091\
        );

    \I__3080\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22088\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__22096\,
            I => data_in_3_0
        );

    \I__3078\ : Odrv4
    port map (
            O => \N__22091\,
            I => data_in_3_0
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__22088\,
            I => data_in_3_0
        );

    \I__3076\ : InMux
    port map (
            O => \N__22081\,
            I => \N__22078\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__22074\
        );

    \I__3074\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22070\
        );

    \I__3073\ : Span4Mux_h
    port map (
            O => \N__22074\,
            I => \N__22067\
        );

    \I__3072\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22064\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__22070\,
            I => data_in_0_5
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__22067\,
            I => data_in_0_5
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__22064\,
            I => data_in_0_5
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__22057\,
            I => \N__22054\
        );

    \I__3067\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22050\
        );

    \I__3066\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22045\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__22050\,
            I => \N__22042\
        );

    \I__3064\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22037\
        );

    \I__3063\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22037\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__22045\,
            I => data_in_3_4
        );

    \I__3061\ : Odrv4
    port map (
            O => \N__22042\,
            I => data_in_3_4
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__22037\,
            I => data_in_3_4
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__22030\,
            I => \c0.n9451_cascade_\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__22027\,
            I => \n12933_cascade_\
        );

    \I__3057\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22021\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__22016\
        );

    \I__3055\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22010\
        );

    \I__3054\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22010\
        );

    \I__3053\ : Span4Mux_h
    port map (
            O => \N__22016\,
            I => \N__22005\
        );

    \I__3052\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22002\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__21999\
        );

    \I__3050\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21994\
        );

    \I__3049\ : InMux
    port map (
            O => \N__22008\,
            I => \N__21994\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__22005\,
            I => \c0.n9451\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__22002\,
            I => \c0.n9451\
        );

    \I__3046\ : Odrv12
    port map (
            O => \N__21999\,
            I => \c0.n9451\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__21994\,
            I => \c0.n9451\
        );

    \I__3044\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21982\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__21982\,
            I => \N__21979\
        );

    \I__3042\ : Span4Mux_v
    port map (
            O => \N__21979\,
            I => \N__21976\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__21976\,
            I => \c0.n9\
        );

    \I__3040\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21970\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__21970\,
            I => \c0.n17258\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__21967\,
            I => \c0.n28_cascade_\
        );

    \I__3037\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21961\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__21961\,
            I => \c0.n60\
        );

    \I__3035\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21955\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__21955\,
            I => \c0.n16879\
        );

    \I__3033\ : InMux
    port map (
            O => \N__21952\,
            I => \N__21949\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__21949\,
            I => \N__21945\
        );

    \I__3031\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21942\
        );

    \I__3030\ : Span4Mux_v
    port map (
            O => \N__21945\,
            I => \N__21939\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__21942\,
            I => \N__21936\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__21939\,
            I => \N__21931\
        );

    \I__3027\ : Span4Mux_h
    port map (
            O => \N__21936\,
            I => \N__21931\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__21931\,
            I => \c0.n33\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__21928\,
            I => \c0.n16879_cascade_\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__21925\,
            I => \N__21922\
        );

    \I__3023\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21919\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21915\
        );

    \I__3021\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21912\
        );

    \I__3020\ : Span4Mux_v
    port map (
            O => \N__21915\,
            I => \N__21907\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__21912\,
            I => \N__21907\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__21907\,
            I => \N__21902\
        );

    \I__3017\ : InMux
    port map (
            O => \N__21906\,
            I => \N__21899\
        );

    \I__3016\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21896\
        );

    \I__3015\ : Span4Mux_s3_h
    port map (
            O => \N__21902\,
            I => \N__21893\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__21899\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__21896\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__21893\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__21886\,
            I => \N__21881\
        );

    \I__3010\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21877\
        );

    \I__3009\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21874\
        );

    \I__3008\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21871\
        );

    \I__3007\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21868\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__21877\,
            I => \N__21865\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__21874\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__21871\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__21868\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__21865\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__21856\,
            I => \N__21852\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__21855\,
            I => \N__21848\
        );

    \I__2999\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21842\
        );

    \I__2998\ : InMux
    port map (
            O => \N__21851\,
            I => \N__21842\
        );

    \I__2997\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21839\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__21847\,
            I => \N__21836\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__21842\,
            I => \N__21831\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__21839\,
            I => \N__21831\
        );

    \I__2993\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21828\
        );

    \I__2992\ : Span4Mux_v
    port map (
            O => \N__21831\,
            I => \N__21825\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__21828\,
            I => \N__21822\
        );

    \I__2990\ : Span4Mux_h
    port map (
            O => \N__21825\,
            I => \N__21819\
        );

    \I__2989\ : Span4Mux_h
    port map (
            O => \N__21822\,
            I => \N__21816\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__21819\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__21816\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__2986\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21807\
        );

    \I__2985\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21804\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__21807\,
            I => n9445
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__21804\,
            I => n9445
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__21799\,
            I => \N__21796\
        );

    \I__2981\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21793\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__21793\,
            I => \N__21790\
        );

    \I__2979\ : Odrv4
    port map (
            O => \N__21790\,
            I => \c0.n9488\
        );

    \I__2978\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21778\
        );

    \I__2977\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21778\
        );

    \I__2976\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21778\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__21778\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__2974\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21771\
        );

    \I__2973\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21767\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__21771\,
            I => \N__21764\
        );

    \I__2971\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21761\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__21767\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__2969\ : Odrv12
    port map (
            O => \N__21764\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__21761\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__2967\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21749\
        );

    \I__2966\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21746\
        );

    \I__2965\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21743\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__21749\,
            I => \N__21738\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__21746\,
            I => \N__21738\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__21743\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__2961\ : Odrv12
    port map (
            O => \N__21738\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__21733\,
            I => \c0.n59_cascade_\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__21730\,
            I => \c0.n5_adj_2262_cascade_\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__21727\,
            I => \c0.n16876_cascade_\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__21724\,
            I => \c0.n60_cascade_\
        );

    \I__2956\ : SRMux
    port map (
            O => \N__21721\,
            I => \N__21718\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__21718\,
            I => \N__21715\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__21715\,
            I => \c0.n16363\
        );

    \I__2953\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21707\
        );

    \I__2952\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21704\
        );

    \I__2951\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21701\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__21707\,
            I => \N__21698\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__21704\,
            I => \N__21695\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__21701\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__2947\ : Odrv4
    port map (
            O => \N__21698\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__2946\ : Odrv12
    port map (
            O => \N__21695\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__2945\ : InMux
    port map (
            O => \N__21688\,
            I => \N__21679\
        );

    \I__2944\ : InMux
    port map (
            O => \N__21687\,
            I => \N__21679\
        );

    \I__2943\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21679\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__21679\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__2941\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21673\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__21673\,
            I => \N__21669\
        );

    \I__2939\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21666\
        );

    \I__2938\ : Span4Mux_h
    port map (
            O => \N__21669\,
            I => \N__21663\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__21666\,
            I => n9453
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__21663\,
            I => n9453
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__21658\,
            I => \N__21654\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__21657\,
            I => \N__21649\
        );

    \I__2933\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21646\
        );

    \I__2932\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21643\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__21652\,
            I => \N__21637\
        );

    \I__2930\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21634\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__21646\,
            I => \N__21628\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21628\
        );

    \I__2927\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21625\
        );

    \I__2926\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21618\
        );

    \I__2925\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21618\
        );

    \I__2924\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21618\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__21634\,
            I => \N__21615\
        );

    \I__2922\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21612\
        );

    \I__2921\ : Span4Mux_v
    port map (
            O => \N__21628\,
            I => \N__21607\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__21625\,
            I => \N__21607\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__21618\,
            I => \N__21602\
        );

    \I__2918\ : Span4Mux_v
    port map (
            O => \N__21615\,
            I => \N__21602\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__21612\,
            I => \N__21597\
        );

    \I__2916\ : Span4Mux_v
    port map (
            O => \N__21607\,
            I => \N__21597\
        );

    \I__2915\ : Span4Mux_h
    port map (
            O => \N__21602\,
            I => \N__21594\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__21597\,
            I => \N__21591\
        );

    \I__2913\ : Span4Mux_s1_h
    port map (
            O => \N__21594\,
            I => \N__21588\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__21591\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__21588\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__2910\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21579\
        );

    \I__2909\ : CascadeMux
    port map (
            O => \N__21582\,
            I => \N__21576\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__21579\,
            I => \N__21573\
        );

    \I__2907\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21570\
        );

    \I__2906\ : Span4Mux_s3_h
    port map (
            O => \N__21573\,
            I => \N__21567\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__21570\,
            I => \N__21564\
        );

    \I__2904\ : Odrv4
    port map (
            O => \N__21567\,
            I => n2275
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__21564\,
            I => n2275
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__21559\,
            I => \n2275_cascade_\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__21556\,
            I => \c0.n7212_cascade_\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__21553\,
            I => \c0.n17452_cascade_\
        );

    \I__2899\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21547\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__21547\,
            I => \c0.n17454\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__21544\,
            I => \c0.n7_cascade_\
        );

    \I__2896\ : SRMux
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__21538\,
            I => \N__21535\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__21535\,
            I => \c0.n16335\
        );

    \I__2893\ : SRMux
    port map (
            O => \N__21532\,
            I => \N__21529\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21526\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__21526\,
            I => \N__21523\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__21523\,
            I => \c0.n16381\
        );

    \I__2889\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21515\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__21519\,
            I => \N__21511\
        );

    \I__2887\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21508\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__21515\,
            I => \N__21505\
        );

    \I__2885\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21502\
        );

    \I__2884\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21499\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__21508\,
            I => \N__21496\
        );

    \I__2882\ : Span4Mux_v
    port map (
            O => \N__21505\,
            I => \N__21493\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__21502\,
            I => \N__21488\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__21499\,
            I => \N__21488\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__21496\,
            I => \N__21485\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__21493\,
            I => \N__21480\
        );

    \I__2877\ : Span4Mux_v
    port map (
            O => \N__21488\,
            I => \N__21480\
        );

    \I__2876\ : Span4Mux_h
    port map (
            O => \N__21485\,
            I => \N__21477\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__21480\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__21477\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__21472\,
            I => \N__21467\
        );

    \I__2872\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21463\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21460\
        );

    \I__2870\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21457\
        );

    \I__2869\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21454\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__21463\,
            I => \N__21451\
        );

    \I__2867\ : InMux
    port map (
            O => \N__21460\,
            I => \N__21448\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__21457\,
            I => \N__21445\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__21454\,
            I => \N__21442\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__21451\,
            I => \N__21439\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__21448\,
            I => \N__21436\
        );

    \I__2862\ : Span12Mux_s9_v
    port map (
            O => \N__21445\,
            I => \N__21433\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__21442\,
            I => \N__21426\
        );

    \I__2860\ : Span4Mux_v
    port map (
            O => \N__21439\,
            I => \N__21426\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__21436\,
            I => \N__21426\
        );

    \I__2858\ : Odrv12
    port map (
            O => \N__21433\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__21426\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__2856\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21418\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__21418\,
            I => \N__21415\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__21415\,
            I => \N__21412\
        );

    \I__2853\ : Span4Mux_v
    port map (
            O => \N__21412\,
            I => \N__21409\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__21409\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_16\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__21406\,
            I => \n1716_cascade_\
        );

    \I__2850\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21400\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__21400\,
            I => n14
        );

    \I__2848\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21394\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__21394\,
            I => \N__21391\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__21391\,
            I => n16775
        );

    \I__2845\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21384\
        );

    \I__2844\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21381\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__21384\,
            I => \N__21378\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__21381\,
            I => \N__21375\
        );

    \I__2841\ : Span4Mux_h
    port map (
            O => \N__21378\,
            I => \N__21372\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__21375\,
            I => n3977
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__21372\,
            I => n3977
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__21367\,
            I => \n16775_cascade_\
        );

    \I__2837\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21360\
        );

    \I__2836\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21356\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__21360\,
            I => \N__21353\
        );

    \I__2834\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21350\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__21356\,
            I => \c0.delay_counter_10\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__21353\,
            I => \c0.delay_counter_10\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__21350\,
            I => \c0.delay_counter_10\
        );

    \I__2830\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21340\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__21340\,
            I => \N__21337\
        );

    \I__2828\ : Odrv12
    port map (
            O => \N__21337\,
            I => \c0.n6522\
        );

    \I__2827\ : InMux
    port map (
            O => \N__21334\,
            I => \c0.n15523\
        );

    \I__2826\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21328\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21323\
        );

    \I__2824\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21318\
        );

    \I__2823\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21318\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__21323\,
            I => \c0.delay_counter_11\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__21318\,
            I => \c0.delay_counter_11\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__21313\,
            I => \N__21310\
        );

    \I__2819\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21307\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21304\
        );

    \I__2817\ : Span4Mux_v
    port map (
            O => \N__21304\,
            I => \N__21301\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__21301\,
            I => \c0.n6521\
        );

    \I__2815\ : InMux
    port map (
            O => \N__21298\,
            I => \c0.n15524\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__21295\,
            I => \N__21292\
        );

    \I__2813\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21286\
        );

    \I__2812\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21283\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__21290\,
            I => \N__21280\
        );

    \I__2810\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21277\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__21286\,
            I => \N__21274\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__21283\,
            I => \N__21271\
        );

    \I__2807\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21268\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__21277\,
            I => \c0.delay_counter_12\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__21274\,
            I => \c0.delay_counter_12\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__21271\,
            I => \c0.delay_counter_12\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__21268\,
            I => \c0.delay_counter_12\
        );

    \I__2802\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21256\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__21256\,
            I => \N__21253\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__21253\,
            I => \c0.n17575\
        );

    \I__2799\ : InMux
    port map (
            O => \N__21250\,
            I => \c0.n15525\
        );

    \I__2798\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21244\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21241\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__21241\,
            I => \c0.n17639\
        );

    \I__2795\ : InMux
    port map (
            O => \N__21238\,
            I => \c0.n15526\
        );

    \I__2794\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21230\
        );

    \I__2793\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21227\
        );

    \I__2792\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21224\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__21230\,
            I => \N__21221\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__21227\,
            I => \N__21217\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21212\
        );

    \I__2788\ : Span4Mux_s2_v
    port map (
            O => \N__21221\,
            I => \N__21212\
        );

    \I__2787\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21209\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__21217\,
            I => \c0.delay_counter_14\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__21212\,
            I => \c0.delay_counter_14\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__21209\,
            I => \c0.delay_counter_14\
        );

    \I__2783\ : InMux
    port map (
            O => \N__21202\,
            I => \c0.n15527\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__21199\,
            I => \N__21196\
        );

    \I__2781\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21193\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__21193\,
            I => \N__21190\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__21190\,
            I => \c0.n17635\
        );

    \I__2778\ : SRMux
    port map (
            O => \N__21187\,
            I => \N__21184\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__21184\,
            I => \N__21181\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__21181\,
            I => \c0.n16331\
        );

    \I__2775\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21175\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__21175\,
            I => \c0.n6530\
        );

    \I__2773\ : InMux
    port map (
            O => \N__21172\,
            I => \c0.n15515\
        );

    \I__2772\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21164\
        );

    \I__2771\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21159\
        );

    \I__2770\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21159\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__21164\,
            I => \c0.delay_counter_3\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__21159\,
            I => \c0.delay_counter_3\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__21154\,
            I => \N__21151\
        );

    \I__2766\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21148\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__21148\,
            I => \c0.n6529\
        );

    \I__2764\ : InMux
    port map (
            O => \N__21145\,
            I => \c0.n15516\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__21142\,
            I => \N__21139\
        );

    \I__2762\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21136\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__21136\,
            I => \c0.n6528\
        );

    \I__2760\ : InMux
    port map (
            O => \N__21133\,
            I => \c0.n15517\
        );

    \I__2759\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21124\
        );

    \I__2758\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21121\
        );

    \I__2757\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21118\
        );

    \I__2756\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21115\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__21124\,
            I => \c0.delay_counter_5\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__21121\,
            I => \c0.delay_counter_5\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__21118\,
            I => \c0.delay_counter_5\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__21115\,
            I => \c0.delay_counter_5\
        );

    \I__2751\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21103\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__21103\,
            I => \c0.n17574\
        );

    \I__2749\ : InMux
    port map (
            O => \N__21100\,
            I => \c0.n15518\
        );

    \I__2748\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21092\
        );

    \I__2747\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21089\
        );

    \I__2746\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21086\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__21092\,
            I => \N__21083\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__21089\,
            I => \c0.delay_counter_6\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__21086\,
            I => \c0.delay_counter_6\
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__21083\,
            I => \c0.delay_counter_6\
        );

    \I__2741\ : InMux
    port map (
            O => \N__21076\,
            I => \N__21073\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__21073\,
            I => \c0.n6526\
        );

    \I__2739\ : InMux
    port map (
            O => \N__21070\,
            I => \c0.n15519\
        );

    \I__2738\ : InMux
    port map (
            O => \N__21067\,
            I => \N__21061\
        );

    \I__2737\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21058\
        );

    \I__2736\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21055\
        );

    \I__2735\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21052\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__21061\,
            I => \c0.delay_counter_7\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__21058\,
            I => \c0.delay_counter_7\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__21055\,
            I => \c0.delay_counter_7\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__21052\,
            I => \c0.delay_counter_7\
        );

    \I__2730\ : InMux
    port map (
            O => \N__21043\,
            I => \N__21040\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__21040\,
            I => \c0.n17638\
        );

    \I__2728\ : InMux
    port map (
            O => \N__21037\,
            I => \c0.n15520\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__21034\,
            I => \N__21031\
        );

    \I__2726\ : InMux
    port map (
            O => \N__21031\,
            I => \N__21028\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__21028\,
            I => \N__21025\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__21025\,
            I => \c0.n6524\
        );

    \I__2723\ : InMux
    port map (
            O => \N__21022\,
            I => \bfn_5_32_0_\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21019\,
            I => \N__21014\
        );

    \I__2721\ : InMux
    port map (
            O => \N__21018\,
            I => \N__21011\
        );

    \I__2720\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21008\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__21014\,
            I => \c0.delay_counter_9\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__21011\,
            I => \c0.delay_counter_9\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21008\,
            I => \c0.delay_counter_9\
        );

    \I__2716\ : InMux
    port map (
            O => \N__21001\,
            I => \N__20998\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__20998\,
            I => \c0.n6523\
        );

    \I__2714\ : InMux
    port map (
            O => \N__20995\,
            I => \c0.n15522\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__20992\,
            I => \c0.n1419_cascade_\
        );

    \I__2712\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20971\
        );

    \I__2711\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20971\
        );

    \I__2710\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20964\
        );

    \I__2709\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20964\
        );

    \I__2708\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20964\
        );

    \I__2707\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20957\
        );

    \I__2706\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20957\
        );

    \I__2705\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20957\
        );

    \I__2704\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20944\
        );

    \I__2703\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20944\
        );

    \I__2702\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20944\
        );

    \I__2701\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20944\
        );

    \I__2700\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20944\
        );

    \I__2699\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20944\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__20971\,
            I => \c0.n1419\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__20964\,
            I => \c0.n1419\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__20957\,
            I => \c0.n1419\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__20944\,
            I => \c0.n1419\
        );

    \I__2694\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20932\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__20932\,
            I => n53
        );

    \I__2692\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20925\
        );

    \I__2691\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20920\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__20925\,
            I => \N__20917\
        );

    \I__2689\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20914\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__20923\,
            I => \N__20911\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__20920\,
            I => \N__20906\
        );

    \I__2686\ : Span4Mux_s3_v
    port map (
            O => \N__20917\,
            I => \N__20906\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20903\
        );

    \I__2684\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20900\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__20906\,
            I => \c0.delay_counter_0\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__20903\,
            I => \c0.delay_counter_0\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__20900\,
            I => \c0.delay_counter_0\
        );

    \I__2680\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20890\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__20890\,
            I => \N__20887\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__20887\,
            I => \c0.n17637\
        );

    \I__2677\ : InMux
    port map (
            O => \N__20884\,
            I => \bfn_5_31_0_\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__20881\,
            I => \N__20878\
        );

    \I__2675\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20873\
        );

    \I__2674\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20870\
        );

    \I__2673\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20867\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__20873\,
            I => \c0.delay_counter_1\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__20870\,
            I => \c0.delay_counter_1\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__20867\,
            I => \c0.delay_counter_1\
        );

    \I__2669\ : InMux
    port map (
            O => \N__20860\,
            I => \N__20857\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__20857\,
            I => \c0.n6531\
        );

    \I__2667\ : InMux
    port map (
            O => \N__20854\,
            I => \c0.n15514\
        );

    \I__2666\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20842\
        );

    \I__2665\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20839\
        );

    \I__2664\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20830\
        );

    \I__2663\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20830\
        );

    \I__2662\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20830\
        );

    \I__2661\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20830\
        );

    \I__2660\ : InMux
    port map (
            O => \N__20845\,
            I => \N__20827\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__20842\,
            I => n16893
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__20839\,
            I => n16893
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__20830\,
            I => n16893
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__20827\,
            I => n16893
        );

    \I__2655\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20815\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__20815\,
            I => \c0.tx.n17462\
        );

    \I__2653\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20805\
        );

    \I__2652\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20802\
        );

    \I__2651\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20799\
        );

    \I__2650\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20796\
        );

    \I__2649\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20793\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20790\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__20802\,
            I => \N__20783\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__20799\,
            I => \N__20783\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__20796\,
            I => \N__20783\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__20793\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__2643\ : Odrv12
    port map (
            O => \N__20790\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__20783\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__2641\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20773\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__20773\,
            I => \N__20770\
        );

    \I__2639\ : Span4Mux_h
    port map (
            O => \N__20770\,
            I => \N__20767\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__20767\,
            I => n17397
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__20764\,
            I => \N__20758\
        );

    \I__2636\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20755\
        );

    \I__2635\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20750\
        );

    \I__2634\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20750\
        );

    \I__2633\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20747\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__20755\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__20750\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__20747\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__20740\,
            I => \c0.tx.n17975_cascade_\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__20737\,
            I => \c0.tx.o_Tx_Serial_N_2064_cascade_\
        );

    \I__2627\ : InMux
    port map (
            O => \N__20734\,
            I => \N__20731\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__20731\,
            I => \N__20728\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__20728\,
            I => n3_adj_2406
        );

    \I__2624\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20722\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20719\
        );

    \I__2622\ : Span4Mux_h
    port map (
            O => \N__20719\,
            I => \N__20715\
        );

    \I__2621\ : InMux
    port map (
            O => \N__20718\,
            I => \N__20712\
        );

    \I__2620\ : Span4Mux_v
    port map (
            O => \N__20715\,
            I => \N__20709\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__20712\,
            I => \N__20706\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__20709\,
            I => n13082
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__20706\,
            I => n13082
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__20701\,
            I => \c0.n16891_cascade_\
        );

    \I__2615\ : InMux
    port map (
            O => \N__20698\,
            I => \N__20694\
        );

    \I__2614\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20690\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__20694\,
            I => \N__20687\
        );

    \I__2612\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20682\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__20690\,
            I => \N__20679\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__20687\,
            I => \N__20676\
        );

    \I__2609\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20671\
        );

    \I__2608\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20671\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__20682\,
            I => \r_Bit_Index_0\
        );

    \I__2606\ : Odrv12
    port map (
            O => \N__20679\,
            I => \r_Bit_Index_0\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__20676\,
            I => \r_Bit_Index_0\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__20671\,
            I => \r_Bit_Index_0\
        );

    \I__2603\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20659\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__20659\,
            I => \N__20655\
        );

    \I__2601\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20652\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__20655\,
            I => \c0.rx.n9323\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__20652\,
            I => \c0.rx.n9323\
        );

    \I__2598\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20641\
        );

    \I__2597\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20641\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__20641\,
            I => \N__20637\
        );

    \I__2595\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20634\
        );

    \I__2594\ : Odrv12
    port map (
            O => \N__20637\,
            I => n9477
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__20634\,
            I => n9477
        );

    \I__2592\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20626\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__20626\,
            I => \N__20622\
        );

    \I__2590\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20619\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__20622\,
            I => n4_adj_2409
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__20619\,
            I => n4_adj_2409
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__20614\,
            I => \n9477_cascade_\
        );

    \I__2586\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20607\
        );

    \I__2585\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20604\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__20607\,
            I => data_in_0_2
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__20604\,
            I => data_in_0_2
        );

    \I__2582\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20596\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__20596\,
            I => \N__20591\
        );

    \I__2580\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20586\
        );

    \I__2579\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20586\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__20591\,
            I => data_in_1_3
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__20586\,
            I => data_in_1_3
        );

    \I__2576\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20578\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__20578\,
            I => \N__20575\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__20575\,
            I => \c0.n12_adj_2200\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__20572\,
            I => \N__20569\
        );

    \I__2572\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20566\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__20566\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_31\
        );

    \I__2570\ : InMux
    port map (
            O => \N__20563\,
            I => \N__20559\
        );

    \I__2569\ : InMux
    port map (
            O => \N__20562\,
            I => \N__20556\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__20559\,
            I => \N__20553\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__20556\,
            I => \N__20550\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__20553\,
            I => \N__20547\
        );

    \I__2565\ : Span4Mux_h
    port map (
            O => \N__20550\,
            I => \N__20544\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__20547\,
            I => n4_adj_2460
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__20544\,
            I => n4_adj_2460
        );

    \I__2562\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20536\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__20536\,
            I => \N__20532\
        );

    \I__2560\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20529\
        );

    \I__2559\ : Span4Mux_h
    port map (
            O => \N__20532\,
            I => \N__20524\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__20529\,
            I => \N__20524\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__20524\,
            I => n4_adj_2417
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__20521\,
            I => \c0.n127_adj_2136_cascade_\
        );

    \I__2555\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20515\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__20515\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_27\
        );

    \I__2553\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20509\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__20509\,
            I => \N__20504\
        );

    \I__2551\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20499\
        );

    \I__2550\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20499\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__20504\,
            I => \N__20496\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__20499\,
            I => \N__20493\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__20496\,
            I => n9472
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__20493\,
            I => n9472
        );

    \I__2545\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20485\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__20485\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_30\
        );

    \I__2543\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20479\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__20479\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_25\
        );

    \I__2541\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20473\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__20473\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_28\
        );

    \I__2539\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__20467\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_24\
        );

    \I__2537\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__20461\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_26\
        );

    \I__2535\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20455\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__20455\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_22\
        );

    \I__2533\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20449\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__20449\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_9\
        );

    \I__2531\ : SRMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__20443\,
            I => \N__20440\
        );

    \I__2529\ : Span4Mux_h
    port map (
            O => \N__20440\,
            I => \N__20437\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__20437\,
            I => \c0.n3_adj_2248\
        );

    \I__2527\ : InMux
    port map (
            O => \N__20434\,
            I => \N__20431\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__20431\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_8\
        );

    \I__2525\ : InMux
    port map (
            O => \N__20428\,
            I => \N__20425\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__20425\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_19\
        );

    \I__2523\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20419\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__20419\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_20\
        );

    \I__2521\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20413\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__20413\,
            I => \N__20410\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__20410\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_21\
        );

    \I__2518\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20404\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__20404\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_23\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__20401\,
            I => \c0.n18_adj_2198_cascade_\
        );

    \I__2515\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__20395\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_6\
        );

    \I__2513\ : SRMux
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__20389\,
            I => \c0.n3_adj_2253\
        );

    \I__2511\ : SRMux
    port map (
            O => \N__20386\,
            I => \N__20383\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__20383\,
            I => \N__20380\
        );

    \I__2509\ : Span4Mux_h
    port map (
            O => \N__20380\,
            I => \N__20377\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__20377\,
            I => \c0.n3_adj_2237\
        );

    \I__2507\ : SRMux
    port map (
            O => \N__20374\,
            I => \N__20371\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__20371\,
            I => \N__20368\
        );

    \I__2505\ : Span4Mux_s1_h
    port map (
            O => \N__20368\,
            I => \N__20365\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__20365\,
            I => \N__20362\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__20362\,
            I => \c0.n3_adj_2235\
        );

    \I__2502\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20356\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__20356\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_11\
        );

    \I__2500\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20350\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__20350\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_11\
        );

    \I__2498\ : SRMux
    port map (
            O => \N__20347\,
            I => \N__20344\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__20344\,
            I => \N__20341\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__20341\,
            I => \c0.n3_adj_2246\
        );

    \I__2495\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20335\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__20335\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_10\
        );

    \I__2493\ : SRMux
    port map (
            O => \N__20332\,
            I => \N__20329\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__20329\,
            I => \N__20326\
        );

    \I__2491\ : Span4Mux_v
    port map (
            O => \N__20326\,
            I => \N__20323\
        );

    \I__2490\ : Span4Mux_s1_h
    port map (
            O => \N__20323\,
            I => \N__20320\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__20320\,
            I => \c0.n3_adj_2231\
        );

    \I__2488\ : SRMux
    port map (
            O => \N__20317\,
            I => \N__20314\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__20314\,
            I => \N__20311\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__20311\,
            I => \N__20308\
        );

    \I__2485\ : Span4Mux_v
    port map (
            O => \N__20308\,
            I => \N__20305\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__20305\,
            I => \c0.n3_adj_2227\
        );

    \I__2483\ : SRMux
    port map (
            O => \N__20302\,
            I => \N__20299\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20296\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__20296\,
            I => \N__20293\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__20293\,
            I => \c0.n3_adj_2223\
        );

    \I__2479\ : SRMux
    port map (
            O => \N__20290\,
            I => \N__20287\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__20287\,
            I => \N__20284\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__20284\,
            I => \N__20281\
        );

    \I__2476\ : Span4Mux_s2_h
    port map (
            O => \N__20281\,
            I => \N__20278\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__20278\,
            I => \c0.n3_adj_2225\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__20275\,
            I => \c0.n1439_cascade_\
        );

    \I__2473\ : SRMux
    port map (
            O => \N__20272\,
            I => \N__20269\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__20269\,
            I => \N__20266\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__20266\,
            I => \N__20263\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__20263\,
            I => \N__20260\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__20260\,
            I => \c0.n3_adj_2221\
        );

    \I__2468\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20254\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__20254\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_7\
        );

    \I__2466\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20248\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__20248\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_7\
        );

    \I__2464\ : SRMux
    port map (
            O => \N__20245\,
            I => \N__20242\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__20242\,
            I => \N__20239\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__20239\,
            I => \c0.n3_adj_2250\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__20236\,
            I => \n3977_cascade_\
        );

    \I__2460\ : SRMux
    port map (
            O => \N__20233\,
            I => \N__20230\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__20230\,
            I => \c0.n3_adj_2233\
        );

    \I__2458\ : SRMux
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__20224\,
            I => \N__20221\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__20221\,
            I => \c0.n3_adj_2219\
        );

    \I__2455\ : SRMux
    port map (
            O => \N__20218\,
            I => \N__20215\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__20215\,
            I => \N__20212\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__20212\,
            I => \N__20209\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__20209\,
            I => \c0.n16441\
        );

    \I__2451\ : SRMux
    port map (
            O => \N__20206\,
            I => \N__20203\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__20203\,
            I => \N__20200\
        );

    \I__2449\ : Span4Mux_s2_h
    port map (
            O => \N__20200\,
            I => \N__20197\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__20197\,
            I => \c0.n3_adj_2229\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__20194\,
            I => \n29_cascade_\
        );

    \I__2446\ : IoInMux
    port map (
            O => \N__20191\,
            I => \N__20188\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__20188\,
            I => tx_enable
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__20185\,
            I => \N__20182\
        );

    \I__2443\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20179\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__20179\,
            I => \c0.n12991\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__20176\,
            I => \c0.n12991_cascade_\
        );

    \I__2440\ : InMux
    port map (
            O => \N__20173\,
            I => \N__20170\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__20170\,
            I => \c0.n19_adj_2270\
        );

    \I__2438\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20164\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__20164\,
            I => \N__20161\
        );

    \I__2436\ : Odrv4
    port map (
            O => \N__20161\,
            I => n16859
        );

    \I__2435\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20155\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__20155\,
            I => \N__20151\
        );

    \I__2433\ : InMux
    port map (
            O => \N__20154\,
            I => \N__20148\
        );

    \I__2432\ : Span4Mux_v
    port map (
            O => \N__20151\,
            I => \N__20142\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__20148\,
            I => \N__20142\
        );

    \I__2430\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20134\
        );

    \I__2429\ : Span4Mux_s2_v
    port map (
            O => \N__20142\,
            I => \N__20131\
        );

    \I__2428\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20126\
        );

    \I__2427\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20126\
        );

    \I__2426\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20123\
        );

    \I__2425\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20120\
        );

    \I__2424\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20117\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__20134\,
            I => \N__20114\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__20131\,
            I => n17_adj_2416
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__20126\,
            I => n17_adj_2416
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__20123\,
            I => n17_adj_2416
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__20120\,
            I => n17_adj_2416
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__20117\,
            I => n17_adj_2416
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__20114\,
            I => n17_adj_2416
        );

    \I__2416\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20097\
        );

    \I__2415\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20093\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__20097\,
            I => \N__20090\
        );

    \I__2413\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20087\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__20093\,
            I => \N__20084\
        );

    \I__2411\ : Span4Mux_s3_h
    port map (
            O => \N__20090\,
            I => \N__20081\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__20087\,
            I => \r_Clock_Count_0_adj_2437\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__20084\,
            I => \r_Clock_Count_0_adj_2437\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__20081\,
            I => \r_Clock_Count_0_adj_2437\
        );

    \I__2407\ : IoInMux
    port map (
            O => \N__20074\,
            I => \N__20069\
        );

    \I__2406\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20064\
        );

    \I__2405\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20064\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__20069\,
            I => tx_o
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__20064\,
            I => tx_o
        );

    \I__2402\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20056\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__20056\,
            I => \N__20053\
        );

    \I__2400\ : Span4Mux_h
    port map (
            O => \N__20053\,
            I => \N__20049\
        );

    \I__2399\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20045\
        );

    \I__2398\ : Sp12to4
    port map (
            O => \N__20049\,
            I => \N__20042\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20048\,
            I => \N__20039\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__20045\,
            I => data_in_1_0
        );

    \I__2395\ : Odrv12
    port map (
            O => \N__20042\,
            I => data_in_1_0
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__20039\,
            I => data_in_1_0
        );

    \I__2393\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20029\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__20029\,
            I => \c0.n12993\
        );

    \I__2391\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20022\
        );

    \I__2390\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20019\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__20022\,
            I => \c0.n13298\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__20019\,
            I => \c0.n13298\
        );

    \I__2387\ : InMux
    port map (
            O => \N__20014\,
            I => \N__20011\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__20011\,
            I => \c0.n20_adj_2267\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__20008\,
            I => \c0.n21_adj_2271_cascade_\
        );

    \I__2384\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19998\
        );

    \I__2383\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19995\
        );

    \I__2382\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19990\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19990\
        );

    \I__2380\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19987\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__19998\,
            I => \N__19984\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__19995\,
            I => \r_SM_Main_2_N_2033_1\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__19990\,
            I => \r_SM_Main_2_N_2033_1\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__19987\,
            I => \r_SM_Main_2_N_2033_1\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__19984\,
            I => \r_SM_Main_2_N_2033_1\
        );

    \I__2374\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19972\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__19972\,
            I => \N__19966\
        );

    \I__2372\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19963\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__19970\,
            I => \N__19958\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__19969\,
            I => \N__19954\
        );

    \I__2369\ : Sp12to4
    port map (
            O => \N__19966\,
            I => \N__19949\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__19963\,
            I => \N__19949\
        );

    \I__2367\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19946\
        );

    \I__2366\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19941\
        );

    \I__2365\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19941\
        );

    \I__2364\ : InMux
    port map (
            O => \N__19957\,
            I => \N__19936\
        );

    \I__2363\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19936\
        );

    \I__2362\ : Odrv12
    port map (
            O => \N__19949\,
            I => \r_Bit_Index_2\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__19946\,
            I => \r_Bit_Index_2\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__19941\,
            I => \r_Bit_Index_2\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__19936\,
            I => \r_Bit_Index_2\
        );

    \I__2358\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19922\
        );

    \I__2357\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19919\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__19925\,
            I => \N__19914\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__19922\,
            I => \N__19910\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19907\
        );

    \I__2353\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19904\
        );

    \I__2352\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19901\
        );

    \I__2351\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19896\
        );

    \I__2350\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19896\
        );

    \I__2349\ : Span12Mux_v
    port map (
            O => \N__19910\,
            I => \N__19893\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__19907\,
            I => \N__19890\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19885\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19885\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__19896\,
            I => \N__19882\
        );

    \I__2344\ : Odrv12
    port map (
            O => \N__19893\,
            I => \r_Bit_Index_1_adj_2438\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__19890\,
            I => \r_Bit_Index_1_adj_2438\
        );

    \I__2342\ : Odrv12
    port map (
            O => \N__19885\,
            I => \r_Bit_Index_1_adj_2438\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__19882\,
            I => \r_Bit_Index_1_adj_2438\
        );

    \I__2340\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19869\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__19872\,
            I => \N__19866\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__19869\,
            I => \N__19860\
        );

    \I__2337\ : InMux
    port map (
            O => \N__19866\,
            I => \N__19855\
        );

    \I__2336\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19855\
        );

    \I__2335\ : InMux
    port map (
            O => \N__19864\,
            I => \N__19852\
        );

    \I__2334\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19849\
        );

    \I__2333\ : Span4Mux_h
    port map (
            O => \N__19860\,
            I => \N__19846\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__19855\,
            I => \N__19843\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__19852\,
            I => \r_Clock_Count_7\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__19849\,
            I => \r_Clock_Count_7\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__19846\,
            I => \r_Clock_Count_7\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__19843\,
            I => \r_Clock_Count_7\
        );

    \I__2327\ : InMux
    port map (
            O => \N__19834\,
            I => \N__19831\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__19831\,
            I => \N__19828\
        );

    \I__2325\ : Span4Mux_s3_h
    port map (
            O => \N__19828\,
            I => \N__19821\
        );

    \I__2324\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19816\
        );

    \I__2323\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19816\
        );

    \I__2322\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19811\
        );

    \I__2321\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19811\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__19821\,
            I => \r_Clock_Count_6\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__19816\,
            I => \r_Clock_Count_6\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__19811\,
            I => \r_Clock_Count_6\
        );

    \I__2317\ : InMux
    port map (
            O => \N__19804\,
            I => \N__19797\
        );

    \I__2316\ : InMux
    port map (
            O => \N__19803\,
            I => \N__19797\
        );

    \I__2315\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19794\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__19797\,
            I => \N__19787\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__19794\,
            I => \N__19787\
        );

    \I__2312\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19782\
        );

    \I__2311\ : InMux
    port map (
            O => \N__19792\,
            I => \N__19782\
        );

    \I__2310\ : Span4Mux_h
    port map (
            O => \N__19787\,
            I => \N__19779\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__19782\,
            I => \r_Clock_Count_8\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__19779\,
            I => \r_Clock_Count_8\
        );

    \I__2307\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19771\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__2305\ : Span4Mux_s3_h
    port map (
            O => \N__19768\,
            I => \N__19764\
        );

    \I__2304\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19761\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__19764\,
            I => n9937
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__19761\,
            I => n9937
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__19756\,
            I => \c0.tx.n15683_cascade_\
        );

    \I__2300\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19749\
        );

    \I__2299\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19745\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__19749\,
            I => \N__19742\
        );

    \I__2297\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19739\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__19745\,
            I => \c0.tx.n14082\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__19742\,
            I => \c0.tx.n14082\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__19739\,
            I => \c0.tx.n14082\
        );

    \I__2293\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__19729\,
            I => \N__19726\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__19726\,
            I => n17573
        );

    \I__2290\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19718\
        );

    \I__2289\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19715\
        );

    \I__2288\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19712\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__19718\,
            I => \N__19709\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19706\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__19712\,
            I => \r_Clock_Count_4\
        );

    \I__2284\ : Odrv12
    port map (
            O => \N__19709\,
            I => \r_Clock_Count_4\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__19706\,
            I => \r_Clock_Count_4\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__19699\,
            I => \c0.n12993_cascade_\
        );

    \I__2281\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19693\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__19693\,
            I => \N__19690\
        );

    \I__2279\ : Span12Mux_v
    port map (
            O => \N__19690\,
            I => \N__19687\
        );

    \I__2278\ : Odrv12
    port map (
            O => \N__19687\,
            I => n16856
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__19684\,
            I => \N__19681\
        );

    \I__2276\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19673\
        );

    \I__2275\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19673\
        );

    \I__2274\ : InMux
    port map (
            O => \N__19679\,
            I => \N__19669\
        );

    \I__2273\ : InMux
    port map (
            O => \N__19678\,
            I => \N__19666\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__19673\,
            I => \N__19663\
        );

    \I__2271\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19660\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__19669\,
            I => \N__19656\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__19666\,
            I => \N__19649\
        );

    \I__2268\ : Span4Mux_s2_h
    port map (
            O => \N__19663\,
            I => \N__19649\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__19660\,
            I => \N__19649\
        );

    \I__2266\ : InMux
    port map (
            O => \N__19659\,
            I => \N__19646\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__19656\,
            I => \N__19643\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__19649\,
            I => \N__19640\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__19646\,
            I => \r_Clock_Count_6_adj_2431\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__19643\,
            I => \r_Clock_Count_6_adj_2431\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__19640\,
            I => \r_Clock_Count_6_adj_2431\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__19633\,
            I => \n16893_cascade_\
        );

    \I__2259\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19627\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__19627\,
            I => n5
        );

    \I__2257\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19621\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19618\
        );

    \I__2255\ : Span4Mux_h
    port map (
            O => \N__19618\,
            I => \N__19615\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__19615\,
            I => n17636
        );

    \I__2253\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19603\
        );

    \I__2252\ : InMux
    port map (
            O => \N__19611\,
            I => \N__19603\
        );

    \I__2251\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19603\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__19603\,
            I => data_in_2_4
        );

    \I__2249\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19592\
        );

    \I__2248\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19592\
        );

    \I__2247\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19587\
        );

    \I__2246\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19587\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__19592\,
            I => data_in_1_4
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__19587\,
            I => data_in_1_4
        );

    \I__2243\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19579\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__19579\,
            I => \N__19576\
        );

    \I__2241\ : Span4Mux_h
    port map (
            O => \N__19576\,
            I => \N__19573\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__19573\,
            I => n17567
        );

    \I__2239\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19566\
        );

    \I__2238\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19563\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__19566\,
            I => \N__19559\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__19563\,
            I => \N__19556\
        );

    \I__2235\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19553\
        );

    \I__2234\ : Span4Mux_s3_h
    port map (
            O => \N__19559\,
            I => \N__19548\
        );

    \I__2233\ : Span4Mux_s3_h
    port map (
            O => \N__19556\,
            I => \N__19548\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__19553\,
            I => \r_Clock_Count_4_adj_2450\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__19548\,
            I => \r_Clock_Count_4_adj_2450\
        );

    \I__2230\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19537\
        );

    \I__2229\ : InMux
    port map (
            O => \N__19542\,
            I => \N__19532\
        );

    \I__2228\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19532\
        );

    \I__2227\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19529\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__19537\,
            I => data_in_2_3
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__19532\,
            I => data_in_2_3
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__19529\,
            I => data_in_2_3
        );

    \I__2223\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19519\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__19519\,
            I => \N__19516\
        );

    \I__2221\ : Odrv12
    port map (
            O => \N__19516\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_29\
        );

    \I__2220\ : InMux
    port map (
            O => \N__19513\,
            I => \c0.n15650\
        );

    \I__2219\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19507\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__19507\,
            I => \N__19504\
        );

    \I__2217\ : Sp12to4
    port map (
            O => \N__19504\,
            I => \N__19501\
        );

    \I__2216\ : Odrv12
    port map (
            O => \N__19501\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_30\
        );

    \I__2215\ : InMux
    port map (
            O => \N__19498\,
            I => \c0.n15651\
        );

    \I__2214\ : InMux
    port map (
            O => \N__19495\,
            I => \c0.n15652\
        );

    \I__2213\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19489\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19486\
        );

    \I__2211\ : Span4Mux_s2_h
    port map (
            O => \N__19486\,
            I => \N__19483\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__19483\,
            I => \N__19480\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__19480\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_31\
        );

    \I__2208\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19472\
        );

    \I__2207\ : InMux
    port map (
            O => \N__19476\,
            I => \N__19469\
        );

    \I__2206\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19466\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__19472\,
            I => data_in_0_6
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__19469\,
            I => data_in_0_6
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__19466\,
            I => data_in_0_6
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__19459\,
            I => \c0.n17274_cascade_\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__19456\,
            I => \N__19433\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__19455\,
            I => \N__19430\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__19454\,
            I => \N__19427\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__19453\,
            I => \N__19424\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__19452\,
            I => \N__19421\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__19451\,
            I => \N__19417\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__19450\,
            I => \N__19414\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__19449\,
            I => \N__19410\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__19448\,
            I => \N__19407\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__19447\,
            I => \N__19404\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__19446\,
            I => \N__19399\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__19445\,
            I => \N__19395\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__19444\,
            I => \N__19391\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__19443\,
            I => \N__19387\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__19442\,
            I => \N__19384\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__19441\,
            I => \N__19380\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__19440\,
            I => \N__19376\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__19439\,
            I => \N__19372\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__19438\,
            I => \N__19368\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__19437\,
            I => \N__19365\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__19436\,
            I => \N__19362\
        );

    \I__2180\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19355\
        );

    \I__2179\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19355\
        );

    \I__2178\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19355\
        );

    \I__2177\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19344\
        );

    \I__2176\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19344\
        );

    \I__2175\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19344\
        );

    \I__2174\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19344\
        );

    \I__2173\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19344\
        );

    \I__2172\ : InMux
    port map (
            O => \N__19413\,
            I => \N__19333\
        );

    \I__2171\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19333\
        );

    \I__2170\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19333\
        );

    \I__2169\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19333\
        );

    \I__2168\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19333\
        );

    \I__2167\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19316\
        );

    \I__2166\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19316\
        );

    \I__2165\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19316\
        );

    \I__2164\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19316\
        );

    \I__2163\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19316\
        );

    \I__2162\ : InMux
    port map (
            O => \N__19391\,
            I => \N__19316\
        );

    \I__2161\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19316\
        );

    \I__2160\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19316\
        );

    \I__2159\ : InMux
    port map (
            O => \N__19384\,
            I => \N__19299\
        );

    \I__2158\ : InMux
    port map (
            O => \N__19383\,
            I => \N__19299\
        );

    \I__2157\ : InMux
    port map (
            O => \N__19380\,
            I => \N__19299\
        );

    \I__2156\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19299\
        );

    \I__2155\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19299\
        );

    \I__2154\ : InMux
    port map (
            O => \N__19375\,
            I => \N__19299\
        );

    \I__2153\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19299\
        );

    \I__2152\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19299\
        );

    \I__2151\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19292\
        );

    \I__2150\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19292\
        );

    \I__2149\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19292\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__19355\,
            I => \N__19287\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__19344\,
            I => \N__19287\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__19333\,
            I => \N__19280\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19280\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__19299\,
            I => \N__19280\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__19292\,
            I => \c0.n17889\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__19287\,
            I => \c0.n17889\
        );

    \I__2141\ : Odrv12
    port map (
            O => \N__19280\,
            I => \c0.n17889\
        );

    \I__2140\ : InMux
    port map (
            O => \N__19273\,
            I => \N__19268\
        );

    \I__2139\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19265\
        );

    \I__2138\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19262\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__19268\,
            I => \N__19259\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__19265\,
            I => data_in_3_1
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__19262\,
            I => data_in_3_1
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__19259\,
            I => data_in_3_1
        );

    \I__2133\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19247\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__19251\,
            I => \N__19244\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__19250\,
            I => \N__19241\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__19247\,
            I => \N__19238\
        );

    \I__2129\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19233\
        );

    \I__2128\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19233\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__19238\,
            I => data_in_2_1
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__19233\,
            I => data_in_2_1
        );

    \I__2125\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19225\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__19225\,
            I => \N__19222\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__19222\,
            I => \N__19219\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__19219\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_20\
        );

    \I__2121\ : InMux
    port map (
            O => \N__19216\,
            I => \c0.n15641\
        );

    \I__2120\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19210\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__19210\,
            I => \N__19207\
        );

    \I__2118\ : Span4Mux_h
    port map (
            O => \N__19207\,
            I => \N__19204\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__19204\,
            I => \N__19201\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__19201\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_21\
        );

    \I__2115\ : InMux
    port map (
            O => \N__19198\,
            I => \c0.n15642\
        );

    \I__2114\ : InMux
    port map (
            O => \N__19195\,
            I => \N__19192\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__19192\,
            I => \N__19189\
        );

    \I__2112\ : Span4Mux_s3_h
    port map (
            O => \N__19189\,
            I => \N__19186\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__19186\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_22\
        );

    \I__2110\ : InMux
    port map (
            O => \N__19183\,
            I => \c0.n15643\
        );

    \I__2109\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19177\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__19177\,
            I => \N__19174\
        );

    \I__2107\ : Span4Mux_s1_h
    port map (
            O => \N__19174\,
            I => \N__19171\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__19171\,
            I => \N__19168\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__19168\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_23\
        );

    \I__2104\ : InMux
    port map (
            O => \N__19165\,
            I => \c0.n15644\
        );

    \I__2103\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19159\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__19159\,
            I => \N__19156\
        );

    \I__2101\ : Odrv12
    port map (
            O => \N__19156\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_24\
        );

    \I__2100\ : InMux
    port map (
            O => \N__19153\,
            I => \bfn_4_25_0_\
        );

    \I__2099\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19147\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__19147\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_25\
        );

    \I__2097\ : InMux
    port map (
            O => \N__19144\,
            I => \c0.n15646\
        );

    \I__2096\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19138\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__19138\,
            I => \N__19135\
        );

    \I__2094\ : Span4Mux_s3_h
    port map (
            O => \N__19135\,
            I => \N__19132\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__19132\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_26\
        );

    \I__2092\ : InMux
    port map (
            O => \N__19129\,
            I => \c0.n15647\
        );

    \I__2091\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19123\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__19123\,
            I => \N__19120\
        );

    \I__2089\ : Span4Mux_s3_h
    port map (
            O => \N__19120\,
            I => \N__19117\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__19117\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_27\
        );

    \I__2087\ : InMux
    port map (
            O => \N__19114\,
            I => \c0.n15648\
        );

    \I__2086\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19108\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__2084\ : Sp12to4
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__2083\ : Odrv12
    port map (
            O => \N__19102\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_28\
        );

    \I__2082\ : InMux
    port map (
            O => \N__19099\,
            I => \c0.n15649\
        );

    \I__2081\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__19093\,
            I => \N__19090\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__19090\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_12\
        );

    \I__2078\ : InMux
    port map (
            O => \N__19087\,
            I => \c0.n15633\
        );

    \I__2077\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19081\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__19081\,
            I => \N__19078\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__19078\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_13\
        );

    \I__2074\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19072\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__19072\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_13\
        );

    \I__2072\ : InMux
    port map (
            O => \N__19069\,
            I => \c0.n15634\
        );

    \I__2071\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19063\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__19063\,
            I => \N__19060\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__19060\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_14\
        );

    \I__2068\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19054\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__19054\,
            I => \N__19051\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__19051\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_14\
        );

    \I__2065\ : InMux
    port map (
            O => \N__19048\,
            I => \c0.n15635\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19042\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__19042\,
            I => \N__19039\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__19039\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_15\
        );

    \I__2061\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19033\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__19033\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_15\
        );

    \I__2059\ : InMux
    port map (
            O => \N__19030\,
            I => \c0.n15636\
        );

    \I__2058\ : InMux
    port map (
            O => \N__19027\,
            I => \bfn_4_24_0_\
        );

    \I__2057\ : InMux
    port map (
            O => \N__19024\,
            I => \c0.n15638\
        );

    \I__2056\ : InMux
    port map (
            O => \N__19021\,
            I => \c0.n15639\
        );

    \I__2055\ : InMux
    port map (
            O => \N__19018\,
            I => \N__19015\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__19015\,
            I => \N__19012\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__19012\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_19\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19009\,
            I => \c0.n15640\
        );

    \I__2051\ : InMux
    port map (
            O => \N__19006\,
            I => \c0.n15624\
        );

    \I__2050\ : InMux
    port map (
            O => \N__19003\,
            I => \N__19000\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__19000\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_4\
        );

    \I__2048\ : InMux
    port map (
            O => \N__18997\,
            I => \c0.n15625\
        );

    \I__2047\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18991\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__18991\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_5\
        );

    \I__2045\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18985\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__18985\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_5\
        );

    \I__2043\ : InMux
    port map (
            O => \N__18982\,
            I => \c0.n15626\
        );

    \I__2042\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18976\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__18976\,
            I => \N__18973\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__18973\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_6\
        );

    \I__2039\ : InMux
    port map (
            O => \N__18970\,
            I => \c0.n15627\
        );

    \I__2038\ : InMux
    port map (
            O => \N__18967\,
            I => \c0.n15628\
        );

    \I__2037\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18961\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18958\
        );

    \I__2035\ : Odrv12
    port map (
            O => \N__18958\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_8\
        );

    \I__2034\ : InMux
    port map (
            O => \N__18955\,
            I => \bfn_4_23_0_\
        );

    \I__2033\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18949\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__18949\,
            I => \N__18946\
        );

    \I__2031\ : Span4Mux_s3_h
    port map (
            O => \N__18946\,
            I => \N__18943\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__18943\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_9\
        );

    \I__2029\ : InMux
    port map (
            O => \N__18940\,
            I => \c0.n15630\
        );

    \I__2028\ : InMux
    port map (
            O => \N__18937\,
            I => \c0.n15631\
        );

    \I__2027\ : InMux
    port map (
            O => \N__18934\,
            I => \c0.n15632\
        );

    \I__2026\ : SRMux
    port map (
            O => \N__18931\,
            I => \N__18928\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__18928\,
            I => \N__18925\
        );

    \I__2024\ : Span4Mux_h
    port map (
            O => \N__18925\,
            I => \N__18922\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__18922\,
            I => \c0.n3_adj_2259\
        );

    \I__2022\ : InMux
    port map (
            O => \N__18919\,
            I => \N__18916\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__18916\,
            I => \c0.n10_adj_2329\
        );

    \I__2020\ : InMux
    port map (
            O => \N__18913\,
            I => \N__18910\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__18910\,
            I => \c0.n16895\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__18907\,
            I => \c0.n16895_cascade_\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__18904\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_1_cascade_\
        );

    \I__2016\ : SRMux
    port map (
            O => \N__18901\,
            I => \N__18898\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18895\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__18895\,
            I => \N__18892\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__18892\,
            I => \c0.n3_adj_2260\
        );

    \I__2012\ : InMux
    port map (
            O => \N__18889\,
            I => \bfn_4_22_0_\
        );

    \I__2011\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18883\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__18883\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_1\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__18880\,
            I => \N__18877\
        );

    \I__2008\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18874\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__18874\,
            I => \N__18871\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__18871\,
            I => \N__18868\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__18868\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_1\
        );

    \I__2004\ : InMux
    port map (
            O => \N__18865\,
            I => \c0.n15622\
        );

    \I__2003\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18859\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__18859\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_2\
        );

    \I__2001\ : InMux
    port map (
            O => \N__18856\,
            I => \N__18853\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__18853\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_2\
        );

    \I__1999\ : InMux
    port map (
            O => \N__18850\,
            I => \c0.n15623\
        );

    \I__1998\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18844\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__18844\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_3\
        );

    \I__1996\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18838\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__18838\,
            I => \N__18835\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__18835\,
            I => \c0.FRAME_MATCHER_i_31_N_1280_3\
        );

    \I__1993\ : SRMux
    port map (
            O => \N__18832\,
            I => \N__18829\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__18829\,
            I => \N__18826\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__18826\,
            I => \c0.n3_adj_2217\
        );

    \I__1990\ : SRMux
    port map (
            O => \N__18823\,
            I => \N__18820\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__18820\,
            I => \c0.n3_adj_2215\
        );

    \I__1988\ : SRMux
    port map (
            O => \N__18817\,
            I => \N__18814\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__18814\,
            I => \N__18811\
        );

    \I__1986\ : Span4Mux_s3_h
    port map (
            O => \N__18811\,
            I => \N__18808\
        );

    \I__1985\ : Span4Mux_h
    port map (
            O => \N__18808\,
            I => \N__18805\
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__18805\,
            I => \c0.n3_adj_2210\
        );

    \I__1983\ : SRMux
    port map (
            O => \N__18802\,
            I => \N__18799\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__18799\,
            I => \N__18796\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__18796\,
            I => \N__18793\
        );

    \I__1980\ : Span4Mux_s0_h
    port map (
            O => \N__18793\,
            I => \N__18790\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__18790\,
            I => \c0.n3_adj_2249\
        );

    \I__1978\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18784\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__18784\,
            I => \c0.n9393\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__18781\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_2_cascade_\
        );

    \I__1975\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__18775\,
            I => n16857
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__18772\,
            I => \N__18766\
        );

    \I__1972\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18763\
        );

    \I__1971\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18758\
        );

    \I__1970\ : InMux
    port map (
            O => \N__18769\,
            I => \N__18758\
        );

    \I__1969\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18753\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__18763\,
            I => \N__18748\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__18758\,
            I => \N__18748\
        );

    \I__1966\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18744\
        );

    \I__1965\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18741\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__18753\,
            I => \N__18736\
        );

    \I__1963\ : Span4Mux_s1_v
    port map (
            O => \N__18748\,
            I => \N__18736\
        );

    \I__1962\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18733\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__18744\,
            I => \r_Clock_Count_5_adj_2432\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__18741\,
            I => \r_Clock_Count_5_adj_2432\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__18736\,
            I => \r_Clock_Count_5_adj_2432\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__18733\,
            I => \r_Clock_Count_5_adj_2432\
        );

    \I__1957\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18721\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__18721\,
            I => n16858
        );

    \I__1955\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18714\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__18717\,
            I => \N__18710\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__18714\,
            I => \N__18707\
        );

    \I__1952\ : InMux
    port map (
            O => \N__18713\,
            I => \N__18704\
        );

    \I__1951\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18701\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__18707\,
            I => \r_Clock_Count_3_adj_2434\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__18704\,
            I => \r_Clock_Count_3_adj_2434\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__18701\,
            I => \r_Clock_Count_3_adj_2434\
        );

    \I__1947\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18691\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__18691\,
            I => \N__18688\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__18688\,
            I => n9406
        );

    \I__1944\ : InMux
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__18679\,
            I => n17461
        );

    \I__1941\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18672\
        );

    \I__1940\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18668\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__18672\,
            I => \N__18665\
        );

    \I__1938\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18662\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__18668\,
            I => \r_Clock_Count_1\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__18665\,
            I => \r_Clock_Count_1\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__18662\,
            I => \r_Clock_Count_1\
        );

    \I__1934\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18652\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__18652\,
            I => \N__18649\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__18649\,
            I => \N__18646\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__18646\,
            I => n17601
        );

    \I__1930\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18640\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__18640\,
            I => \N__18637\
        );

    \I__1928\ : Span4Mux_h
    port map (
            O => \N__18637\,
            I => \N__18634\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__18634\,
            I => n17602
        );

    \I__1926\ : InMux
    port map (
            O => \N__18631\,
            I => \N__18627\
        );

    \I__1925\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18623\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__18627\,
            I => \N__18620\
        );

    \I__1923\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18617\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__18623\,
            I => \r_Clock_Count_4_adj_2433\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__18620\,
            I => \r_Clock_Count_4_adj_2433\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__18617\,
            I => \r_Clock_Count_4_adj_2433\
        );

    \I__1919\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18607\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__18607\,
            I => \c0.rx.n6\
        );

    \I__1917\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18601\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__18601\,
            I => \N__18598\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__18598\,
            I => n16853
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__18595\,
            I => \N__18592\
        );

    \I__1913\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18589\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__18589\,
            I => \N__18584\
        );

    \I__1911\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18579\
        );

    \I__1910\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18579\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__18584\,
            I => \r_Clock_Count_1_adj_2436\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__18579\,
            I => \r_Clock_Count_1_adj_2436\
        );

    \I__1907\ : InMux
    port map (
            O => \N__18574\,
            I => \N__18569\
        );

    \I__1906\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18564\
        );

    \I__1905\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18564\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__18569\,
            I => \N__18561\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__18564\,
            I => \N__18558\
        );

    \I__1902\ : Odrv12
    port map (
            O => \N__18561\,
            I => n4_adj_2411
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__18558\,
            I => n4_adj_2411
        );

    \I__1900\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18547\
        );

    \I__1899\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18544\
        );

    \I__1898\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18539\
        );

    \I__1897\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18539\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18534\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__18544\,
            I => \N__18534\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__18539\,
            I => \N__18531\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__18534\,
            I => \N__18528\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__18531\,
            I => \N__18525\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__18528\,
            I => n17260
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__18525\,
            I => n17260
        );

    \I__1889\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18516\
        );

    \I__1888\ : InMux
    port map (
            O => \N__18519\,
            I => \N__18513\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18508\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__18513\,
            I => \N__18508\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__18508\,
            I => n10425
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__18505\,
            I => \n7866_cascade_\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__18502\,
            I => \n10425_cascade_\
        );

    \I__1882\ : InMux
    port map (
            O => \N__18499\,
            I => \N__18494\
        );

    \I__1881\ : InMux
    port map (
            O => \N__18498\,
            I => \N__18489\
        );

    \I__1880\ : InMux
    port map (
            O => \N__18497\,
            I => \N__18489\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__18494\,
            I => \N__18486\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__18489\,
            I => n12
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__18486\,
            I => n12
        );

    \I__1876\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18478\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__18478\,
            I => n13276
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__18475\,
            I => \n10_adj_2415_cascade_\
        );

    \I__1873\ : InMux
    port map (
            O => \N__18472\,
            I => \N__18467\
        );

    \I__1872\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18464\
        );

    \I__1871\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18461\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__18467\,
            I => n15701
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__18464\,
            I => n15701
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__18461\,
            I => n15701
        );

    \I__1867\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18451\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__18451\,
            I => \N__18446\
        );

    \I__1865\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18443\
        );

    \I__1864\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18440\
        );

    \I__1863\ : Span4Mux_s3_h
    port map (
            O => \N__18446\,
            I => \N__18437\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__18443\,
            I => \N__18432\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__18440\,
            I => \N__18432\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__18437\,
            I => n16844
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__18432\,
            I => n16844
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__18427\,
            I => \n9472_cascade_\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__18424\,
            I => \c0.rx.n10086_cascade_\
        );

    \I__1856\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18417\
        );

    \I__1855\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18414\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__18417\,
            I => \N__18409\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__18414\,
            I => \N__18406\
        );

    \I__1852\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18403\
        );

    \I__1851\ : InMux
    port map (
            O => \N__18412\,
            I => \N__18400\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__18409\,
            I => \N__18397\
        );

    \I__1849\ : Span4Mux_h
    port map (
            O => \N__18406\,
            I => \N__18392\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__18403\,
            I => \N__18392\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__18400\,
            I => \N__18389\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__18397\,
            I => \c0.rx.r_SM_Main_2_N_2090_2\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__18392\,
            I => \c0.rx.r_SM_Main_2_N_2090_2\
        );

    \I__1844\ : Odrv12
    port map (
            O => \N__18389\,
            I => \c0.rx.r_SM_Main_2_N_2090_2\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__18382\,
            I => \n14060_cascade_\
        );

    \I__1842\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18375\
        );

    \I__1841\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18372\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__18375\,
            I => data_in_0_7
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__18372\,
            I => data_in_0_7
        );

    \I__1838\ : InMux
    port map (
            O => \N__18367\,
            I => \N__18362\
        );

    \I__1837\ : InMux
    port map (
            O => \N__18366\,
            I => \N__18359\
        );

    \I__1836\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18356\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__18362\,
            I => data_in_1_5
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__18359\,
            I => data_in_1_5
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__18356\,
            I => data_in_1_5
        );

    \I__1832\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18343\
        );

    \I__1831\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18343\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__18343\,
            I => data_in_0_4
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__18340\,
            I => \c0.n17172_cascade_\
        );

    \I__1828\ : SRMux
    port map (
            O => \N__18337\,
            I => \N__18334\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__18334\,
            I => \N__18331\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__18331\,
            I => \c0.n3_adj_2242\
        );

    \I__1825\ : SRMux
    port map (
            O => \N__18328\,
            I => \N__18325\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__18325\,
            I => \c0.n3_adj_2243\
        );

    \I__1823\ : SRMux
    port map (
            O => \N__18322\,
            I => \N__18319\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__18319\,
            I => \N__18316\
        );

    \I__1821\ : Span4Mux_s3_h
    port map (
            O => \N__18316\,
            I => \N__18313\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__18313\,
            I => \c0.n3_adj_2244\
        );

    \I__1819\ : SRMux
    port map (
            O => \N__18310\,
            I => \N__18307\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__18307\,
            I => \N__18304\
        );

    \I__1817\ : Span4Mux_s3_h
    port map (
            O => \N__18304\,
            I => \N__18301\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__18301\,
            I => \c0.n3_adj_2256\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__18298\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_4_cascade_\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__18295\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_3_cascade_\
        );

    \I__1813\ : SRMux
    port map (
            O => \N__18292\,
            I => \N__18289\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__18289\,
            I => \N__18286\
        );

    \I__1811\ : Span4Mux_s2_h
    port map (
            O => \N__18286\,
            I => \N__18283\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__18283\,
            I => \c0.n3_adj_2258\
        );

    \I__1809\ : SRMux
    port map (
            O => \N__18280\,
            I => \N__18277\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__18277\,
            I => \N__18274\
        );

    \I__1807\ : Span4Mux_s3_h
    port map (
            O => \N__18274\,
            I => \N__18271\
        );

    \I__1806\ : Odrv4
    port map (
            O => \N__18271\,
            I => \c0.n16379\
        );

    \I__1805\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18265\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__18265\,
            I => n1651
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__18262\,
            I => \n6_cascade_\
        );

    \I__1802\ : InMux
    port map (
            O => \N__18259\,
            I => \N__18256\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__18256\,
            I => n4
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__18253\,
            I => \n8_adj_2459_cascade_\
        );

    \I__1799\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18247\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__18247\,
            I => \FRAME_MATCHER_state_31_N_1440_1\
        );

    \I__1797\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18241\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__18241\,
            I => n3_adj_2408
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__18238\,
            I => \c0.FRAME_MATCHER_i_31_N_1312_5_cascade_\
        );

    \I__1794\ : InMux
    port map (
            O => \N__18235\,
            I => \N__18232\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__18232\,
            I => \N__18229\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__18229\,
            I => n16854
        );

    \I__1791\ : InMux
    port map (
            O => \N__18226\,
            I => \c0.rx.n15671\
        );

    \I__1790\ : InMux
    port map (
            O => \N__18223\,
            I => \c0.rx.n15672\
        );

    \I__1789\ : InMux
    port map (
            O => \N__18220\,
            I => \c0.rx.n15673\
        );

    \I__1788\ : InMux
    port map (
            O => \N__18217\,
            I => \N__18214\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__18214\,
            I => \N__18206\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18213\,
            I => \N__18203\
        );

    \I__1785\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18200\
        );

    \I__1784\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18197\
        );

    \I__1783\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18192\
        );

    \I__1782\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18192\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__18206\,
            I => \r_Clock_Count_7_adj_2430\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__18203\,
            I => \r_Clock_Count_7_adj_2430\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__18200\,
            I => \r_Clock_Count_7_adj_2430\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__18197\,
            I => \r_Clock_Count_7_adj_2430\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__18192\,
            I => \r_Clock_Count_7_adj_2430\
        );

    \I__1776\ : InMux
    port map (
            O => \N__18181\,
            I => \N__18167\
        );

    \I__1775\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18167\
        );

    \I__1774\ : InMux
    port map (
            O => \N__18179\,
            I => \N__18167\
        );

    \I__1773\ : InMux
    port map (
            O => \N__18178\,
            I => \N__18156\
        );

    \I__1772\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18156\
        );

    \I__1771\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18156\
        );

    \I__1770\ : InMux
    port map (
            O => \N__18175\,
            I => \N__18156\
        );

    \I__1769\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18156\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__18167\,
            I => n16852
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__18156\,
            I => n16852
        );

    \I__1766\ : InMux
    port map (
            O => \N__18151\,
            I => \c0.rx.n15674\
        );

    \I__1765\ : InMux
    port map (
            O => \N__18148\,
            I => \N__18145\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__18145\,
            I => n16855
        );

    \I__1763\ : InMux
    port map (
            O => \N__18142\,
            I => \N__18137\
        );

    \I__1762\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18132\
        );

    \I__1761\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18132\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__18137\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__18132\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__1758\ : SRMux
    port map (
            O => \N__18127\,
            I => \N__18124\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__18124\,
            I => \c0.n16349\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__18121\,
            I => \n1651_cascade_\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__18118\,
            I => \c0.rx.r_SM_Main_2_N_2096_0_cascade_\
        );

    \I__1754\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18112\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__18112\,
            I => n6_adj_2461
        );

    \I__1752\ : InMux
    port map (
            O => \N__18109\,
            I => \N__18106\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__18106\,
            I => n17641
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__18103\,
            I => \n17144_cascade_\
        );

    \I__1749\ : InMux
    port map (
            O => \N__18100\,
            I => \N__18088\
        );

    \I__1748\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18088\
        );

    \I__1747\ : InMux
    port map (
            O => \N__18098\,
            I => \N__18088\
        );

    \I__1746\ : InMux
    port map (
            O => \N__18097\,
            I => \N__18081\
        );

    \I__1745\ : InMux
    port map (
            O => \N__18096\,
            I => \N__18081\
        );

    \I__1744\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18081\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__18088\,
            I => n16828
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__18081\,
            I => n16828
        );

    \I__1741\ : InMux
    port map (
            O => \N__18076\,
            I => \bfn_2_32_0_\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18073\,
            I => \c0.rx.n15668\
        );

    \I__1739\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18066\
        );

    \I__1738\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18062\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__18066\,
            I => \N__18059\
        );

    \I__1736\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18056\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__18062\,
            I => \r_Clock_Count_2_adj_2435\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__18059\,
            I => \r_Clock_Count_2_adj_2435\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__18056\,
            I => \r_Clock_Count_2_adj_2435\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18046\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__18046\,
            I => \N__18043\
        );

    \I__1730\ : Odrv4
    port map (
            O => \N__18043\,
            I => n16860
        );

    \I__1729\ : InMux
    port map (
            O => \N__18040\,
            I => \c0.rx.n15669\
        );

    \I__1728\ : InMux
    port map (
            O => \N__18037\,
            I => \c0.rx.n15670\
        );

    \I__1727\ : InMux
    port map (
            O => \N__18034\,
            I => \N__18031\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__18031\,
            I => n17494
        );

    \I__1725\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18025\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__18025\,
            I => n17542
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__18022\,
            I => \N__18019\
        );

    \I__1722\ : InMux
    port map (
            O => \N__18019\,
            I => \N__18016\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__18016\,
            I => n17484
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__18013\,
            I => \n17_adj_2416_cascade_\
        );

    \I__1719\ : InMux
    port map (
            O => \N__18010\,
            I => \N__18005\
        );

    \I__1718\ : InMux
    port map (
            O => \N__18009\,
            I => \N__18000\
        );

    \I__1717\ : InMux
    port map (
            O => \N__18008\,
            I => \N__18000\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__18005\,
            I => \r_Clock_Count_2\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__18000\,
            I => \r_Clock_Count_2\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__17995\,
            I => \N__17990\
        );

    \I__1713\ : InMux
    port map (
            O => \N__17994\,
            I => \N__17987\
        );

    \I__1712\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17982\
        );

    \I__1711\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17982\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__17987\,
            I => \r_Clock_Count_3\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__17982\,
            I => \r_Clock_Count_3\
        );

    \I__1708\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17972\
        );

    \I__1707\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17967\
        );

    \I__1706\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17967\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__17972\,
            I => \r_Clock_Count_0\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__17967\,
            I => \r_Clock_Count_0\
        );

    \I__1703\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17957\
        );

    \I__1702\ : InMux
    port map (
            O => \N__17961\,
            I => \N__17954\
        );

    \I__1701\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17951\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__17957\,
            I => \r_Clock_Count_5\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__17954\,
            I => \r_Clock_Count_5\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__17951\,
            I => \r_Clock_Count_5\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__17944\,
            I => \c0.tx.n10_cascade_\
        );

    \I__1696\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17935\
        );

    \I__1695\ : InMux
    port map (
            O => \N__17940\,
            I => \N__17928\
        );

    \I__1694\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17928\
        );

    \I__1693\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17928\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__17935\,
            I => n16863
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__17928\,
            I => n16863
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__17923\,
            I => \n16863_cascade_\
        );

    \I__1689\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17917\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__17917\,
            I => n9403
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__17914\,
            I => \n17140_cascade_\
        );

    \I__1686\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17899\
        );

    \I__1685\ : InMux
    port map (
            O => \N__17910\,
            I => \N__17899\
        );

    \I__1684\ : InMux
    port map (
            O => \N__17909\,
            I => \N__17899\
        );

    \I__1683\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17892\
        );

    \I__1682\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17892\
        );

    \I__1681\ : InMux
    port map (
            O => \N__17906\,
            I => \N__17892\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__17899\,
            I => n16817
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__17892\,
            I => n16817
        );

    \I__1678\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17882\
        );

    \I__1677\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17877\
        );

    \I__1676\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17877\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__17882\,
            I => n12_adj_2410
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__17877\,
            I => n12_adj_2410
        );

    \I__1673\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17867\
        );

    \I__1672\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17864\
        );

    \I__1671\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17861\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__17867\,
            I => \r_Clock_Count_5_adj_2449\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__17864\,
            I => \r_Clock_Count_5_adj_2449\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__17861\,
            I => \r_Clock_Count_5_adj_2449\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__17854\,
            I => \N__17851\
        );

    \I__1666\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17846\
        );

    \I__1665\ : InMux
    port map (
            O => \N__17850\,
            I => \N__17843\
        );

    \I__1664\ : InMux
    port map (
            O => \N__17849\,
            I => \N__17840\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__17846\,
            I => \r_Clock_Count_1_adj_2453\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__17843\,
            I => \r_Clock_Count_1_adj_2453\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__17840\,
            I => \r_Clock_Count_1_adj_2453\
        );

    \I__1660\ : InMux
    port map (
            O => \N__17833\,
            I => \N__17830\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__17830\,
            I => \c0.tx2.n10\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__17827\,
            I => \N__17824\
        );

    \I__1657\ : InMux
    port map (
            O => \N__17824\,
            I => \N__17820\
        );

    \I__1656\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17817\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__17820\,
            I => n15837
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__17817\,
            I => n15837
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__17812\,
            I => \n15837_cascade_\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__17809\,
            I => \r_SM_Main_2_N_2033_1_cascade_\
        );

    \I__1651\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17799\
        );

    \I__1650\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17796\
        );

    \I__1649\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17789\
        );

    \I__1648\ : InMux
    port map (
            O => \N__17803\,
            I => \N__17789\
        );

    \I__1647\ : InMux
    port map (
            O => \N__17802\,
            I => \N__17789\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__17799\,
            I => \r_Clock_Count_7_adj_2447\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__17796\,
            I => \r_Clock_Count_7_adj_2447\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__17789\,
            I => \r_Clock_Count_7_adj_2447\
        );

    \I__1643\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17773\
        );

    \I__1642\ : InMux
    port map (
            O => \N__17781\,
            I => \N__17773\
        );

    \I__1641\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17766\
        );

    \I__1640\ : InMux
    port map (
            O => \N__17779\,
            I => \N__17766\
        );

    \I__1639\ : InMux
    port map (
            O => \N__17778\,
            I => \N__17766\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__17773\,
            I => \r_Clock_Count_8_adj_2446\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__17766\,
            I => \r_Clock_Count_8_adj_2446\
        );

    \I__1636\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17757\
        );

    \I__1635\ : InMux
    port map (
            O => \N__17760\,
            I => \N__17754\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__17757\,
            I => n9929
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__17754\,
            I => n9929
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__17749\,
            I => \N__17745\
        );

    \I__1631\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17739\
        );

    \I__1630\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17739\
        );

    \I__1629\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17736\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__17739\,
            I => blink_counter_23
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__17736\,
            I => blink_counter_23
        );

    \I__1626\ : InMux
    port map (
            O => \N__17731\,
            I => n15612
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__17728\,
            I => \N__17725\
        );

    \I__1624\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17718\
        );

    \I__1623\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17718\
        );

    \I__1622\ : InMux
    port map (
            O => \N__17723\,
            I => \N__17715\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__17718\,
            I => blink_counter_24
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__17715\,
            I => blink_counter_24
        );

    \I__1619\ : InMux
    port map (
            O => \N__17710\,
            I => \bfn_2_28_0_\
        );

    \I__1618\ : InMux
    port map (
            O => \N__17707\,
            I => n15614
        );

    \I__1617\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17700\
        );

    \I__1616\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17697\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__17700\,
            I => blink_counter_25
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__17697\,
            I => blink_counter_25
        );

    \I__1613\ : InMux
    port map (
            O => \N__17692\,
            I => \N__17689\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__17689\,
            I => n17570
        );

    \I__1611\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17683\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__17683\,
            I => n17629
        );

    \I__1609\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17677\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__17677\,
            I => n17504
        );

    \I__1607\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17669\
        );

    \I__1606\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17664\
        );

    \I__1605\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17664\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__17669\,
            I => \r_Clock_Count_2_adj_2452\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__17664\,
            I => \r_Clock_Count_2_adj_2452\
        );

    \I__1602\ : InMux
    port map (
            O => \N__17659\,
            I => \N__17654\
        );

    \I__1601\ : InMux
    port map (
            O => \N__17658\,
            I => \N__17651\
        );

    \I__1600\ : InMux
    port map (
            O => \N__17657\,
            I => \N__17648\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__17654\,
            I => \r_Clock_Count_3_adj_2451\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__17651\,
            I => \r_Clock_Count_3_adj_2451\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__17648\,
            I => \r_Clock_Count_3_adj_2451\
        );

    \I__1596\ : InMux
    port map (
            O => \N__17641\,
            I => n15603
        );

    \I__1595\ : InMux
    port map (
            O => \N__17638\,
            I => \N__17635\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__17635\,
            I => n11
        );

    \I__1593\ : InMux
    port map (
            O => \N__17632\,
            I => n15604
        );

    \I__1592\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17626\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__17626\,
            I => n10_adj_2420
        );

    \I__1590\ : InMux
    port map (
            O => \N__17623\,
            I => \bfn_2_27_0_\
        );

    \I__1589\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17617\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__17617\,
            I => n9
        );

    \I__1587\ : InMux
    port map (
            O => \N__17614\,
            I => n15606
        );

    \I__1586\ : InMux
    port map (
            O => \N__17611\,
            I => \N__17608\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__17608\,
            I => n8
        );

    \I__1584\ : InMux
    port map (
            O => \N__17605\,
            I => n15607
        );

    \I__1583\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17599\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__17599\,
            I => n7
        );

    \I__1581\ : InMux
    port map (
            O => \N__17596\,
            I => n15608
        );

    \I__1580\ : InMux
    port map (
            O => \N__17593\,
            I => \N__17590\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__17590\,
            I => n6_adj_2421
        );

    \I__1578\ : InMux
    port map (
            O => \N__17587\,
            I => n15609
        );

    \I__1577\ : InMux
    port map (
            O => \N__17584\,
            I => \N__17578\
        );

    \I__1576\ : InMux
    port map (
            O => \N__17583\,
            I => \N__17578\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17574\
        );

    \I__1574\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17571\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__17574\,
            I => blink_counter_21
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__17571\,
            I => blink_counter_21
        );

    \I__1571\ : InMux
    port map (
            O => \N__17566\,
            I => n15610
        );

    \I__1570\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17556\
        );

    \I__1569\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17556\
        );

    \I__1568\ : InMux
    port map (
            O => \N__17561\,
            I => \N__17553\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__17556\,
            I => blink_counter_22
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__17553\,
            I => blink_counter_22
        );

    \I__1565\ : InMux
    port map (
            O => \N__17548\,
            I => n15611
        );

    \I__1564\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17542\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__17542\,
            I => n20
        );

    \I__1562\ : InMux
    port map (
            O => \N__17539\,
            I => n15595
        );

    \I__1561\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17533\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__17533\,
            I => n19
        );

    \I__1559\ : InMux
    port map (
            O => \N__17530\,
            I => n15596
        );

    \I__1558\ : InMux
    port map (
            O => \N__17527\,
            I => \N__17524\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__17524\,
            I => n18
        );

    \I__1556\ : InMux
    port map (
            O => \N__17521\,
            I => \bfn_2_26_0_\
        );

    \I__1555\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17515\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__17515\,
            I => n17_adj_2422
        );

    \I__1553\ : InMux
    port map (
            O => \N__17512\,
            I => n15598
        );

    \I__1552\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17506\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__17506\,
            I => n16
        );

    \I__1550\ : InMux
    port map (
            O => \N__17503\,
            I => n15599
        );

    \I__1549\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17497\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__17497\,
            I => n15
        );

    \I__1547\ : InMux
    port map (
            O => \N__17494\,
            I => n15600
        );

    \I__1546\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17488\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__17488\,
            I => n14_adj_2424
        );

    \I__1544\ : InMux
    port map (
            O => \N__17485\,
            I => n15601
        );

    \I__1543\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17479\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__17479\,
            I => n13
        );

    \I__1541\ : InMux
    port map (
            O => \N__17476\,
            I => n15602
        );

    \I__1540\ : InMux
    port map (
            O => \N__17473\,
            I => \N__17470\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__17470\,
            I => n12_adj_2419
        );

    \I__1538\ : InMux
    port map (
            O => \N__17467\,
            I => \N__17464\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__17464\,
            I => n26
        );

    \I__1536\ : InMux
    port map (
            O => \N__17461\,
            I => \bfn_2_25_0_\
        );

    \I__1535\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17455\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__17455\,
            I => n25
        );

    \I__1533\ : InMux
    port map (
            O => \N__17452\,
            I => n15590
        );

    \I__1532\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17446\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__17446\,
            I => n24
        );

    \I__1530\ : InMux
    port map (
            O => \N__17443\,
            I => n15591
        );

    \I__1529\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17437\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__17437\,
            I => n23
        );

    \I__1527\ : InMux
    port map (
            O => \N__17434\,
            I => n15592
        );

    \I__1526\ : InMux
    port map (
            O => \N__17431\,
            I => \N__17428\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__17428\,
            I => n22
        );

    \I__1524\ : InMux
    port map (
            O => \N__17425\,
            I => n15593
        );

    \I__1523\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17419\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__17419\,
            I => n21
        );

    \I__1521\ : InMux
    port map (
            O => \N__17416\,
            I => n15594
        );

    \I__1520\ : InMux
    port map (
            O => \N__17413\,
            I => \N__17404\
        );

    \I__1519\ : InMux
    port map (
            O => \N__17412\,
            I => \N__17404\
        );

    \I__1518\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17404\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__17404\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__1516\ : SRMux
    port map (
            O => \N__17401\,
            I => \N__17398\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__17398\,
            I => \N__17395\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__17395\,
            I => \c0.n16443\
        );

    \I__1513\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17387\
        );

    \I__1512\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17382\
        );

    \I__1511\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17382\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__17387\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__17382\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__1508\ : SRMux
    port map (
            O => \N__17377\,
            I => \N__17374\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__17374\,
            I => \N__17371\
        );

    \I__1506\ : Span4Mux_s1_h
    port map (
            O => \N__17371\,
            I => \N__17368\
        );

    \I__1505\ : Span4Mux_h
    port map (
            O => \N__17368\,
            I => \N__17365\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__17365\,
            I => \c0.n16447\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__17362\,
            I => \N__17358\
        );

    \I__1502\ : InMux
    port map (
            O => \N__17361\,
            I => \N__17353\
        );

    \I__1501\ : InMux
    port map (
            O => \N__17358\,
            I => \N__17353\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__17353\,
            I => \N__17349\
        );

    \I__1499\ : InMux
    port map (
            O => \N__17352\,
            I => \N__17346\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__17349\,
            I => \N__17343\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__17346\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__17343\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__1495\ : SRMux
    port map (
            O => \N__17338\,
            I => \N__17335\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__17335\,
            I => \c0.n16451\
        );

    \I__1493\ : SRMux
    port map (
            O => \N__17332\,
            I => \N__17329\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__17329\,
            I => \N__17326\
        );

    \I__1491\ : Odrv12
    port map (
            O => \N__17326\,
            I => \c0.n16445\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__17323\,
            I => \c0.rx.r_SM_Main_2_N_2090_2_cascade_\
        );

    \I__1489\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17317\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__17317\,
            I => n17631
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__17314\,
            I => \n16810_cascade_\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__17311\,
            I => \c0.rx.n13452_cascade_\
        );

    \I__1485\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17305\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__17305\,
            I => n16867
        );

    \I__1483\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17296\
        );

    \I__1482\ : InMux
    port map (
            O => \N__17301\,
            I => \N__17296\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__17296\,
            I => n17222
        );

    \I__1480\ : SRMux
    port map (
            O => \N__17293\,
            I => \N__17290\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__17290\,
            I => \N__17287\
        );

    \I__1478\ : Span4Mux_s3_v
    port map (
            O => \N__17287\,
            I => \N__17284\
        );

    \I__1477\ : Span4Mux_s1_h
    port map (
            O => \N__17284\,
            I => \N__17281\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__17281\,
            I => \c0.rx.n16850\
        );

    \I__1475\ : InMux
    port map (
            O => \N__17278\,
            I => \c0.tx.n15662\
        );

    \I__1474\ : InMux
    port map (
            O => \N__17275\,
            I => \c0.tx.n15663\
        );

    \I__1473\ : InMux
    port map (
            O => \N__17272\,
            I => \c0.tx.n15664\
        );

    \I__1472\ : InMux
    port map (
            O => \N__17269\,
            I => \c0.tx.n15665\
        );

    \I__1471\ : InMux
    port map (
            O => \N__17266\,
            I => \c0.tx.n15666\
        );

    \I__1470\ : InMux
    port map (
            O => \N__17263\,
            I => \bfn_1_31_0_\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__17260\,
            I => \n17537_cascade_\
        );

    \I__1468\ : InMux
    port map (
            O => \N__17257\,
            I => \bfn_1_29_0_\
        );

    \I__1467\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17251\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__17251\,
            I => n17640
        );

    \I__1465\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17243\
        );

    \I__1464\ : InMux
    port map (
            O => \N__17247\,
            I => \N__17240\
        );

    \I__1463\ : InMux
    port map (
            O => \N__17246\,
            I => \N__17237\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__17243\,
            I => n16824
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__17240\,
            I => n16824
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__17237\,
            I => n16824
        );

    \I__1459\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17227\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__17227\,
            I => n10_adj_2412
        );

    \I__1457\ : InMux
    port map (
            O => \N__17224\,
            I => \N__17221\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__17221\,
            I => n17458
        );

    \I__1455\ : InMux
    port map (
            O => \N__17218\,
            I => \bfn_1_30_0_\
        );

    \I__1454\ : InMux
    port map (
            O => \N__17215\,
            I => \c0.tx.n15660\
        );

    \I__1453\ : InMux
    port map (
            O => \N__17212\,
            I => \c0.tx.n15661\
        );

    \I__1452\ : InMux
    port map (
            O => \N__17209\,
            I => \N__17206\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__17206\,
            I => n17298
        );

    \I__1450\ : InMux
    port map (
            O => \N__17203\,
            I => \bfn_1_28_0_\
        );

    \I__1449\ : InMux
    port map (
            O => \N__17200\,
            I => \c0.tx2.n15675\
        );

    \I__1448\ : InMux
    port map (
            O => \N__17197\,
            I => \c0.tx2.n15676\
        );

    \I__1447\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17191\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__17191\,
            I => n17457
        );

    \I__1445\ : InMux
    port map (
            O => \N__17188\,
            I => \c0.tx2.n15677\
        );

    \I__1444\ : InMux
    port map (
            O => \N__17185\,
            I => \c0.tx2.n15678\
        );

    \I__1443\ : InMux
    port map (
            O => \N__17182\,
            I => \c0.tx2.n15679\
        );

    \I__1442\ : InMux
    port map (
            O => \N__17179\,
            I => \c0.tx2.n15680\
        );

    \I__1441\ : InMux
    port map (
            O => \N__17176\,
            I => \c0.tx2.n15681\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__17173\,
            I => \n17299_cascade_\
        );

    \I__1439\ : IoInMux
    port map (
            O => \N__17170\,
            I => \N__17167\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__17167\,
            I => \N__17164\
        );

    \I__1437\ : Span4Mux_s1_v
    port map (
            O => \N__17164\,
            I => \N__17161\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__17161\,
            I => \N__17158\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__17158\,
            I => \LED_c\
        );

    \I__1434\ : IoInMux
    port map (
            O => \N__17155\,
            I => \N__17152\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__17152\,
            I => tx2_enable
        );

    \I__1432\ : IoInMux
    port map (
            O => \N__17149\,
            I => \N__17146\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__17146\,
            I => \N__17143\
        );

    \I__1430\ : IoSpan4Mux
    port map (
            O => \N__17143\,
            I => \N__17140\
        );

    \I__1429\ : IoSpan4Mux
    port map (
            O => \N__17140\,
            I => \N__17137\
        );

    \I__1428\ : IoSpan4Mux
    port map (
            O => \N__17137\,
            I => \N__17134\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__17134\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_13_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_29_0_\
        );

    \IN_MUX_bfv_13_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15566,
            carryinitout => \bfn_13_30_0_\
        );

    \IN_MUX_bfv_13_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15574,
            carryinitout => \bfn_13_31_0_\
        );

    \IN_MUX_bfv_13_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15582,
            carryinitout => \bfn_13_32_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15535,
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_13_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15543,
            carryinitout => \bfn_13_27_0_\
        );

    \IN_MUX_bfv_13_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15551,
            carryinitout => \bfn_13_28_0_\
        );

    \IN_MUX_bfv_1_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_28_0_\
        );

    \IN_MUX_bfv_1_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx2.n15682\,
            carryinitout => \bfn_1_29_0_\
        );

    \IN_MUX_bfv_1_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_30_0_\
        );

    \IN_MUX_bfv_1_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n15667\,
            carryinitout => \bfn_1_31_0_\
        );

    \IN_MUX_bfv_2_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_32_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_4_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_22_0_\
        );

    \IN_MUX_bfv_4_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n15629\,
            carryinitout => \bfn_4_23_0_\
        );

    \IN_MUX_bfv_4_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n15637\,
            carryinitout => \bfn_4_24_0_\
        );

    \IN_MUX_bfv_4_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n15645\,
            carryinitout => \bfn_4_25_0_\
        );

    \IN_MUX_bfv_5_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_31_0_\
        );

    \IN_MUX_bfv_5_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n15521\,
            carryinitout => \bfn_5_32_0_\
        );

    \IN_MUX_bfv_6_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_30_0_\
        );

    \IN_MUX_bfv_2_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_25_0_\
        );

    \IN_MUX_bfv_2_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15597,
            carryinitout => \bfn_2_26_0_\
        );

    \IN_MUX_bfv_2_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15605,
            carryinitout => \bfn_2_27_0_\
        );

    \IN_MUX_bfv_2_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15613,
            carryinitout => \bfn_2_28_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17149\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i11_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__34663\,
            in1 => \N__17352\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_state_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50377\,
            ce => 'H',
            sr => \N__17338\
        );

    \c0.FRAME_MATCHER_state_i8_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34655\,
            in2 => \_gnd_net_\,
            in3 => \N__30110\,
            lcout => \c0.FRAME_MATCHER_state_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50378\,
            ce => 'H',
            sr => \N__17332\
        );

    \c0.FRAME_MATCHER_state_i13_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__34660\,
            in1 => \N__17392\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_state_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50380\,
            ce => 'H',
            sr => \N__17377\
        );

    \c0.FRAME_MATCHER_i_i23_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33226\,
            in1 => \N__33004\,
            in2 => \_gnd_net_\,
            in3 => \N__19180\,
            lcout => \c0.FRAME_MATCHER_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50383\,
            ce => 'H',
            sr => \N__20206\
        );

    \c0.FRAME_MATCHER_i_i20_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33257\,
            in1 => \N__32911\,
            in2 => \_gnd_net_\,
            in3 => \N__19228\,
            lcout => \c0.FRAME_MATCHER_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50387\,
            ce => 'H',
            sr => \N__20374\
        );

    \c0.FRAME_MATCHER_i_i22_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33266\,
            in1 => \N__33003\,
            in2 => \_gnd_net_\,
            in3 => \N__19195\,
            lcout => \c0.FRAME_MATCHER_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50393\,
            ce => 'H',
            sr => \N__20332\
        );

    \c0.FRAME_MATCHER_i_i8_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__32999\,
            in1 => \N__33268\,
            in2 => \_gnd_net_\,
            in3 => \N__18964\,
            lcout => \c0.FRAME_MATCHER_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50400\,
            ce => 'H',
            sr => \N__18802\
        );

    \c0.FRAME_MATCHER_i_i26_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33000\,
            in1 => \N__33269\,
            in2 => \_gnd_net_\,
            in3 => \N__19141\,
            lcout => \c0.FRAME_MATCHER_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50406\,
            ce => 'H',
            sr => \N__20302\
        );

    \c0.FRAME_MATCHER_i_i1_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33279\,
            in2 => \N__18880\,
            in3 => \N__33001\,
            lcout => \c0.FRAME_MATCHER_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50413\,
            ce => 'H',
            sr => \N__18901\
        );

    \c0.FRAME_MATCHER_i_i27_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33280\,
            in1 => \N__33002\,
            in2 => \_gnd_net_\,
            in3 => \N__19126\,
            lcout => \c0.FRAME_MATCHER_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50423\,
            ce => 'H',
            sr => \N__20272\
        );

    \c0.tx2.r_Clock_Count__i3_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17194\,
            in1 => \N__31532\,
            in2 => \_gnd_net_\,
            in3 => \N__17659\,
            lcout => \r_Clock_Count_3_adj_2451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i14822_4_lut_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__30779\,
            in1 => \N__30852\,
            in2 => \N__33874\,
            in3 => \N__18412\,
            lcout => n17260,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14861_4_lut_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011000100"
        )
    port map (
            in0 => \N__17563\,
            in1 => \N__17748\,
            in2 => \N__17728\,
            in3 => \N__17584\,
            lcout => OPEN,
            ltout => \n17299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14862_3_lut_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__17704\,
            in1 => \_gnd_net_\,
            in2 => \N__17173\,
            in3 => \N__17209\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i81_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__25602\,
            in1 => \N__31924\,
            in2 => \N__23664\,
            in3 => \N__31137\,
            lcout => \c0.data_in_frame_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15447_2_lut_3_lut_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__30780\,
            in1 => \_gnd_net_\,
            in2 => \N__33875\,
            in3 => \N__30853\,
            lcout => \c0.rx.n16850\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx2_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14860_4_lut_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000100010"
        )
    port map (
            in0 => \N__17583\,
            in1 => \N__17724\,
            in2 => \N__17749\,
            in3 => \N__17562\,
            lcout => n17298,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_2_lut_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17906\,
            in1 => \N__31407\,
            in2 => \_gnd_net_\,
            in3 => \N__17203\,
            lcout => n17544,
            ltout => OPEN,
            carryin => \bfn_1_28_0_\,
            carryout => \c0.tx2.n15675\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_3_lut_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17910\,
            in1 => \N__17850\,
            in2 => \_gnd_net_\,
            in3 => \N__17200\,
            lcout => n17504,
            ltout => OPEN,
            carryin => \c0.tx2.n15675\,
            carryout => \c0.tx2.n15676\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_4_lut_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17908\,
            in1 => \N__17674\,
            in2 => \_gnd_net_\,
            in3 => \N__17197\,
            lcout => n17570,
            ltout => OPEN,
            carryin => \c0.tx2.n15676\,
            carryout => \c0.tx2.n15677\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_5_lut_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17909\,
            in1 => \N__17658\,
            in2 => \_gnd_net_\,
            in3 => \N__17188\,
            lcout => n17457,
            ltout => OPEN,
            carryin => \c0.tx2.n15677\,
            carryout => \c0.tx2.n15678\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_6_lut_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17907\,
            in1 => \N__19570\,
            in2 => \_gnd_net_\,
            in3 => \N__17185\,
            lcout => n17567,
            ltout => OPEN,
            carryin => \c0.tx2.n15678\,
            carryout => \c0.tx2.n15679\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_7_lut_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17911\,
            in1 => \N__17871\,
            in2 => \_gnd_net_\,
            in3 => \N__17182\,
            lcout => n17629,
            ltout => OPEN,
            carryin => \c0.tx2.n15679\,
            carryout => \c0.tx2.n15680\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_8_lut_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17246\,
            in1 => \N__26382\,
            in2 => \_gnd_net_\,
            in3 => \N__17179\,
            lcout => n17634,
            ltout => OPEN,
            carryin => \c0.tx2.n15680\,
            carryout => \c0.tx2.n15681\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_9_lut_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17247\,
            in1 => \N__17805\,
            in2 => \_gnd_net_\,
            in3 => \N__17176\,
            lcout => n17640,
            ltout => OPEN,
            carryin => \c0.tx2.n15681\,
            carryout => \c0.tx2.n15682\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_10_lut_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17248\,
            in1 => \N__17781\,
            in2 => \_gnd_net_\,
            in3 => \N__17257\,
            lcout => n17458,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i7_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31513\,
            in1 => \N__17806\,
            in2 => \_gnd_net_\,
            in3 => \N__17254\,
            lcout => \r_Clock_Count_7_adj_2447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50447\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_777_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001110"
        )
    port map (
            in0 => \N__17886\,
            in1 => \N__17230\,
            in2 => \N__17827\,
            in3 => \N__30996\,
            lcout => n16824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_797_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__30995\,
            in1 => \N__17760\,
            in2 => \N__31514\,
            in3 => \N__17885\,
            lcout => n10_adj_2412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30994\,
            lcout => n9403,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i8_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17782\,
            in1 => \N__31485\,
            in2 => \_gnd_net_\,
            in3 => \N__17224\,
            lcout => \r_Clock_Count_8_adj_2446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50447\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18099\,
            in1 => \N__17977\,
            in2 => \_gnd_net_\,
            in3 => \N__17218\,
            lcout => n17542,
            ltout => OPEN,
            carryin => \bfn_1_30_0_\,
            carryout => \c0.tx.n15660\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_3_lut_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18095\,
            in1 => \N__18676\,
            in2 => \_gnd_net_\,
            in3 => \N__17215\,
            lcout => n17461,
            ltout => OPEN,
            carryin => \c0.tx.n15660\,
            carryout => \c0.tx.n15661\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_4_lut_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18100\,
            in1 => \N__18010\,
            in2 => \_gnd_net_\,
            in3 => \N__17212\,
            lcout => n17484,
            ltout => OPEN,
            carryin => \c0.tx.n15661\,
            carryout => \c0.tx.n15662\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_5_lut_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18096\,
            in1 => \N__17994\,
            in2 => \_gnd_net_\,
            in3 => \N__17278\,
            lcout => n17494,
            ltout => OPEN,
            carryin => \c0.tx.n15662\,
            carryout => \c0.tx.n15663\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_6_lut_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18098\,
            in1 => \N__19723\,
            in2 => \_gnd_net_\,
            in3 => \N__17275\,
            lcout => n17573,
            ltout => OPEN,
            carryin => \c0.tx.n15663\,
            carryout => \c0.tx.n15664\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_7_lut_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18097\,
            in1 => \N__17961\,
            in2 => \_gnd_net_\,
            in3 => \N__17272\,
            lcout => n17631,
            ltout => OPEN,
            carryin => \c0.tx.n15664\,
            carryout => \c0.tx.n15665\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_8_lut_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18449\,
            in1 => \N__19834\,
            in2 => \_gnd_net_\,
            in3 => \N__17269\,
            lcout => n17636,
            ltout => OPEN,
            carryin => \c0.tx.n15665\,
            carryout => \c0.tx.n15666\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_9_lut_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18450\,
            in1 => \N__19863\,
            in2 => \_gnd_net_\,
            in3 => \N__17266\,
            lcout => n17641,
            ltout => OPEN,
            carryin => \c0.tx.n15666\,
            carryout => \c0.tx.n15667\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_10_lut_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__19792\,
            in1 => \N__18454\,
            in2 => \_gnd_net_\,
            in3 => \N__17263\,
            lcout => OPEN,
            ltout => \n17537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i8_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23969\,
            in1 => \_gnd_net_\,
            in2 => \N__17260\,
            in3 => \N__19793\,
            lcout => \r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15303_3_lut_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__33880\,
            in1 => \N__33780\,
            in2 => \_gnd_net_\,
            in3 => \N__33754\,
            lcout => n17601,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__19679\,
            in1 => \N__18212\,
            in2 => \N__18772\,
            in3 => \N__17941\,
            lcout => \c0.rx.r_SM_Main_2_N_2090_2\,
            ltout => \c0.rx.r_SM_Main_2_N_2090_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15361_2_lut_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__33881\,
            in1 => \_gnd_net_\,
            in2 => \N__17323\,
            in3 => \_gnd_net_\,
            lcout => n17602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i5_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23968\,
            in1 => \N__17962\,
            in2 => \_gnd_net_\,
            in3 => \N__17320\,
            lcout => \r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_796_LC_1_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__17302\,
            in1 => \N__17939\,
            in2 => \N__33885\,
            in3 => \N__18770\,
            lcout => OPEN,
            ltout => \n16810_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_1_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__20147\,
            in1 => \N__30770\,
            in2 => \N__17314\,
            in3 => \N__17308\,
            lcout => n16852,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i11107_2_lut_LC_1_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17938\,
            in2 => \_gnd_net_\,
            in3 => \N__18769\,
            lcout => OPEN,
            ltout => \c0.rx.n13452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_adj_398_LC_1_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__30769\,
            in1 => \N__30830\,
            in2 => \N__17311\,
            in3 => \N__17301\,
            lcout => n16867,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i14784_2_lut_LC_1_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18211\,
            in2 => \_gnd_net_\,
            in3 => \N__19680\,
            lcout => n17222,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_1_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__17940\,
            in1 => \N__18771\,
            in2 => \N__19684\,
            in3 => \N__18217\,
            lcout => \r_SM_Main_2_adj_2439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50482\,
            ce => 'H',
            sr => \N__17293\
        );

    \c0.i3_4_lut_adj_457_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17390\,
            in1 => \N__17411\,
            in2 => \N__17362\,
            in3 => \N__18140\,
            lcout => \c0.n16772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i7_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34661\,
            lcout => \c0.FRAME_MATCHER_state_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50381\,
            ce => 'H',
            sr => \N__17401\
        );

    \c0.i1_2_lut_adj_711_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17412\,
            in2 => \_gnd_net_\,
            in3 => \N__32567\,
            lcout => \c0.n16443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_726_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32584\,
            in3 => \N__17391\,
            lcout => \c0.n16447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_721_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32571\,
            lcout => \c0.n16451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_730_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18141\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29966\,
            lcout => \c0.n16349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_709_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21775\,
            in2 => \_gnd_net_\,
            in3 => \N__32566\,
            lcout => \c0.n16441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_713_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30109\,
            in2 => \N__32583\,
            in3 => \_gnd_net_\,
            lcout => \c0.n16445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i9_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33225\,
            in1 => \N__33005\,
            in2 => \_gnd_net_\,
            in3 => \N__18952\,
            lcout => \c0.FRAME_MATCHER_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50384\,
            ce => 'H',
            sr => \N__20446\
        );

    \c0.FRAME_MATCHER_state_i30_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__34659\,
            in1 => \N__21710\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_state_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50388\,
            ce => 'H',
            sr => \N__18280\
        );

    \c0.FRAME_MATCHER_i_i31_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33256\,
            in1 => \N__32910\,
            in2 => \_gnd_net_\,
            in3 => \N__19492\,
            lcout => \c0.FRAME_MATCHER_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50394\,
            ce => 'H',
            sr => \N__18817\
        );

    \c0.FRAME_MATCHER_i_i3_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33260\,
            in1 => \N__32960\,
            in2 => \_gnd_net_\,
            in3 => \N__18841\,
            lcout => \c0.FRAME_MATCHER_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50401\,
            ce => 'H',
            sr => \N__18292\
        );

    \c0.FRAME_MATCHER_i_i14_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33265\,
            in1 => \N__32997\,
            in2 => \_gnd_net_\,
            in3 => \N__19057\,
            lcout => \c0.FRAME_MATCHER_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50407\,
            ce => 'H',
            sr => \N__18328\
        );

    \c0.FRAME_MATCHER_i_i19_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33267\,
            in1 => \N__32998\,
            in2 => \_gnd_net_\,
            in3 => \N__19018\,
            lcout => \c0.FRAME_MATCHER_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50414\,
            ce => 'H',
            sr => \N__20386\
        );

    \blink_counter_2352__i0_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17467\,
            in2 => \_gnd_net_\,
            in3 => \N__17461\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_2_25_0_\,
            carryout => n15590,
            clk => \N__50424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i1_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17458\,
            in2 => \_gnd_net_\,
            in3 => \N__17452\,
            lcout => n25,
            ltout => OPEN,
            carryin => n15590,
            carryout => n15591,
            clk => \N__50424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i2_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17449\,
            in2 => \_gnd_net_\,
            in3 => \N__17443\,
            lcout => n24,
            ltout => OPEN,
            carryin => n15591,
            carryout => n15592,
            clk => \N__50424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i3_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17440\,
            in2 => \_gnd_net_\,
            in3 => \N__17434\,
            lcout => n23,
            ltout => OPEN,
            carryin => n15592,
            carryout => n15593,
            clk => \N__50424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i4_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17431\,
            in2 => \_gnd_net_\,
            in3 => \N__17425\,
            lcout => n22,
            ltout => OPEN,
            carryin => n15593,
            carryout => n15594,
            clk => \N__50424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i5_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17422\,
            in2 => \_gnd_net_\,
            in3 => \N__17416\,
            lcout => n21,
            ltout => OPEN,
            carryin => n15594,
            carryout => n15595,
            clk => \N__50424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i6_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17545\,
            in2 => \_gnd_net_\,
            in3 => \N__17539\,
            lcout => n20,
            ltout => OPEN,
            carryin => n15595,
            carryout => n15596,
            clk => \N__50424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i7_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17536\,
            in2 => \_gnd_net_\,
            in3 => \N__17530\,
            lcout => n19,
            ltout => OPEN,
            carryin => n15596,
            carryout => n15597,
            clk => \N__50424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i8_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17527\,
            in2 => \_gnd_net_\,
            in3 => \N__17521\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_2_26_0_\,
            carryout => n15598,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i9_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17518\,
            in2 => \_gnd_net_\,
            in3 => \N__17512\,
            lcout => n17_adj_2422,
            ltout => OPEN,
            carryin => n15598,
            carryout => n15599,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i10_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17509\,
            in2 => \_gnd_net_\,
            in3 => \N__17503\,
            lcout => n16,
            ltout => OPEN,
            carryin => n15599,
            carryout => n15600,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i11_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17500\,
            in2 => \_gnd_net_\,
            in3 => \N__17494\,
            lcout => n15,
            ltout => OPEN,
            carryin => n15600,
            carryout => n15601,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i12_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17491\,
            in2 => \_gnd_net_\,
            in3 => \N__17485\,
            lcout => n14_adj_2424,
            ltout => OPEN,
            carryin => n15601,
            carryout => n15602,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i13_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17482\,
            in2 => \_gnd_net_\,
            in3 => \N__17476\,
            lcout => n13,
            ltout => OPEN,
            carryin => n15602,
            carryout => n15603,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i14_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17473\,
            in2 => \_gnd_net_\,
            in3 => \N__17641\,
            lcout => n12_adj_2419,
            ltout => OPEN,
            carryin => n15603,
            carryout => n15604,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i15_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17638\,
            in2 => \_gnd_net_\,
            in3 => \N__17632\,
            lcout => n11,
            ltout => OPEN,
            carryin => n15604,
            carryout => n15605,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i16_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17629\,
            in2 => \_gnd_net_\,
            in3 => \N__17623\,
            lcout => n10_adj_2420,
            ltout => OPEN,
            carryin => \bfn_2_27_0_\,
            carryout => n15606,
            clk => \N__50439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i17_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17620\,
            in2 => \_gnd_net_\,
            in3 => \N__17614\,
            lcout => n9,
            ltout => OPEN,
            carryin => n15606,
            carryout => n15607,
            clk => \N__50439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i18_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17611\,
            in2 => \_gnd_net_\,
            in3 => \N__17605\,
            lcout => n8,
            ltout => OPEN,
            carryin => n15607,
            carryout => n15608,
            clk => \N__50439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i19_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17602\,
            in2 => \_gnd_net_\,
            in3 => \N__17596\,
            lcout => n7,
            ltout => OPEN,
            carryin => n15608,
            carryout => n15609,
            clk => \N__50439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i20_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17593\,
            in2 => \_gnd_net_\,
            in3 => \N__17587\,
            lcout => n6_adj_2421,
            ltout => OPEN,
            carryin => n15609,
            carryout => n15610,
            clk => \N__50439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i21_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17577\,
            in2 => \_gnd_net_\,
            in3 => \N__17566\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n15610,
            carryout => n15611,
            clk => \N__50439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i22_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17561\,
            in2 => \_gnd_net_\,
            in3 => \N__17548\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n15611,
            carryout => n15612,
            clk => \N__50439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i23_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17744\,
            in2 => \_gnd_net_\,
            in3 => \N__17731\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n15612,
            carryout => n15613,
            clk => \N__50439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i24_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17723\,
            in2 => \_gnd_net_\,
            in3 => \N__17710\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_2_28_0_\,
            carryout => n15614,
            clk => \N__50448\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2352__i25_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17703\,
            in2 => \_gnd_net_\,
            in3 => \N__17707\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50448\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__30759\,
            in1 => \N__30864\,
            in2 => \N__33886\,
            in3 => \N__18413\,
            lcout => \c0.rx.n9323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i2_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31497\,
            in1 => \N__17692\,
            in2 => \_gnd_net_\,
            in3 => \N__17673\,
            lcout => \r_Clock_Count_2_adj_2452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50448\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000101000"
        )
    port map (
            in0 => \N__24065\,
            in1 => \N__20812\,
            in2 => \N__31361\,
            in3 => \N__19752\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50448\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i5_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31498\,
            in1 => \N__17872\,
            in2 => \_gnd_net_\,
            in3 => \N__17686\,
            lcout => \r_Clock_Count_5_adj_2449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50448\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i1_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__31496\,
            in1 => \N__17680\,
            in2 => \N__17854\,
            in3 => \_gnd_net_\,
            lcout => \r_Clock_Count_1_adj_2453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50448\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4_4_lut_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19569\,
            in1 => \N__17672\,
            in2 => \N__31408\,
            in3 => \N__17657\,
            lcout => \c0.tx2.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14702_3_lut_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__31486\,
            in1 => \N__30997\,
            in2 => \_gnd_net_\,
            in3 => \N__17887\,
            lcout => OPEN,
            ltout => \n17140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14847_4_lut_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101111"
        )
    port map (
            in0 => \N__17920\,
            in1 => \N__17761\,
            in2 => \N__17914\,
            in3 => \N__17823\,
            lcout => n16817,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_4_lut_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__26390\,
            in1 => \N__17802\,
            in2 => \N__29344\,
            in3 => \N__17778\,
            lcout => n12_adj_2410,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5_3_lut_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17870\,
            in1 => \N__17849\,
            in2 => \_gnd_net_\,
            in3 => \N__17833\,
            lcout => n15837,
            ltout => \n15837_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_4_lut_adj_399_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26392\,
            in1 => \N__17804\,
            in2 => \N__17812\,
            in3 => \N__17780\,
            lcout => \r_SM_Main_2_N_2033_1\,
            ltout => \r_SM_Main_2_N_2033_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i1_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__29325\,
            in1 => \N__31014\,
            in2 => \N__17809\,
            in3 => \N__31488\,
            lcout => \r_SM_Main_1_adj_2444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_4_lut_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26391\,
            in1 => \N__17803\,
            in2 => \N__29343\,
            in3 => \N__17779\,
            lcout => n9929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i2_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29326\,
            in1 => \N__31487\,
            in2 => \N__31021\,
            in3 => \N__20004\,
            lcout => \r_SM_Main_2_adj_2443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i2_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__18069\,
            in1 => \N__18049\,
            in2 => \_gnd_net_\,
            in3 => \N__20137\,
            lcout => \r_Clock_Count_2_adj_2435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i3_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23970\,
            in1 => \N__18034\,
            in2 => \_gnd_net_\,
            in3 => \N__17993\,
            lcout => \r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23959\,
            in1 => \N__18028\,
            in2 => \_gnd_net_\,
            in3 => \N__17976\,
            lcout => \r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i2_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__18009\,
            in1 => \_gnd_net_\,
            in2 => \N__18022\,
            in3 => \N__23960\,
            lcout => \r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_793_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__30848\,
            in1 => \N__30735\,
            in2 => \N__33876\,
            in3 => \N__18115\,
            lcout => n17_adj_2416,
            ltout => \n17_adj_2416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i4_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18630\,
            in2 => \N__18013\,
            in3 => \N__18235\,
            lcout => \r_Clock_Count_4_adj_2433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4_4_lut_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19722\,
            in1 => \N__18008\,
            in2 => \N__17995\,
            in3 => \N__17975\,
            lcout => OPEN,
            ltout => \c0.tx.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5_3_lut_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17960\,
            in2 => \N__17944\,
            in3 => \N__18671\,
            lcout => n15701,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18065\,
            in1 => \N__20101\,
            in2 => \N__18717\,
            in3 => \N__18610\,
            lcout => n16863,
            ltout => \n16863_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__18747\,
            in1 => \N__18209\,
            in2 => \N__17923\,
            in3 => \N__19672\,
            lcout => \c0.rx.r_SM_Main_2_N_2096_0\,
            ltout => \c0.rx.r_SM_Main_2_N_2096_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_adj_397_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18118\,
            in3 => \N__33747\,
            lcout => n6_adj_2461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i7_LC_2_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23961\,
            in1 => \N__19864\,
            in2 => \_gnd_net_\,
            in3 => \N__18109\,
            lcout => \r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i7_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__18210\,
            in1 => \N__18148\,
            in2 => \_gnd_net_\,
            in3 => \N__20139\,
            lcout => \r_Clock_Count_7_adj_2430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14706_3_lut_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__24066\,
            in1 => \N__23957\,
            in2 => \_gnd_net_\,
            in3 => \N__18499\,
            lcout => OPEN,
            ltout => \n17144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14845_4_lut_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101000101"
        )
    port map (
            in0 => \N__18471\,
            in1 => \N__18694\,
            in2 => \N__18103\,
            in3 => \N__19774\,
            lcout => n16828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_2_lut_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18175\,
            in1 => \N__20100\,
            in2 => \_gnd_net_\,
            in3 => \N__18076\,
            lcout => n16859,
            ltout => OPEN,
            carryin => \bfn_2_32_0_\,
            carryout => \c0.rx.n15668\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_3_lut_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18179\,
            in1 => \_gnd_net_\,
            in2 => \N__18595\,
            in3 => \N__18073\,
            lcout => n16853,
            ltout => OPEN,
            carryin => \c0.rx.n15668\,
            carryout => \c0.rx.n15669\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_4_lut_LC_2_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18176\,
            in1 => \N__18070\,
            in2 => \_gnd_net_\,
            in3 => \N__18040\,
            lcout => n16860,
            ltout => OPEN,
            carryin => \c0.rx.n15669\,
            carryout => \c0.rx.n15670\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_5_lut_LC_2_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18180\,
            in1 => \N__18713\,
            in2 => \_gnd_net_\,
            in3 => \N__18037\,
            lcout => n16858,
            ltout => OPEN,
            carryin => \c0.rx.n15670\,
            carryout => \c0.rx.n15671\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_6_lut_LC_2_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18177\,
            in1 => \N__18631\,
            in2 => \_gnd_net_\,
            in3 => \N__18226\,
            lcout => n16854,
            ltout => OPEN,
            carryin => \c0.rx.n15671\,
            carryout => \c0.rx.n15672\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_7_lut_LC_2_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18181\,
            in1 => \N__18756\,
            in2 => \_gnd_net_\,
            in3 => \N__18223\,
            lcout => n16857,
            ltout => OPEN,
            carryin => \c0.rx.n15672\,
            carryout => \c0.rx.n15673\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_8_lut_LC_2_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18174\,
            in1 => \N__19678\,
            in2 => \_gnd_net_\,
            in3 => \N__18220\,
            lcout => n16856,
            ltout => OPEN,
            carryin => \c0.rx.n15673\,
            carryout => \c0.rx.n15674\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_9_lut_LC_2_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__18213\,
            in1 => \N__18178\,
            in2 => \_gnd_net_\,
            in3 => \N__18151\,
            lcout => n16855,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__5__2252_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31228\,
            in1 => \N__27801\,
            in2 => \_gnd_net_\,
            in3 => \N__25908\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i15_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18142\,
            in2 => \_gnd_net_\,
            in3 => \N__34642\,
            lcout => \c0.FRAME_MATCHER_state_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50385\,
            ce => 'H',
            sr => \N__18127\
        );

    \c0.i10728_2_lut_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32260\,
            in2 => \_gnd_net_\,
            in3 => \N__23253\,
            lcout => n1651,
            ltout => \n1651_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_776_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__21388\,
            in1 => \N__21676\,
            in2 => \N__18121\,
            in3 => \N__22279\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10657_3_lut_4_lut_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__21583\,
            in1 => \N__32261\,
            in2 => \N__22287\,
            in3 => \N__23254\,
            lcout => \FRAME_MATCHER_state_31_N_1440_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_775_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__27907\,
            in1 => \N__28036\,
            in2 => \N__22309\,
            in3 => \N__22280\,
            lcout => OPEN,
            ltout => \n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010101"
        )
    port map (
            in0 => \N__32454\,
            in1 => \N__18268\,
            in2 => \N__18262\,
            in3 => \N__18259\,
            lcout => OPEN,
            ltout => \n8_adj_2459_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i1_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__33278\,
            in1 => \N__18244\,
            in2 => \N__18253\,
            in3 => \N__18250\,
            lcout => \FRAME_MATCHER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_798_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110000"
        )
    port map (
            in0 => \N__32268\,
            in1 => \N__22354\,
            in2 => \N__22288\,
            in3 => \N__23255\,
            lcout => n3_adj_2408,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_725_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__18787\,
            in1 => \N__32892\,
            in2 => \N__22702\,
            in3 => \N__22324\,
            lcout => \c0.n4_adj_2360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i27_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25328\,
            in2 => \_gnd_net_\,
            in3 => \N__34643\,
            lcout => \c0.FRAME_MATCHER_state_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50395\,
            ce => 'H',
            sr => \N__25309\
        );

    \c0.i10765_2_lut_3_lut_4_lut_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23428\,
            in1 => \N__23258\,
            in2 => \N__24440\,
            in3 => \N__23049\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_5\,
            ltout => \c0.FRAME_MATCHER_i_31_N_1312_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_5_i3_2_lut_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__29728\,
            in1 => \_gnd_net_\,
            in2 => \N__18238\,
            in3 => \_gnd_net_\,
            lcout => \c0.n3_adj_2256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i5_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33255\,
            in1 => \N__32896\,
            in2 => \_gnd_net_\,
            in3 => \N__18988\,
            lcout => \c0.FRAME_MATCHER_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50402\,
            ce => 'H',
            sr => \N__18310\
        );

    \c0.i10766_2_lut_3_lut_4_lut_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23259\,
            in1 => \N__24491\,
            in2 => \N__23064\,
            in3 => \N__23426\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_4\,
            ltout => \c0.FRAME_MATCHER_i_31_N_1312_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_4_i3_2_lut_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18298\,
            in3 => \N__29727\,
            lcout => \c0.n3_adj_2257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10767_2_lut_3_lut_4_lut_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23260\,
            in1 => \N__25120\,
            in2 => \N__23065\,
            in3 => \N__23427\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_3\,
            ltout => \c0.FRAME_MATCHER_i_31_N_1312_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_3_i3_2_lut_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18295\,
            in3 => \N__29726\,
            lcout => \c0.n3_adj_2258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_42_i10_2_lut_3_lut_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__25116\,
            in1 => \N__24490\,
            in2 => \_gnd_net_\,
            in3 => \N__24429\,
            lcout => \c0.n10_adj_2329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i13_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__32912\,
            in1 => \N__33258\,
            in2 => \_gnd_net_\,
            in3 => \N__19075\,
            lcout => \c0.FRAME_MATCHER_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50408\,
            ce => 'H',
            sr => \N__18322\
        );

    \c0.i1_2_lut_adj_762_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21712\,
            in2 => \_gnd_net_\,
            in3 => \N__29941\,
            lcout => \c0.n16379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30027\,
            in2 => \_gnd_net_\,
            in3 => \N__30117\,
            lcout => \c0.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i10739_2_lut_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19927\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19975\,
            lcout => n13082,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_400_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31728\,
            in2 => \_gnd_net_\,
            in3 => \N__31672\,
            lcout => n445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10755_2_lut_3_lut_4_lut_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23417\,
            in1 => \N__22996\,
            in2 => \N__28249\,
            in3 => \N__23236\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i15_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__32913\,
            in1 => \N__33259\,
            in2 => \_gnd_net_\,
            in3 => \N__19036\,
            lcout => \c0.FRAME_MATCHER_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50415\,
            ce => 'H',
            sr => \N__18337\
        );

    \c0.select_238_Select_15_i3_2_lut_3_lut_4_lut_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29735\,
            in1 => \N__23008\,
            in2 => \N__28250\,
            in3 => \N__22704\,
            lcout => \c0.n3_adj_2242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10756_2_lut_3_lut_4_lut_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23237\,
            in1 => \N__28283\,
            in2 => \N__23046\,
            in3 => \N__23415\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_14_i3_2_lut_3_lut_4_lut_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29734\,
            in1 => \N__23007\,
            in2 => \N__28290\,
            in3 => \N__22705\,
            lcout => \c0.n3_adj_2243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10757_2_lut_3_lut_4_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23238\,
            in1 => \N__24337\,
            in2 => \N__23047\,
            in3 => \N__23418\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_13_i3_2_lut_3_lut_4_lut_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29733\,
            in1 => \N__23006\,
            in2 => \N__24347\,
            in3 => \N__22703\,
            lcout => \c0.n3_adj_2244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10758_2_lut_3_lut_4_lut_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23239\,
            in1 => \N__25470\,
            in2 => \N__23048\,
            in3 => \N__23416\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i25_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__32914\,
            in1 => \N__33261\,
            in2 => \_gnd_net_\,
            in3 => \N__19150\,
            lcout => \c0.FRAME_MATCHER_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50425\,
            ce => 'H',
            sr => \N__20290\
        );

    \c0.data_in_1__0__2273_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27744\,
            in1 => \N__23572\,
            in2 => \_gnd_net_\,
            in3 => \N__20052\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_54_i4_2_lut_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__19918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19971\,
            lcout => n4_adj_2460,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20718\,
            in1 => \N__33764\,
            in2 => \N__26490\,
            in3 => \N__20508\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__0__2265_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23573\,
            in1 => \N__22110\,
            in2 => \_gnd_net_\,
            in3 => \N__27746\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__20539\,
            in1 => \N__33763\,
            in2 => \N__31202\,
            in3 => \N__20507\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__1__2272_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19252\,
            in1 => \N__22408\,
            in2 => \_gnd_net_\,
            in3 => \N__27745\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__5__2276_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27743\,
            in1 => \N__22077\,
            in2 => \_gnd_net_\,
            in3 => \N__18367\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__3__2270_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20595\,
            in1 => \N__27708\,
            in2 => \_gnd_net_\,
            in3 => \N__19542\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14734_2_lut_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20048\,
            in2 => \_gnd_net_\,
            in3 => \N__20594\,
            lcout => OPEN,
            ltout => \c0.n17172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14824_4_lut_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18348\,
            in1 => \N__18365\,
            in2 => \N__18340\,
            in3 => \N__18378\,
            lcout => \c0.n17262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_567_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__25084\,
            in1 => \N__21653\,
            in2 => \_gnd_net_\,
            in3 => \N__32705\,
            lcout => \c0.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__7__2274_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18379\,
            in1 => \N__23539\,
            in2 => \_gnd_net_\,
            in3 => \N__27709\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14826_3_lut_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19541\,
            in1 => \N__19476\,
            in2 => \_gnd_net_\,
            in3 => \N__19599\,
            lcout => \c0.n17264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__5__2268_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18366\,
            in1 => \N__25894\,
            in2 => \_gnd_net_\,
            in3 => \N__27710\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__4__2277_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27707\,
            in1 => \N__19600\,
            in2 => \_gnd_net_\,
            in3 => \N__18349\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i75_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__26936\,
            in1 => \N__28803\,
            in2 => \N__22563\,
            in3 => \N__31135\,
            lcout => \c0.data_in_frame_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__1__2256_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27705\,
            in1 => \_gnd_net_\,
            in2 => \N__30665\,
            in3 => \N__19272\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4216_2_lut_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27248\,
            in2 => \_gnd_net_\,
            in3 => \N__29342\,
            lcout => \c0.tx2.n6480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__6__2275_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27704\,
            in1 => \N__19477\,
            in2 => \_gnd_net_\,
            in3 => \N__27610\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20697\,
            in2 => \_gnd_net_\,
            in3 => \N__20658\,
            lcout => n9472,
            ltout => \n9472_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__30649\,
            in1 => \N__20625\,
            in2 => \N__18427\,
            in3 => \N__33753\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13_4_lut_4_lut_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000101"
        )
    port map (
            in0 => \N__30760\,
            in1 => \N__30875\,
            in2 => \N__33859\,
            in3 => \N__18420\,
            lcout => OPEN,
            ltout => \c0.rx.n10086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__27706\,
            in1 => \N__30761\,
            in2 => \N__18424\,
            in3 => \N__30876\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i57_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25585\,
            in1 => \N__25770\,
            in2 => \_gnd_net_\,
            in3 => \N__20845\,
            lcout => data_in_frame_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50459\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14959_3_lut_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31343\,
            in1 => \N__35443\,
            in2 => \_gnd_net_\,
            in3 => \N__29368\,
            lcout => n17397,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i10646_2_lut_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29320\,
            in2 => \_gnd_net_\,
            in3 => \N__20001\,
            lcout => \c0.tx2.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_56_i4_2_lut_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19961\,
            in2 => \_gnd_net_\,
            in3 => \N__19917\,
            lcout => n4_adj_2409,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100110011"
        )
    port map (
            in0 => \N__18574\,
            in1 => \N__33858\,
            in2 => \N__19970\,
            in3 => \N__18421\,
            lcout => n13440,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_4_lut_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19804\,
            in1 => \N__19825\,
            in2 => \N__19872\,
            in3 => \N__18470\,
            lcout => n14060,
            ltout => \n14060_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i14754_4_lut_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__24156\,
            in1 => \N__24043\,
            in2 => \N__18382\,
            in3 => \N__23892\,
            lcout => \c0.tx.n14082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001110"
        )
    port map (
            in0 => \N__24169\,
            in1 => \N__19630\,
            in2 => \N__23933\,
            in3 => \N__24103\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5592_4_lut_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__31013\,
            in1 => \N__27249\,
            in2 => \N__29239\,
            in3 => \N__20002\,
            lcout => OPEN,
            ltout => \n7866_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i0_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100110000"
        )
    port map (
            in0 => \N__20003\,
            in1 => \N__31499\,
            in2 => \N__18505\,
            in3 => \N__29327\,
            lcout => \r_SM_Main_0_adj_2445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i14832_3_lut_4_lut_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__18572\,
            in1 => \N__30749\,
            in2 => \N__19969\,
            in3 => \N__18550\,
            lcout => n10425,
            ltout => \n10425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000011000000"
        )
    port map (
            in0 => \N__18551\,
            in1 => \N__19957\,
            in2 => \N__18502\,
            in3 => \N__18573\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_4_lut_adj_402_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__19824\,
            in1 => \N__19865\,
            in2 => \N__24171\,
            in3 => \N__19803\,
            lcout => n12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i10933_2_lut_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24039\,
            in2 => \_gnd_net_\,
            in3 => \N__23953\,
            lcout => n13276,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__23954\,
            in1 => \N__19767\,
            in2 => \N__24064\,
            in3 => \N__18497\,
            lcout => OPEN,
            ltout => \n10_adj_2415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_789_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110010"
        )
    port map (
            in0 => \N__18498\,
            in1 => \N__18481\,
            in2 => \N__18475\,
            in3 => \N__18472\,
            lcout => n16844,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__20693\,
            in1 => \N__18552\,
            in2 => \_gnd_net_\,
            in3 => \N__18520\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23958\,
            in1 => \N__18675\,
            in2 => \_gnd_net_\,
            in3 => \N__18685\,
            lcout => \r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000101010001"
        )
    port map (
            in0 => \N__30874\,
            in1 => \N__18655\,
            in2 => \N__30768\,
            in3 => \N__18643\,
            lcout => \r_SM_Main_1_adj_2440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18626\,
            in2 => \_gnd_net_\,
            in3 => \N__18587\,
            lcout => \c0.rx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i1_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__18588\,
            in1 => \N__18604\,
            in2 => \_gnd_net_\,
            in3 => \N__20138\,
            lcout => \r_Clock_Count_1_adj_2436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_3_lut_4_lut_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__31706\,
            in1 => \N__23956\,
            in2 => \N__24049\,
            in3 => \N__24172\,
            lcout => n8730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14840_4_lut_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21235\,
            in1 => \N__20929\,
            in2 => \N__20185\,
            in3 => \N__20026\,
            lcout => \c0.n17278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_395_LC_3_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19913\,
            in2 => \_gnd_net_\,
            in3 => \N__20685\,
            lcout => n4_adj_2411,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_3_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001000000000"
        )
    port map (
            in0 => \N__20686\,
            in1 => \N__18553\,
            in2 => \N__19925\,
            in3 => \N__18519\,
            lcout => \r_Bit_Index_1_adj_2438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i5_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__20141\,
            in1 => \N__18757\,
            in2 => \_gnd_net_\,
            in3 => \N__18778\,
            lcout => \r_Clock_Count_5_adj_2432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i3_LC_3_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__18718\,
            in1 => \N__18724\,
            in2 => \_gnd_net_\,
            in3 => \N__20140\,
            lcout => \r_Clock_Count_3_adj_2434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_3_lut_4_lut_LC_3_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__27532\,
            in1 => \N__24250\,
            in2 => \N__31721\,
            in3 => \N__31670\,
            lcout => n16886,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_401_LC_3_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__23955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24023\,
            lcout => n9406,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_2156_LC_3_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000010"
        )
    port map (
            in0 => \N__42607\,
            in1 => \N__27064\,
            in2 => \N__31612\,
            in3 => \N__27280\,
            lcout => \c0.r_SM_Main_2_N_2036_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50506\,
            ce => 'H',
            sr => \N__45550\
        );

    \c0.FRAME_MATCHER_i_i24_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33185\,
            in1 => \N__33007\,
            in2 => \_gnd_net_\,
            in3 => \N__19162\,
            lcout => \c0.FRAME_MATCHER_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50396\,
            ce => 'H',
            sr => \N__20317\
        );

    \c0.FRAME_MATCHER_i_i21_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33161\,
            in1 => \N__33006\,
            in2 => \_gnd_net_\,
            in3 => \N__19213\,
            lcout => \c0.FRAME_MATCHER_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50390\,
            ce => 'H',
            sr => \N__20233\
        );

    \c0.FRAME_MATCHER_i_i28_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33098\,
            in1 => \N__32989\,
            in2 => \_gnd_net_\,
            in3 => \N__19111\,
            lcout => \c0.FRAME_MATCHER_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50382\,
            ce => 'H',
            sr => \N__20227\
        );

    \c0.FRAME_MATCHER_i_i30_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33184\,
            in1 => \N__32947\,
            in2 => \_gnd_net_\,
            in3 => \N__19510\,
            lcout => \c0.FRAME_MATCHER_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50391\,
            ce => 'H',
            sr => \N__18823\
        );

    \c0.FRAME_MATCHER_i_i29_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33186\,
            in1 => \N__32893\,
            in2 => \_gnd_net_\,
            in3 => \N__19522\,
            lcout => \c0.FRAME_MATCHER_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50397\,
            ce => 'H',
            sr => \N__18832\
        );

    \c0.select_238_Select_29_i3_2_lut_3_lut_4_lut_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23036\,
            in1 => \N__29679\,
            in2 => \N__22163\,
            in3 => \N__22674\,
            lcout => \c0.n3_adj_2217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_30_i3_2_lut_3_lut_4_lut_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23037\,
            in1 => \N__29680\,
            in2 => \N__24908\,
            in3 => \N__22675\,
            lcout => \c0.n3_adj_2215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_31_i3_2_lut_3_lut_4_lut_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22672\,
            in1 => \N__22494\,
            in2 => \N__29711\,
            in3 => \N__23038\,
            lcout => \c0.n3_adj_2210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_8_i3_2_lut_3_lut_4_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23039\,
            in1 => \N__29684\,
            in2 => \N__24868\,
            in3 => \N__22673\,
            lcout => \c0.n3_adj_2249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_700_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__22493\,
            in1 => \N__25179\,
            in2 => \_gnd_net_\,
            in3 => \N__23035\,
            lcout => \c0.n9393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i6_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33181\,
            in1 => \N__32946\,
            in2 => \_gnd_net_\,
            in3 => \N__18979\,
            lcout => \c0.FRAME_MATCHER_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50403\,
            ce => 'H',
            sr => \N__20392\
        );

    \c0.i10768_2_lut_3_lut_4_lut_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23430\,
            in1 => \N__23256\,
            in2 => \N__25080\,
            in3 => \N__23056\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_2\,
            ltout => \c0.FRAME_MATCHER_i_31_N_1312_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_2_i3_2_lut_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18781\,
            in3 => \N__29649\,
            lcout => \c0.n3_adj_2259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i2_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__32848\,
            in1 => \N__33254\,
            in2 => \_gnd_net_\,
            in3 => \N__18856\,
            lcout => \c0.FRAME_MATCHER_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50409\,
            ce => 'H',
            sr => \N__18931\
        );

    \c0.i1_2_lut_3_lut_adj_681_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__25066\,
            in1 => \N__21641\,
            in2 => \_gnd_net_\,
            in3 => \N__18913\,
            lcout => n16896,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_627_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__32690\,
            in1 => \N__18919\,
            in2 => \_gnd_net_\,
            in3 => \N__23714\,
            lcout => \c0.n16895\,
            ltout => \c0.n16895_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_651_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21640\,
            in2 => \N__18907\,
            in3 => \N__25062\,
            lcout => n16897,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10769_2_lut_3_lut_4_lut_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23429\,
            in1 => \N__23257\,
            in2 => \N__21652\,
            in3 => \N__23057\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_1\,
            ltout => \c0.FRAME_MATCHER_i_31_N_1312_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_1_i3_2_lut_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18904\,
            in3 => \N__29648\,
            lcout => \c0.n3_adj_2260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_2_lut_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__29574\,
            in1 => \N__19371\,
            in2 => \N__32709\,
            in3 => \N__18889\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_0\,
            ltout => OPEN,
            carryin => \bfn_4_22_0_\,
            carryout => \c0.n15622\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_3_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18886\,
            in1 => \N__21642\,
            in2 => \N__19439\,
            in3 => \N__18865\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_1\,
            ltout => OPEN,
            carryin => \c0.n15622\,
            carryout => \c0.n15623\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_4_lut_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__18862\,
            in1 => \N__19375\,
            in2 => \N__25073\,
            in3 => \N__18850\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_2\,
            ltout => OPEN,
            carryin => \c0.n15623\,
            carryout => \c0.n15624\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_5_lut_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18847\,
            in1 => \N__25122\,
            in2 => \N__19440\,
            in3 => \N__19006\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_3\,
            ltout => OPEN,
            carryin => \c0.n15624\,
            carryout => \c0.n15625\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_6_lut_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19003\,
            in1 => \N__19379\,
            in2 => \N__24511\,
            in3 => \N__18997\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_4\,
            ltout => OPEN,
            carryin => \c0.n15625\,
            carryout => \c0.n15626\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_7_lut_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18994\,
            in1 => \N__24433\,
            in2 => \N__19441\,
            in3 => \N__18982\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_5\,
            ltout => OPEN,
            carryin => \c0.n15626\,
            carryout => \c0.n15627\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_8_lut_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20398\,
            in1 => \N__19383\,
            in2 => \N__21925\,
            in3 => \N__18970\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_6\,
            ltout => OPEN,
            carryin => \c0.n15627\,
            carryout => \c0.n15628\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_9_lut_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20257\,
            in1 => \N__21880\,
            in2 => \N__19442\,
            in3 => \N__18967\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_7\,
            ltout => OPEN,
            carryin => \c0.n15628\,
            carryout => \c0.n15629\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_10_lut_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20434\,
            in1 => \N__24847\,
            in2 => \N__19443\,
            in3 => \N__18955\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_8\,
            ltout => OPEN,
            carryin => \bfn_4_23_0_\,
            carryout => \c0.n15630\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_11_lut_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20452\,
            in1 => \N__19390\,
            in2 => \N__21855\,
            in3 => \N__18940\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_9\,
            ltout => OPEN,
            carryin => \c0.n15630\,
            carryout => \c0.n15631\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_12_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20338\,
            in1 => \N__28184\,
            in2 => \N__19444\,
            in3 => \N__18937\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_10\,
            ltout => OPEN,
            carryin => \c0.n15631\,
            carryout => \c0.n15632\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_13_lut_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20359\,
            in1 => \N__19394\,
            in2 => \N__28322\,
            in3 => \N__18934\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_11\,
            ltout => OPEN,
            carryin => \c0.n15632\,
            carryout => \c0.n15633\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_14_lut_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19096\,
            in1 => \N__25469\,
            in2 => \N__19445\,
            in3 => \N__19087\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_12\,
            ltout => OPEN,
            carryin => \c0.n15633\,
            carryout => \c0.n15634\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_15_lut_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19084\,
            in1 => \N__19398\,
            in2 => \N__24349\,
            in3 => \N__19069\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_13\,
            ltout => OPEN,
            carryin => \c0.n15634\,
            carryout => \c0.n15635\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_16_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19066\,
            in1 => \N__28282\,
            in2 => \N__19446\,
            in3 => \N__19048\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_14\,
            ltout => OPEN,
            carryin => \c0.n15635\,
            carryout => \c0.n15636\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_17_lut_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19045\,
            in1 => \N__19402\,
            in2 => \N__28254\,
            in3 => \N__19030\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_15\,
            ltout => OPEN,
            carryin => \c0.n15636\,
            carryout => \c0.n15637\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_18_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23077\,
            in1 => \N__22752\,
            in2 => \N__19450\,
            in3 => \N__19027\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_16\,
            ltout => OPEN,
            carryin => \bfn_4_24_0_\,
            carryout => \c0.n15638\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_19_lut_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23440\,
            in1 => \N__28081\,
            in2 => \N__19454\,
            in3 => \N__19024\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_17\,
            ltout => OPEN,
            carryin => \c0.n15638\,
            carryout => \c0.n15639\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_20_lut_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22258\,
            in1 => \N__23483\,
            in2 => \N__19451\,
            in3 => \N__19021\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_18\,
            ltout => OPEN,
            carryin => \c0.n15639\,
            carryout => \c0.n15640\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_21_lut_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20428\,
            in1 => \N__19420\,
            in2 => \N__21519\,
            in3 => \N__19009\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_19\,
            ltout => OPEN,
            carryin => \c0.n15640\,
            carryout => \c0.n15641\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_22_lut_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20422\,
            in1 => \N__24546\,
            in2 => \N__19452\,
            in3 => \N__19216\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_20\,
            ltout => OPEN,
            carryin => \c0.n15641\,
            carryout => \c0.n15642\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_23_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20416\,
            in1 => \N__24403\,
            in2 => \N__19455\,
            in3 => \N__19198\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_21\,
            ltout => OPEN,
            carryin => \c0.n15642\,
            carryout => \c0.n15643\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_24_lut_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20458\,
            in1 => \N__24761\,
            in2 => \N__19453\,
            in3 => \N__19183\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_22\,
            ltout => OPEN,
            carryin => \c0.n15643\,
            carryout => \c0.n15644\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_25_lut_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20407\,
            in1 => \N__24722\,
            in2 => \N__19456\,
            in3 => \N__19165\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_23\,
            ltout => OPEN,
            carryin => \c0.n15644\,
            carryout => \c0.n15645\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_26_lut_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20470\,
            in1 => \N__19403\,
            in2 => \N__21472\,
            in3 => \N__19153\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_24\,
            ltout => OPEN,
            carryin => \bfn_4_25_0_\,
            carryout => \c0.n15646\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_27_lut_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20482\,
            in1 => \N__24667\,
            in2 => \N__19447\,
            in3 => \N__19144\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_25\,
            ltout => OPEN,
            carryin => \c0.n15646\,
            carryout => \c0.n15647\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_28_lut_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20464\,
            in1 => \N__24818\,
            in2 => \N__19436\,
            in3 => \N__19129\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_26\,
            ltout => OPEN,
            carryin => \c0.n15647\,
            carryout => \c0.n15648\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_29_lut_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20518\,
            in1 => \N__24955\,
            in2 => \N__19448\,
            in3 => \N__19114\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_27\,
            ltout => OPEN,
            carryin => \c0.n15648\,
            carryout => \c0.n15649\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_30_lut_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20476\,
            in1 => \N__25017\,
            in2 => \N__19437\,
            in3 => \N__19099\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_28\,
            ltout => OPEN,
            carryin => \c0.n15649\,
            carryout => \c0.n15650\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_31_lut_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22123\,
            in1 => \N__22162\,
            in2 => \N__19449\,
            in3 => \N__19513\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_29\,
            ltout => OPEN,
            carryin => \c0.n15650\,
            carryout => \c0.n15651\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_32_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20488\,
            in1 => \N__24907\,
            in2 => \N__19438\,
            in3 => \N__19498\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_30\,
            ltout => OPEN,
            carryin => \c0.n15651\,
            carryout => \c0.n15652\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_997_33_lut_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__19413\,
            in1 => \N__22500\,
            in2 => \N__20572\,
            in3 => \N__19495\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1280_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14836_4_lut_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22048\,
            in1 => \N__22099\,
            in2 => \N__26207\,
            in3 => \N__22073\,
            lcout => OPEN,
            ltout => \c0.n17274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_424_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__19540\,
            in1 => \N__19475\,
            in2 => \N__19459\,
            in3 => \N__19597\,
            lcout => \c0.n9490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__1__2264_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__27672\,
            in1 => \_gnd_net_\,
            in2 => \N__19251\,
            in3 => \N__19271\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15448_1_lut_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27671\,
            lcout => \c0.n17889\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_433_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19273\,
            in1 => \N__20610\,
            in2 => \N__19250\,
            in3 => \N__19610\,
            lcout => \c0.n12_adj_2158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i80_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__28764\,
            in1 => \N__23625\,
            in2 => \N__26539\,
            in3 => \N__31141\,
            lcout => \c0.data_in_frame_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__4__2261_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22049\,
            in1 => \_gnd_net_\,
            in2 => \N__27713\,
            in3 => \N__19611\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__4__2269_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19612\,
            in1 => \N__27673\,
            in2 => \_gnd_net_\,
            in3 => \N__19598\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i53_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31796\,
            in1 => \N__25992\,
            in2 => \_gnd_net_\,
            in3 => \N__25712\,
            lcout => data_in_frame_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i4_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19562\,
            in1 => \N__19582\,
            in2 => \_gnd_net_\,
            in3 => \N__31525\,
            lcout => \r_Clock_Count_4_adj_2450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i56_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26532\,
            in1 => \N__26049\,
            in2 => \_gnd_net_\,
            in3 => \N__25713\,
            lcout => data_in_frame_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__0__2257_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27711\,
            in1 => \_gnd_net_\,
            in2 => \N__25589\,
            in3 => \N__22106\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__3__2262_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25801\,
            in1 => \N__19543\,
            in2 => \_gnd_net_\,
            in3 => \N__27712\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i51_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26562\,
            in1 => \N__26911\,
            in2 => \_gnd_net_\,
            in3 => \N__25711\,
            lcout => data_in_frame_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i60_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30522\,
            in1 => \N__20850\,
            in2 => \_gnd_net_\,
            in3 => \N__28953\,
            lcout => data_in_frame_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_4_lut_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31028\,
            in1 => \N__31524\,
            in2 => \N__27259\,
            in3 => \N__29341\,
            lcout => \c0.tx2.n8737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i6_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__19696\,
            in1 => \N__19659\,
            in2 => \_gnd_net_\,
            in3 => \N__20158\,
            lcout => \r_Clock_Count_6_adj_2431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_678_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__32710\,
            in1 => \N__25086\,
            in2 => \N__21658\,
            in3 => \N__31988\,
            lcout => n16893,
            ltout => \n16893_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i62_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31217\,
            in1 => \_gnd_net_\,
            in2 => \N__19633\,
            in3 => \N__28908\,
            lcout => data_in_frame_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001000100"
        )
    port map (
            in0 => \N__20811\,
            in1 => \N__24063\,
            in2 => \_gnd_net_\,
            in3 => \N__19753\,
            lcout => \c0.tx.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i13_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__28802\,
            in1 => \N__28568\,
            in2 => \N__31830\,
            in3 => \N__31989\,
            lcout => \c0.data_in_frame_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i54_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31216\,
            in1 => \N__28851\,
            in2 => \_gnd_net_\,
            in3 => \N__25715\,
            lcout => data_in_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i52_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30523\,
            in1 => \N__26016\,
            in2 => \_gnd_net_\,
            in3 => \N__25714\,
            lcout => data_in_frame_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i9_3_lut_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24044\,
            in1 => \N__20818\,
            in2 => \_gnd_net_\,
            in3 => \N__31735\,
            lcout => n5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i6_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19827\,
            in1 => \N__23971\,
            in2 => \_gnd_net_\,
            in3 => \N__19624\,
            lcout => \r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i14756_4_lut_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__31022\,
            in1 => \N__29321\,
            in2 => \N__31546\,
            in3 => \N__20005\,
            lcout => n17194,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_52_i4_2_lut_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__19962\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19926\,
            lcout => n4_adj_2417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_4_lut_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19873\,
            in1 => \N__19826\,
            in2 => \N__24170\,
            in3 => \N__19802\,
            lcout => n9937,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i13245_2_lut_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20808\,
            in2 => \_gnd_net_\,
            in3 => \N__31383\,
            lcout => OPEN,
            ltout => \c0.tx.n15683_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001001000"
        )
    port map (
            in0 => \N__20763\,
            in1 => \N__24045\,
            in2 => \N__19756\,
            in3 => \N__19748\,
            lcout => \c0.tx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_483_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26725\,
            in1 => \N__21220\,
            in2 => \N__20923\,
            in3 => \N__26668\,
            lcout => \c0.n20_adj_2267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i4_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23962\,
            in1 => \N__19732\,
            in2 => \_gnd_net_\,
            in3 => \N__19721\,
            lcout => \r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_461_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21359\,
            in2 => \_gnd_net_\,
            in3 => \N__21326\,
            lcout => \c0.n12993\,
            ltout => \c0.n12993_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14838_4_lut_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21291\,
            in1 => \N__21129\,
            in2 => \N__19699\,
            in3 => \N__21066\,
            lcout => \c0.n17276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_462_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20876\,
            in2 => \_gnd_net_\,
            in3 => \N__21167\,
            lcout => \c0.n13298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i3_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__21168\,
            in1 => \N__27552\,
            in2 => \N__21154\,
            in3 => \N__20983\,
            lcout => \c0.delay_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i4_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__20984\,
            in1 => \N__26669\,
            in2 => \N__21142\,
            in3 => \N__27559\,
            lcout => \c0.delay_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i11_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__21327\,
            in1 => \N__27551\,
            in2 => \N__21313\,
            in3 => \N__20982\,
            lcout => \c0.delay_counter_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i1_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__27534\,
            in1 => \N__20860\,
            in2 => \N__20881\,
            in3 => \N__20985\,
            lcout => \c0.delay_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i5_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20987\,
            in1 => \N__21106\,
            in2 => \_gnd_net_\,
            in3 => \N__21130\,
            lcout => \c0.delay_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_1_lut_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27533\,
            lcout => n53,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_491_LC_4_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21064\,
            in1 => \N__20032\,
            in2 => \N__21290\,
            in3 => \N__20025\,
            lcout => OPEN,
            ltout => \c0.n21_adj_2271_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_540_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20014\,
            in2 => \N__20008\,
            in3 => \N__20173\,
            lcout => n29,
            ltout => \n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i9_LC_4_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__21001\,
            in1 => \N__21019\,
            in2 => \N__20194\,
            in3 => \N__20986\,
            lcout => \c0.delay_counter_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20073\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_464_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21097\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21017\,
            lcout => \c0.n12991\,
            ltout => \c0.n12991_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_489_LC_4_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26649\,
            in1 => \N__21127\,
            in2 => \N__20176\,
            in3 => \N__26699\,
            lcout => \c0.n19_adj_2270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__42592\,
            in1 => \N__46362\,
            in2 => \N__45952\,
            in3 => \N__27402\,
            lcout => n9361,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_4_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__24038\,
            in1 => \N__23964\,
            in2 => \N__24187\,
            in3 => \N__24115\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_4_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__20167\,
            in1 => \N__20096\,
            in2 => \_gnd_net_\,
            in3 => \N__20154\,
            lcout => \r_Clock_Count_0_adj_2437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_4_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20734\,
            in1 => \N__23963\,
            in2 => \_gnd_net_\,
            in3 => \N__20072\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i3_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33397\,
            in2 => \_gnd_net_\,
            in3 => \N__34652\,
            lcout => \c0.FRAME_MATCHER_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50416\,
            ce => 'H',
            sr => \N__21187\
        );

    \c0.data_in_0__0__2281_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__27800\,
            in1 => \_gnd_net_\,
            in2 => \N__22205\,
            in3 => \N__20059\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10680_2_lut_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22496\,
            in2 => \_gnd_net_\,
            in3 => \N__25180\,
            lcout => n3977,
            ltout => \n3977_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i2_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111111011"
        )
    port map (
            in0 => \N__21403\,
            in1 => \N__32447\,
            in2 => \N__20236\,
            in3 => \N__32996\,
            lcout => \FRAME_MATCHER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__32299\,
            in1 => \N__33476\,
            in2 => \_gnd_net_\,
            in3 => \N__29475\,
            lcout => \c0.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_21_i3_2_lut_3_lut_4_lut_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22691\,
            in1 => \N__29712\,
            in2 => \N__24388\,
            in3 => \N__23044\,
            lcout => \c0.n3_adj_2233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_28_i3_2_lut_3_lut_4_lut_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23045\,
            in1 => \N__24997\,
            in2 => \N__29732\,
            in3 => \N__22690\,
            lcout => \c0.n3_adj_2219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i6_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21774\,
            in2 => \_gnd_net_\,
            in3 => \N__34564\,
            lcout => \c0.FRAME_MATCHER_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50398\,
            ce => 'H',
            sr => \N__20218\
        );

    \c0.FRAME_MATCHER_state_i4_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30018\,
            in2 => \_gnd_net_\,
            in3 => \N__34561\,
            lcout => \c0.FRAME_MATCHER_state_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50404\,
            ce => 'H',
            sr => \N__29836\
        );

    \c0.select_238_Select_23_i3_2_lut_3_lut_4_lut_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29657\,
            in1 => \N__22667\,
            in2 => \N__24726\,
            in3 => \N__23059\,
            lcout => \c0.n3_adj_2229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14770_3_lut_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__32306\,
            in1 => \N__37387\,
            in2 => \_gnd_net_\,
            in3 => \N__21811\,
            lcout => n17208,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_22_i3_2_lut_3_lut_4_lut_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29656\,
            in1 => \N__22665\,
            in2 => \N__24772\,
            in3 => \N__23058\,
            lcout => \c0.n3_adj_2231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_24_i3_2_lut_3_lut_4_lut_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23060\,
            in1 => \N__21466\,
            in2 => \N__22700\,
            in3 => \N__29658\,
            lcout => \c0.n3_adj_2227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_26_i3_2_lut_3_lut_4_lut_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29660\,
            in1 => \N__22666\,
            in2 => \N__24822\,
            in3 => \N__23062\,
            lcout => \c0.n3_adj_2223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_25_i3_2_lut_3_lut_4_lut_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23061\,
            in1 => \N__24682\,
            in2 => \N__22701\,
            in3 => \N__29659\,
            lcout => \c0.n3_adj_2225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11115_2_lut_3_lut_4_lut_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__33530\,
            in1 => \N__22015\,
            in2 => \N__21799\,
            in3 => \N__32790\,
            lcout => \c0.n1439\,
            ltout => \c0.n1439_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_27_i3_2_lut_3_lut_4_lut_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23063\,
            in1 => \N__22668\,
            in2 => \N__20275\,
            in3 => \N__24960\,
            lcout => \c0.n3_adj_2221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10763_2_lut_3_lut_4_lut_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23422\,
            in1 => \N__23233\,
            in2 => \N__21886\,
            in3 => \N__22971\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i7_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33195\,
            in1 => \N__32803\,
            in2 => \_gnd_net_\,
            in3 => \N__20251\,
            lcout => \c0.FRAME_MATCHER_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50417\,
            ce => 'H',
            sr => \N__20245\
        );

    \c0.select_238_Select_7_i3_2_lut_3_lut_4_lut_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22695\,
            in1 => \N__21884\,
            in2 => \N__29707\,
            in3 => \N__22979\,
            lcout => \c0.n3_adj_2250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10764_2_lut_3_lut_4_lut_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23234\,
            in1 => \N__21905\,
            in2 => \N__23042\,
            in3 => \N__23421\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_6_i3_2_lut_3_lut_4_lut_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22696\,
            in1 => \N__21906\,
            in2 => \N__29706\,
            in3 => \N__22978\,
            lcout => \c0.n3_adj_2253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_12_i3_2_lut_3_lut_4_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22975\,
            in1 => \N__29661\,
            in2 => \N__25477\,
            in3 => \N__22694\,
            lcout => \c0.n3_adj_2245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_19_i3_2_lut_3_lut_4_lut_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22693\,
            in1 => \N__21514\,
            in2 => \N__29705\,
            in3 => \N__22976\,
            lcout => \c0.n3_adj_2237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_20_i3_2_lut_3_lut_4_lut_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22977\,
            in1 => \N__29665\,
            in2 => \N__24545\,
            in3 => \N__22692\,
            lcout => \c0.n3_adj_2235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10759_2_lut_3_lut_4_lut_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23367\,
            in1 => \N__23202\,
            in2 => \N__28323\,
            in3 => \N__22915\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i11_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__32826\,
            in1 => \N__33182\,
            in2 => \_gnd_net_\,
            in3 => \N__20353\,
            lcout => \c0.FRAME_MATCHER_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50426\,
            ce => 'H',
            sr => \N__20347\
        );

    \c0.select_238_Select_11_i3_2_lut_3_lut_4_lut_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22699\,
            in1 => \N__29709\,
            in2 => \N__28324\,
            in3 => \N__22926\,
            lcout => \c0.n3_adj_2246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10760_2_lut_3_lut_4_lut_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23203\,
            in1 => \N__28185\,
            in2 => \N__22993\,
            in3 => \N__23364\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_10_i3_2_lut_3_lut_4_lut_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22697\,
            in1 => \N__29708\,
            in2 => \N__28189\,
            in3 => \N__22925\,
            lcout => \c0.n3_adj_2247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10761_2_lut_3_lut_4_lut_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23204\,
            in1 => \N__21851\,
            in2 => \N__22994\,
            in3 => \N__23365\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_9_i3_2_lut_3_lut_4_lut_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22698\,
            in1 => \N__29710\,
            in2 => \N__21856\,
            in3 => \N__22927\,
            lcout => \c0.n3_adj_2248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10762_2_lut_3_lut_4_lut_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23205\,
            in1 => \N__24860\,
            in2 => \N__22995\,
            in3 => \N__23366\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10751_2_lut_3_lut_4_lut_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23188\,
            in1 => \N__21520\,
            in2 => \N__22989\,
            in3 => \N__23378\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10750_2_lut_3_lut_4_lut_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23377\,
            in1 => \N__23187\,
            in2 => \N__24550\,
            in3 => \N__22891\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10749_2_lut_3_lut_4_lut_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23186\,
            in1 => \N__24402\,
            in2 => \N__22988\,
            in3 => \N__23376\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10747_2_lut_3_lut_4_lut_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23375\,
            in1 => \N__23185\,
            in2 => \N__24727\,
            in3 => \N__22887\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_454_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23581\,
            in1 => \N__22371\,
            in2 => \N__25294\,
            in3 => \N__22183\,
            lcout => OPEN,
            ltout => \c0.n18_adj_2198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_456_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__23494\,
            in1 => \N__20581\,
            in2 => \N__20401\,
            in3 => \N__22213\,
            lcout => \c0.n127_adj_2136\,
            ltout => \c0.n127_adj_2136_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10568_2_lut_3_lut_4_lut_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32691\,
            in1 => \N__23184\,
            in2 => \N__20521\,
            in3 => \N__22886\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10743_2_lut_3_lut_4_lut_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23370\,
            in1 => \N__23197\,
            in2 => \N__24961\,
            in3 => \N__22904\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__20563\,
            in1 => \N__33758\,
            in2 => \N__30487\,
            in3 => \N__20512\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10736_2_lut_3_lut_4_lut_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23368\,
            in1 => \N__23195\,
            in2 => \N__24913\,
            in3 => \N__22902\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10745_2_lut_3_lut_4_lut_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23199\,
            in1 => \N__24680\,
            in2 => \N__22990\,
            in3 => \N__23374\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10742_2_lut_3_lut_4_lut_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23369\,
            in1 => \N__23196\,
            in2 => \N__25018\,
            in3 => \N__22903\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10746_2_lut_3_lut_4_lut_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23200\,
            in1 => \N__21471\,
            in2 => \N__22991\,
            in3 => \N__23373\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10744_2_lut_3_lut_4_lut_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23371\,
            in1 => \N__23198\,
            in2 => \N__24823\,
            in3 => \N__22905\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10748_2_lut_3_lut_4_lut_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23201\,
            in1 => \N__24768\,
            in2 => \N__22992\,
            in3 => \N__23372\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_425_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29085\,
            in1 => \N__28977\,
            in2 => \N__23734\,
            in3 => \N__25969\,
            lcout => \c0.n9743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_698_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__23605\,
            in1 => \N__26152\,
            in2 => \N__22418\,
            in3 => \N__25860\,
            lcout => \c0.n12_adj_2200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_437_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__26151\,
            in1 => \N__22409\,
            in2 => \_gnd_net_\,
            in3 => \N__23604\,
            lcout => \c0.n9493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__7__2266_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27761\,
            in1 => \N__25861\,
            in2 => \_gnd_net_\,
            in3 => \N__23535\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__2__2255_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26901\,
            in1 => \N__27762\,
            in2 => \_gnd_net_\,
            in3 => \N__26203\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10733_2_lut_3_lut_4_lut_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23240\,
            in1 => \N__23402\,
            in2 => \N__22501\,
            in3 => \N__23016\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__4__2253_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31795\,
            in1 => \N__27763\,
            in2 => \_gnd_net_\,
            in3 => \N__22053\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_40_i8_2_lut_3_lut_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__21633\,
            in1 => \N__32704\,
            in2 => \_gnd_net_\,
            in3 => \N__25085\,
            lcout => \c0.n8_adj_2310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__20562\,
            in1 => \N__33759\,
            in2 => \N__26918\,
            in3 => \N__20646\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__20647\,
            in1 => \N__31794\,
            in2 => \N__33766\,
            in3 => \N__20535\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i16_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__31995\,
            in1 => \N__28762\,
            in2 => \N__28611\,
            in3 => \N__26525\,
            lcout => \c0.data_in_frame_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__2__2279_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27768\,
            in1 => \N__26150\,
            in2 => \_gnd_net_\,
            in3 => \N__20611\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__3__2278_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20599\,
            in1 => \N__23511\,
            in2 => \_gnd_net_\,
            in3 => \N__27769\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i9_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__28761\,
            in1 => \N__25594\,
            in2 => \N__26436\,
            in3 => \N__31997\,
            lcout => \c0.data_in_frame_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i22_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31996\,
            in1 => \N__31877\,
            in2 => \N__31229\,
            in3 => \N__26286\,
            lcout => \c0.data_in_frame_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i12_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__28760\,
            in1 => \N__30505\,
            in2 => \N__28524\,
            in3 => \N__31994\,
            lcout => \c0.data_in_frame_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i24_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__31918\,
            in1 => \N__23811\,
            in2 => \N__26537\,
            in3 => \N__31991\,
            lcout => \c0.data_in_frame_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_435_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23745\,
            in1 => \N__28393\,
            in2 => \_gnd_net_\,
            in3 => \N__28514\,
            lcout => \c0.n15939\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i17_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__31917\,
            in1 => \N__30219\,
            in2 => \N__25593\,
            in3 => \N__31990\,
            lcout => \c0.data_in_frame_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_423_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28561\,
            in2 => \_gnd_net_\,
            in3 => \N__28513\,
            lcout => \c0.n17004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__25638\,
            in1 => \N__20725\,
            in2 => \N__33765\,
            in3 => \N__20640\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_585_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__24453\,
            in1 => \N__24509\,
            in2 => \N__25140\,
            in3 => \N__23721\,
            lcout => \c0.n16891\,
            ltout => \c0.n16891_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i14_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__28785\,
            in1 => \N__31212\,
            in2 => \N__20701\,
            in3 => \N__26249\,
            lcout => \c0.data_in_frame_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i63_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20848\,
            in1 => \N__25639\,
            in2 => \_gnd_net_\,
            in3 => \N__25749\,
            lcout => data_in_frame_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i59_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26577\,
            in1 => \N__26919\,
            in2 => \_gnd_net_\,
            in3 => \N__20847\,
            lcout => data_in_frame_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i11_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__28801\,
            in1 => \N__28397\,
            in2 => \N__26932\,
            in3 => \N__31993\,
            lcout => \c0.data_in_frame_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_396_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20698\,
            in2 => \_gnd_net_\,
            in3 => \N__20662\,
            lcout => n9477,
            ltout => \n9477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__25562\,
            in1 => \N__20629\,
            in2 => \N__20614\,
            in3 => \N__33746\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i64_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20849\,
            in1 => \N__26521\,
            in2 => \_gnd_net_\,
            in3 => \N__26070\,
            lcout => data_in_frame_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i58_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30683\,
            in1 => \N__26322\,
            in2 => \_gnd_net_\,
            in3 => \N__20846\,
            lcout => data_in_frame_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i61_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31812\,
            in1 => \N__26304\,
            in2 => \_gnd_net_\,
            in3 => \N__20851\,
            lcout => data_in_frame_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i13_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21247\,
            in1 => \N__26732\,
            in2 => \_gnd_net_\,
            in3 => \N__20989\,
            lcout => \c0.delay_counter_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15371_4_lut_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24104\,
            in1 => \N__20761\,
            in2 => \N__31384\,
            in3 => \N__20809\,
            lcout => \c0.tx.n17462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i0_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20893\,
            in1 => \N__20928\,
            in2 => \_gnd_net_\,
            in3 => \N__20988\,
            lcout => \c0.delay_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__20810\,
            in1 => \N__31315\,
            in2 => \N__20764\,
            in3 => \N__20776\,
            lcout => OPEN,
            ltout => \c0.tx.n17975_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n17975_bdd_4_lut_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__20762\,
            in1 => \N__29419\,
            in2 => \N__20740\,
            in3 => \N__23833\,
            lcout => OPEN,
            ltout => \c0.tx.o_Tx_Serial_N_2064_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24067\,
            in2 => \N__20737\,
            in3 => \N__24173\,
            lcout => n3_adj_2406,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i2_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__20977\,
            in1 => \N__21178\,
            in2 => \N__26650\,
            in3 => \N__27556\,
            lcout => \c0.delay_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i10_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__21363\,
            in1 => \N__21343\,
            in2 => \N__27573\,
            in3 => \N__20976\,
            lcout => \c0.delay_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i14_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__20980\,
            in1 => \_gnd_net_\,
            in2 => \N__21199\,
            in3 => \N__21233\,
            lcout => \c0.delay_counter_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_616_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__35761\,
            in1 => \N__45924\,
            in2 => \_gnd_net_\,
            in3 => \N__24196\,
            lcout => \c0.n1419\,
            ltout => \c0.n1419_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i6_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__21076\,
            in1 => \N__21096\,
            in2 => \N__20992\,
            in3 => \N__27557\,
            lcout => \c0.delay_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i12_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21259\,
            in1 => \N__21289\,
            in2 => \_gnd_net_\,
            in3 => \N__20979\,
            lcout => \c0.delay_counter_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i8_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__20978\,
            in1 => \N__26698\,
            in2 => \N__21034\,
            in3 => \N__27558\,
            lcout => \c0.delay_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i7_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21043\,
            in1 => \N__21067\,
            in2 => \_gnd_net_\,
            in3 => \N__20981\,
            lcout => \c0.delay_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_2_lut_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__20935\,
            in1 => \N__20924\,
            in2 => \_gnd_net_\,
            in3 => \N__20884\,
            lcout => \c0.n17637\,
            ltout => OPEN,
            carryin => \bfn_5_31_0_\,
            carryout => \c0.n15514\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_3_lut_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20877\,
            in2 => \_gnd_net_\,
            in3 => \N__20854\,
            lcout => \c0.n6531\,
            ltout => OPEN,
            carryin => \c0.n15514\,
            carryout => \c0.n15515\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_4_lut_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26635\,
            in2 => \_gnd_net_\,
            in3 => \N__21172\,
            lcout => \c0.n6530\,
            ltout => OPEN,
            carryin => \c0.n15515\,
            carryout => \c0.n15516\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_5_lut_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21169\,
            in2 => \_gnd_net_\,
            in3 => \N__21145\,
            lcout => \c0.n6529\,
            ltout => OPEN,
            carryin => \c0.n15516\,
            carryout => \c0.n15517\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_6_lut_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26670\,
            in2 => \_gnd_net_\,
            in3 => \N__21133\,
            lcout => \c0.n6528\,
            ltout => OPEN,
            carryin => \c0.n15517\,
            carryout => \c0.n15518\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_7_lut_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27569\,
            in1 => \N__21128\,
            in2 => \_gnd_net_\,
            in3 => \N__21100\,
            lcout => \c0.n17574\,
            ltout => OPEN,
            carryin => \c0.n15518\,
            carryout => \c0.n15519\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_8_lut_LC_5_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21095\,
            in2 => \_gnd_net_\,
            in3 => \N__21070\,
            lcout => \c0.n6526\,
            ltout => OPEN,
            carryin => \c0.n15519\,
            carryout => \c0.n15520\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_9_lut_LC_5_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27568\,
            in1 => \N__21065\,
            in2 => \_gnd_net_\,
            in3 => \N__21037\,
            lcout => \c0.n17638\,
            ltout => OPEN,
            carryin => \c0.n15520\,
            carryout => \c0.n15521\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_10_lut_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26703\,
            in2 => \_gnd_net_\,
            in3 => \N__21022\,
            lcout => \c0.n6524\,
            ltout => OPEN,
            carryin => \bfn_5_32_0_\,
            carryout => \c0.n15522\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_11_lut_LC_5_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21018\,
            in2 => \_gnd_net_\,
            in3 => \N__20995\,
            lcout => \c0.n6523\,
            ltout => OPEN,
            carryin => \c0.n15522\,
            carryout => \c0.n15523\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_12_lut_LC_5_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21364\,
            in2 => \_gnd_net_\,
            in3 => \N__21334\,
            lcout => \c0.n6522\,
            ltout => OPEN,
            carryin => \c0.n15523\,
            carryout => \c0.n15524\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_13_lut_LC_5_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21331\,
            in2 => \_gnd_net_\,
            in3 => \N__21298\,
            lcout => \c0.n6521\,
            ltout => OPEN,
            carryin => \c0.n15524\,
            carryout => \c0.n15525\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_14_lut_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27549\,
            in1 => \_gnd_net_\,
            in2 => \N__21295\,
            in3 => \N__21250\,
            lcout => \c0.n17575\,
            ltout => OPEN,
            carryin => \c0.n15525\,
            carryout => \c0.n15526\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_15_lut_LC_5_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27548\,
            in1 => \N__26734\,
            in2 => \_gnd_net_\,
            in3 => \N__21238\,
            lcout => \c0.n17639\,
            ltout => OPEN,
            carryin => \c0.n15526\,
            carryout => \c0.n15527\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2495_16_lut_LC_5_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27550\,
            in1 => \N__21234\,
            in2 => \_gnd_net_\,
            in3 => \N__21202\,
            lcout => \c0.n17635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i29_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__34653\,
            in1 => \N__21752\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_state_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50418\,
            ce => 'H',
            sr => \N__21532\
        );

    \c0.i1_2_lut_adj_738_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29981\,
            in3 => \N__24601\,
            lcout => \c0.n16371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_703_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33402\,
            in2 => \_gnd_net_\,
            in3 => \N__29968\,
            lcout => \c0.n16331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_719_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25259\,
            in2 => \_gnd_net_\,
            in3 => \N__32590\,
            lcout => \c0.n16453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_4_lut_adj_565_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__33493\,
            in1 => \N__34281\,
            in2 => \N__32324\,
            in3 => \N__33401\,
            lcout => \c0.n8603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_760_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21754\,
            in2 => \_gnd_net_\,
            in3 => \N__29967\,
            lcout => \c0.n16381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21518\,
            in1 => \N__23485\,
            in2 => \N__21470\,
            in3 => \N__22726\,
            lcout => \c0.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i16_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111100000000"
        )
    port map (
            in0 => \N__32895\,
            in1 => \_gnd_net_\,
            in2 => \N__33097\,
            in3 => \N__21421\,
            lcout => \c0.FRAME_MATCHER_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50392\,
            ce => 'H',
            sr => \N__22576\
        );

    \c0.i1_2_lut_adj_528_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__33478\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22020\,
            lcout => n9452,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10724_3_lut_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__33517\,
            in1 => \N__23431\,
            in2 => \_gnd_net_\,
            in3 => \N__23225\,
            lcout => OPEN,
            ltout => \n1716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_765_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__21397\,
            in1 => \N__32894\,
            in2 => \N__21406\,
            in3 => \N__23043\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111111"
        )
    port map (
            in0 => \N__33053\,
            in1 => \N__28029\,
            in2 => \N__21582\,
            in3 => \N__22353\,
            lcout => n16775,
            ltout => \n16775_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_802_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110101"
        )
    port map (
            in0 => \N__21387\,
            in1 => \N__27906\,
            in2 => \N__21367\,
            in3 => \N__21672\,
            lcout => n16776,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_406_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__22019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33477\,
            lcout => n9453,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i14_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29816\,
            in2 => \_gnd_net_\,
            in3 => \N__34559\,
            lcout => \c0.FRAME_MATCHER_state_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50405\,
            ce => 'H',
            sr => \N__25426\
        );

    \c0.i10695_4_lut_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__22492\,
            in1 => \N__32669\,
            in2 => \N__21657\,
            in3 => \N__25175\,
            lcout => n2275,
            ltout => \n2275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15357_2_lut_3_lut_4_lut_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23224\,
            in1 => \N__23420\,
            in2 => \N__21559\,
            in3 => \N__23040\,
            lcout => \c0.n17454\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4944_2_lut_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23419\,
            in2 => \_gnd_net_\,
            in3 => \N__23223\,
            lcout => \c0.n7212\,
            ltout => \c0.n7212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15395_3_lut_4_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__27208\,
            in1 => \N__27943\,
            in2 => \N__21556\,
            in3 => \N__23041\,
            lcout => OPEN,
            ltout => \c0.n17452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__33531\,
            in1 => \N__22024\,
            in2 => \N__21553\,
            in3 => \N__21550\,
            lcout => \c0.n7\,
            ltout => \c0.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i5_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21544\,
            in3 => \N__21787\,
            lcout => \c0.FRAME_MATCHER_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50410\,
            ce => 'H',
            sr => \N__21541\
        );

    \c0.i1_2_lut_adj_707_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29920\,
            lcout => \c0.n16335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_467_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21785\,
            in2 => \_gnd_net_\,
            in3 => \N__21770\,
            lcout => \c0.n6_adj_2213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_458_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__25329\,
            in1 => \N__21753\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n59\,
            ltout => \c0.n59_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_476_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29775\,
            in1 => \N__33412\,
            in2 => \N__21733\,
            in3 => \N__24615\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2262_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_479_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28140\,
            in1 => \N__25366\,
            in2 => \N__21730\,
            in3 => \N__24580\,
            lcout => \c0.n16876\,
            ltout => \c0.n16876_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_415_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29509\,
            in2 => \N__21727\,
            in3 => \_gnd_net_\,
            lcout => \c0.n60\,
            ltout => \c0.n60_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14820_4_lut_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24313\,
            in1 => \N__21952\,
            in2 => \N__21724\,
            in3 => \N__32368\,
            lcout => \c0.n17258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i23_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34558\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21688\,
            lcout => \c0.FRAME_MATCHER_state_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50419\,
            ce => 'H',
            sr => \N__21721\
        );

    \c0.i1_2_lut_adj_747_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21687\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29919\,
            lcout => \c0.n16363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_635_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21711\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21686\,
            lcout => \c0.n16898\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30084\,
            in1 => \N__30025\,
            in2 => \N__32341\,
            in3 => \N__21958\,
            lcout => \c0.n9451\,
            ltout => \c0.n9451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10592_2_lut_3_lut_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27937\,
            in1 => \_gnd_net_\,
            in2 => \N__22030\,
            in3 => \N__33522\,
            lcout => n12933,
            ltout => \n12933_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10929_2_lut_3_lut_4_lut_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__22009\,
            in1 => \N__27770\,
            in2 => \N__22027\,
            in3 => \N__33534\,
            lcout => \c0.n13272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i33_3_lut_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27938\,
            in1 => \N__33523\,
            in2 => \_gnd_net_\,
            in3 => \N__22008\,
            lcout => OPEN,
            ltout => \c0.n28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_404_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__21985\,
            in1 => \N__21973\,
            in2 => \N__21967\,
            in3 => \N__32783\,
            lcout => n16795,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__29474\,
            in1 => \N__24312\,
            in2 => \_gnd_net_\,
            in3 => \N__21964\,
            lcout => \c0.n16879\,
            ltout => \c0.n16879_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_419_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33521\,
            in1 => \N__21948\,
            in2 => \N__21928\,
            in3 => \N__32367\,
            lcout => n9445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21918\,
            in1 => \N__21885\,
            in2 => \N__21847\,
            in3 => \N__22164\,
            lcout => \c0.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_422_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__21810\,
            in1 => \N__32292\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n9488\,
            ltout => \c0.n9488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_436_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__25837\,
            in1 => \N__22240\,
            in2 => \N__22228\,
            in3 => \N__22225\,
            lcout => \c0.n9485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_740_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27990\,
            in2 => \_gnd_net_\,
            in3 => \N__29893\,
            lcout => \c0.n16369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14802_2_lut_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23611\,
            lcout => \c0.n17240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__1__2280_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22426\,
            in1 => \N__27782\,
            in2 => \_gnd_net_\,
            in3 => \N__25292\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14818_4_lut_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22207\,
            in1 => \N__25925\,
            in2 => \N__25828\,
            in3 => \N__27609\,
            lcout => \c0.n17256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_410_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27608\,
            in1 => \N__22206\,
            in2 => \N__25929\,
            in3 => \N__22182\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__25824\,
            in1 => \N__25270\,
            in2 => \N__22171\,
            in3 => \N__23548\,
            lcout => \c0.n9482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10741_2_lut_3_lut_4_lut_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23354\,
            in1 => \N__22168\,
            in2 => \N__22954\,
            in3 => \N__23182\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_411_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22111\,
            in1 => \N__22081\,
            in2 => \N__22057\,
            in3 => \N__22383\,
            lcout => OPEN,
            ltout => \c0.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__22531\,
            in1 => \N__22519\,
            in2 => \N__22504\,
            in3 => \N__26208\,
            lcout => n127_adj_2418,
            ltout => \n127_adj_2418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_691_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__22495\,
            in1 => \N__25168\,
            in2 => \N__22435\,
            in3 => \N__23352\,
            lcout => n9435,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__22432\,
            in1 => \N__22425\,
            in2 => \N__22387\,
            in3 => \N__22375\,
            lcout => n127,
            ltout => \n127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_751_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22349\,
            in1 => \N__23351\,
            in2 => \N__22327\,
            in3 => \N__22856\,
            lcout => \c0.n2\,
            ltout => \c0.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__32834\,
            in1 => \N__23183\,
            in2 => \N__22312\,
            in3 => \N__22299\,
            lcout => \c0.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4924_2_lut_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23353\,
            in2 => \_gnd_net_\,
            in3 => \N__22855\,
            lcout => n7198,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10752_2_lut_3_lut_4_lut_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23357\,
            in1 => \N__23189\,
            in2 => \N__23484\,
            in3 => \N__22895\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i18_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33183\,
            in1 => \N__32835\,
            in2 => \_gnd_net_\,
            in3 => \N__22249\,
            lcout => \c0.FRAME_MATCHER_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50452\,
            ce => 'H',
            sr => \N__23449\
        );

    \c0.select_238_Select_18_i3_2_lut_3_lut_4_lut_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22708\,
            in1 => \N__23479\,
            in2 => \N__29749\,
            in3 => \N__22901\,
            lcout => \c0.n3_adj_2239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_764_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22898\,
            in1 => \_gnd_net_\,
            in2 => \N__23235\,
            in3 => \N__23358\,
            lcout => n8828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10753_2_lut_3_lut_4_lut_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23356\,
            in1 => \N__23190\,
            in2 => \N__28082\,
            in3 => \N__22896\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_17_i3_2_lut_3_lut_4_lut_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22900\,
            in1 => \N__29745\,
            in2 => \N__28083\,
            in3 => \N__22707\,
            lcout => \c0.n3_adj_2240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10754_2_lut_3_lut_4_lut_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23355\,
            in1 => \N__23191\,
            in2 => \N__22753\,
            in3 => \N__22897\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1312_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_16_i3_2_lut_3_lut_4_lut_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22899\,
            in1 => \N__29744\,
            in2 => \N__22751\,
            in3 => \N__22706\,
            lcout => \c0.n3_adj_2241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_438_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__29133\,
            in1 => \N__22564\,
            in2 => \N__22543\,
            in3 => \N__26428\,
            lcout => \c0.n21_adj_2171\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i5_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30422\,
            in1 => \N__31797\,
            in2 => \_gnd_net_\,
            in3 => \N__30339\,
            lcout => data_in_frame_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_420_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28603\,
            in2 => \_gnd_net_\,
            in3 => \N__26858\,
            lcout => \c0.n17013\,
            ltout => \c0.n17013_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_440_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23668\,
            in1 => \N__23781\,
            in2 => \N__23644\,
            in3 => \N__26253\,
            lcout => \c0.n17015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__6__2259_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23607\,
            in1 => \_gnd_net_\,
            in2 => \N__27783\,
            in3 => \N__27828\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_430_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23641\,
            in1 => \N__23782\,
            in2 => \N__23632\,
            in3 => \N__26831\,
            lcout => \c0.n17014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i3_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26910\,
            in1 => \N__25951\,
            in2 => \_gnd_net_\,
            in3 => \N__30421\,
            lcout => data_in_frame_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__6__2251_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25672\,
            in1 => \N__27764\,
            in2 => \_gnd_net_\,
            in3 => \N__23606\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14830_3_lut_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23580\,
            in1 => \N__23507\,
            in2 => \_gnd_net_\,
            in3 => \N__23530\,
            lcout => \c0.n17268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i82_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__31111\,
            in1 => \N__30697\,
            in2 => \N__23797\,
            in3 => \N__31878\,
            lcout => \c0.data_in_frame_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i87_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__31879\,
            in1 => \N__23764\,
            in2 => \N__25675\,
            in3 => \N__31112\,
            lcout => \c0.data_in_frame_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23531\,
            in1 => \N__25887\,
            in2 => \N__23512\,
            in3 => \N__26173\,
            lcout => \c0.n19_adj_2199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i79_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__28763\,
            in1 => \N__23680\,
            in2 => \N__25674\,
            in3 => \N__31110\,
            lcout => \c0.data_in_frame_9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_427_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26241\,
            in1 => \N__26832\,
            in2 => \N__23796\,
            in3 => \N__23780\,
            lcout => OPEN,
            ltout => \c0.n16954_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_439_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30575\,
            in2 => \N__23767\,
            in3 => \N__23691\,
            lcout => OPEN,
            ltout => \c0.n18_adj_2174_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_455_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111111"
        )
    port map (
            in0 => \N__23763\,
            in1 => \N__30271\,
            in2 => \N__23755\,
            in3 => \N__23752\,
            lcout => \c0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i77_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31109\,
            in1 => \N__28799\,
            in2 => \N__31826\,
            in3 => \N__23746\,
            lcout => \c0.data_in_frame_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_421_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28392\,
            in1 => \N__29114\,
            in2 => \_gnd_net_\,
            in3 => \N__29049\,
            lcout => \c0.n6_adj_2152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_666_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__24454\,
            in1 => \N__24510\,
            in2 => \N__25144\,
            in3 => \N__23722\,
            lcout => \c0.n16882\,
            ltout => \c0.n16882_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i85_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__31919\,
            in1 => \N__31819\,
            in2 => \N__23695\,
            in3 => \N__23692\,
            lcout => \c0.data_in_frame_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_429_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23679\,
            in1 => \N__26242\,
            in2 => \_gnd_net_\,
            in3 => \N__28575\,
            lcout => \c0.n15938\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i73_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__28796\,
            in1 => \N__28992\,
            in2 => \N__25595\,
            in3 => \N__31107\,
            lcout => \c0.data_in_frame_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i10_LC_6_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__29115\,
            in1 => \N__28798\,
            in2 => \N__30693\,
            in3 => \N__31992\,
            lcout => \c0.data_in_frame_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i76_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__28797\,
            in1 => \N__28356\,
            in2 => \N__30531\,
            in3 => \N__31108\,
            lcout => \c0.data_in_frame_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i15_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__28800\,
            in1 => \N__25649\,
            in2 => \N__26833\,
            in3 => \N__31998\,
            lcout => \c0.data_in_frame_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_adj_566_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__26820\,
            in1 => \N__29036\,
            in2 => \N__23812\,
            in3 => \N__30300\,
            lcout => \c0.n22_adj_2301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i88_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__31923\,
            in1 => \N__28467\,
            in2 => \N__26538\,
            in3 => \N__31114\,
            lcout => \c0.data_in_frame_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i20_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32000\,
            in1 => \N__31921\,
            in2 => \N__30532\,
            in3 => \N__26271\,
            lcout => \c0.data_in_frame_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i49_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28872\,
            in1 => \N__25563\,
            in2 => \_gnd_net_\,
            in3 => \N__25735\,
            lcout => data_in_frame_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i23_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32001\,
            in1 => \N__31922\,
            in2 => \N__25665\,
            in3 => \N__30237\,
            lcout => \c0.data_in_frame_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i19_LC_6_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31999\,
            in1 => \N__31920\,
            in2 => \N__26940\,
            in3 => \N__26349\,
            lcout => \c0.data_in_frame_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i7_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25664\,
            in1 => \N__29045\,
            in2 => \_gnd_net_\,
            in3 => \N__30441\,
            lcout => data_in_frame_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23824\,
            in2 => \_gnd_net_\,
            in3 => \N__31642\,
            lcout => \c0.n65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i43_4_lut_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__46395\,
            in1 => \N__26755\,
            in2 => \N__42749\,
            in3 => \N__24301\,
            lcout => \c0.n25_adj_2324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15400_3_lut_4_lut_4_lut_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010110000000"
        )
    port map (
            in0 => \N__24182\,
            in1 => \N__24113\,
            in2 => \N__24075\,
            in3 => \N__31736\,
            lcout => OPEN,
            ltout => \n4_adj_2458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111010"
        )
    port map (
            in0 => \N__31643\,
            in1 => \N__24074\,
            in2 => \N__24190\,
            in3 => \N__23878\,
            lcout => tx_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24183\,
            in1 => \N__24114\,
            in2 => \N__24076\,
            in3 => \N__23877\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14957_3_lut_LC_6_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26745\,
            in1 => \N__32083\,
            in2 => \_gnd_net_\,
            in3 => \N__31378\,
            lcout => n17395,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_prev_2155_LC_6_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31644\,
            lcout => \c0.tx_active_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2494_2_lut_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23818\,
            in2 => \N__51887\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_transmit_N_1949_0\,
            ltout => OPEN,
            carryin => \bfn_6_30_0_\,
            carryout => \c0.n15653\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2494_3_lut_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52175\,
            in2 => \_gnd_net_\,
            in3 => \N__24217\,
            lcout => \c0.tx_transmit_N_1949_1\,
            ltout => OPEN,
            carryin => \c0.n15653\,
            carryout => \c0.n15654\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2494_4_lut_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52351\,
            in2 => \_gnd_net_\,
            in3 => \N__24214\,
            lcout => \c0.tx_transmit_N_1949_2\,
            ltout => OPEN,
            carryin => \c0.n15654\,
            carryout => \c0.n15655\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2494_5_lut_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43078\,
            in2 => \_gnd_net_\,
            in3 => \N__24211\,
            lcout => \c0.tx_transmit_N_1949_3\,
            ltout => OPEN,
            carryin => \c0.n15655\,
            carryout => \c0.n15656\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2494_6_lut_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35471\,
            in2 => \_gnd_net_\,
            in3 => \N__24208\,
            lcout => \c0.tx_transmit_N_1949_4\,
            ltout => OPEN,
            carryin => \c0.n15656\,
            carryout => \c0.n15657\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2494_7_lut_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26596\,
            in3 => \N__24205\,
            lcout => \c0.tx_transmit_N_1949_5\,
            ltout => OPEN,
            carryin => \c0.n15657\,
            carryout => \c0.n15658\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2494_8_lut_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27012\,
            in2 => \_gnd_net_\,
            in3 => \N__24202\,
            lcout => \c0.tx_transmit_N_1949_6\,
            ltout => OPEN,
            carryin => \c0.n15658\,
            carryout => \c0.n15659\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2494_9_lut_LC_6_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27105\,
            in2 => \_gnd_net_\,
            in3 => \N__24199\,
            lcout => \c0.tx_transmit_N_1949_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i1_LC_6_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__24238\,
            in1 => \N__35745\,
            in2 => \N__52236\,
            in3 => \N__27145\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50526\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i152_2_lut_4_lut_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__27171\,
            in1 => \N__27189\,
            in2 => \N__31737\,
            in3 => \N__31660\,
            lcout => \c0.n456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__26957\,
            in1 => \N__27026\,
            in2 => \_gnd_net_\,
            in3 => \N__27039\,
            lcout => \c0.n8938\,
            ltout => \c0.n8938_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_677_LC_6_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__27170\,
            in1 => \N__27338\,
            in2 => \N__24253\,
            in3 => \N__27308\,
            lcout => \c0.n22_adj_2164\,
            ltout => \c0.n22_adj_2164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_4_lut_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__42574\,
            in1 => \N__46415\,
            in2 => \N__24241\,
            in3 => \N__27385\,
            lcout => \c0.n42_adj_2165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_604_LC_6_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__26973\,
            in1 => \N__24237\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n4_adj_2311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15441_2_lut_3_lut_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__42575\,
            in1 => \_gnd_net_\,
            in2 => \N__45848\,
            in3 => \N__46416\,
            lcout => \data_out_10__7__N_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6219_4_lut_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101100"
        )
    port map (
            in0 => \N__24283\,
            in1 => \N__24300\,
            in2 => \N__42645\,
            in3 => \N__45761\,
            lcout => \c0.n8631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_697_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__46302\,
            in1 => \N__34309\,
            in2 => \N__45549\,
            in3 => \N__27427\,
            lcout => OPEN,
            ltout => \c0.n15868_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_701_LC_6_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__27576\,
            in1 => \N__46303\,
            in2 => \N__24229\,
            in3 => \N__24226\,
            lcout => OPEN,
            ltout => \n10141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state_i0_i1_LC_6_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000001010"
        )
    port map (
            in0 => \N__46304\,
            in1 => \_gnd_net_\,
            in2 => \N__24220\,
            in3 => \N__45907\,
            lcout => \UART_TRANSMITTER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14724_2_lut_LC_6_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__34310\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46301\,
            lcout => n17162,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__6__2214_LC_6_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__46305\,
            in1 => \N__34053\,
            in2 => \N__46150\,
            in3 => \N__42580\,
            lcout => \c0.data_out_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i142_2_lut_4_lut_LC_6_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__27357\,
            in1 => \N__27310\,
            in2 => \N__27464\,
            in3 => \N__27375\,
            lcout => \c0.n446\,
            ltout => \c0.n446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15401_4_lut_LC_6_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__45760\,
            in1 => \N__42576\,
            in2 => \N__24286\,
            in3 => \N__24282\,
            lcout => n10031,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i19_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24602\,
            in2 => \_gnd_net_\,
            in3 => \N__34654\,
            lcout => \c0.FRAME_MATCHER_state_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50420\,
            ce => 'H',
            sr => \N__24274\
        );

    \c0.FRAME_MATCHER_state_i10_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25260\,
            in2 => \_gnd_net_\,
            in3 => \N__34644\,
            lcout => \c0.FRAME_MATCHER_state_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50399\,
            ce => 'H',
            sr => \N__24262\
        );

    \c0.FRAME_MATCHER_state_i21_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25412\,
            in2 => \_gnd_net_\,
            in3 => \N__34562\,
            lcout => \c0.FRAME_MATCHER_state_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50411\,
            ce => 'H',
            sr => \N__25387\
        );

    \c0.FRAME_MATCHER_state_i22_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25515\,
            in2 => \_gnd_net_\,
            in3 => \N__34560\,
            lcout => \c0.FRAME_MATCHER_state_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50421\,
            ce => 'H',
            sr => \N__25498\
        );

    \c0.i4_4_lut_adj_649_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28141\,
            in1 => \N__25374\,
            in2 => \N__29536\,
            in3 => \N__24604\,
            lcout => \c0.n10_adj_2336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_466_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25408\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25514\,
            lcout => OPEN,
            ltout => \c0.n61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_443_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24637\,
            in1 => \N__27991\,
            in2 => \N__24628\,
            in3 => \N__27880\,
            lcout => OPEN,
            ltout => \c0.n16133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_650_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24625\,
            in1 => \N__32403\,
            in2 => \N__24619\,
            in3 => \N__24616\,
            lcout => \c0.n62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_695_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24603\,
            in1 => \N__25513\,
            in2 => \N__25413\,
            in3 => \N__29809\,
            lcout => \c0.n52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_732_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32404\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29945\,
            lcout => \c0.n16347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i26_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25373\,
            in2 => \_gnd_net_\,
            in3 => \N__34563\,
            lcout => \c0.FRAME_MATCHER_state_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50427\,
            ce => 'H',
            sr => \N__25345\
        );

    \c0.FRAME_MATCHER_i_i4_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33247\,
            in1 => \N__32802\,
            in2 => \_gnd_net_\,
            in3 => \N__24574\,
            lcout => \c0.FRAME_MATCHER_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50435\,
            ce => 'H',
            sr => \N__24562\
        );

    \c0.i1_2_lut_adj_408_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__24535\,
            in1 => \N__24475\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24446\,
            in1 => \N__24398\,
            in2 => \N__24352\,
            in3 => \N__24348\,
            lcout => \c0.n51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_441_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27983\,
            in1 => \N__27879\,
            in2 => \N__30064\,
            in3 => \N__25231\,
            lcout => \c0.n56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_468_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25261\,
            in1 => \N__32614\,
            in2 => \N__34441\,
            in3 => \N__25240\,
            lcout => \c0.n16869\,
            ltout => \c0.n16869_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_471_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25225\,
            in3 => \N__30028\,
            lcout => \c0.n16871\,
            ltout => \c0.n16871_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_496_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__29532\,
            in1 => \N__32310\,
            in2 => \N__25222\,
            in3 => \N__25219\,
            lcout => \c0.n12_adj_2189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28213\,
            in1 => \N__24643\,
            in2 => \N__25213\,
            in3 => \N__24778\,
            lcout => OPEN,
            ltout => \c0.n56_adj_2146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24967\,
            in1 => \N__25204\,
            in2 => \N__25189\,
            in3 => \N__25186\,
            lcout => \c0.n9346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25121\,
            in1 => \N__25087\,
            in2 => \N__25016\,
            in3 => \N__25451\,
            lcout => \c0.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_407_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24956\,
            in1 => \N__24909\,
            in2 => \N__24864\,
            in3 => \N__24808\,
            lcout => \c0.n47_adj_2144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24751\,
            in1 => \N__24712\,
            in2 => \N__28084\,
            in3 => \N__24681\,
            lcout => \c0.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_744_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25519\,
            in2 => \_gnd_net_\,
            in3 => \N__29894\,
            lcout => \c0.n16365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i12_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33209\,
            in1 => \N__32847\,
            in2 => \_gnd_net_\,
            in3 => \N__25486\,
            lcout => \c0.FRAME_MATCHER_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50453\,
            ce => 'H',
            sr => \N__25438\
        );

    \c0.i1_2_lut_adj_728_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29824\,
            in2 => \_gnd_net_\,
            in3 => \N__29884\,
            lcout => \c0.n16351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_742_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25414\,
            in2 => \_gnd_net_\,
            in3 => \N__29885\,
            lcout => \c0.n16367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_752_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29917\,
            in3 => \N__28139\,
            lcout => \c0.n16359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_754_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25375\,
            in2 => \_gnd_net_\,
            in3 => \N__29889\,
            lcout => \c0.n16357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_756_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29918\,
            in3 => \N__25333\,
            lcout => \c0.n16355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14828_4_lut_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25293\,
            in1 => \N__26176\,
            in2 => \N__25886\,
            in3 => \N__25850\,
            lcout => \c0.n17266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i50_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30696\,
            in1 => \N__26035\,
            in2 => \_gnd_net_\,
            in3 => \N__25724\,
            lcout => data_in_frame_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__5__2260_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25879\,
            in1 => \N__27803\,
            in2 => \_gnd_net_\,
            in3 => \N__25930\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__7__2258_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25851\,
            in1 => \_gnd_net_\,
            in2 => \N__27808\,
            in3 => \N__25818\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_432_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25790\,
            in2 => \_gnd_net_\,
            in3 => \N__27824\,
            lcout => \c0.n8_adj_2157\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__7__2250_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27802\,
            in1 => \N__26520\,
            in2 => \_gnd_net_\,
            in3 => \N__25817\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__3__2254_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25794\,
            in1 => \N__27804\,
            in2 => \_gnd_net_\,
            in3 => \N__30488\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_412_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__30267\,
            in1 => \N__25774\,
            in2 => \N__25756\,
            in3 => \N__30191\,
            lcout => \c0.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1028_2_lut_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__30377\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25950\,
            lcout => \c0.n2334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i55_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25731\,
            in1 => \N__25673\,
            in2 => \_gnd_net_\,
            in3 => \N__26091\,
            lcout => data_in_frame_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i1_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26852\,
            in1 => \N__25603\,
            in2 => \_gnd_net_\,
            in3 => \N__30436\,
            lcout => data_in_frame_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i2_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30437\,
            in1 => \N__30695\,
            in2 => \_gnd_net_\,
            in3 => \N__26780\,
            lcout => data_in_frame_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_746_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29055\,
            in1 => \N__28649\,
            in2 => \_gnd_net_\,
            in3 => \N__25962\,
            lcout => \c0.n2351\,
            ltout => \c0.n2351_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1046_2_lut_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26056\,
            in3 => \N__26851\,
            lcout => \c0.n2352\,
            ltout => \c0.n2352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011111101101"
        )
    port map (
            in0 => \N__26053\,
            in1 => \N__26034\,
            in2 => \N__26023\,
            in3 => \N__28650\,
            lcout => \c0.n23_adj_2145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__26020\,
            in1 => \N__26545\,
            in2 => \N__26002\,
            in3 => \N__25978\,
            lcout => \c0.n30_adj_2148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i137_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48769\,
            in1 => \N__34785\,
            in2 => \_gnd_net_\,
            in3 => \N__51249\,
            lcout => data_out_frame2_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_416_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25948\,
            in2 => \_gnd_net_\,
            in3 => \N__26773\,
            lcout => \c0.n9541\,
            ltout => \c0.n9541_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_414_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30334\,
            in1 => \N__30378\,
            in2 => \N__25972\,
            in3 => \N__30299\,
            lcout => \c0.n16943\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_715_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28610\,
            in1 => \N__25949\,
            in2 => \N__26109\,
            in3 => \N__26774\,
            lcout => \c0.n15929\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1030_2_lut_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__30335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30379\,
            lcout => \c0.n2336\,
            ltout => \c0.n2336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_655_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__26287\,
            in1 => \N__26272\,
            in2 => \N__26257\,
            in3 => \N__28887\,
            lcout => OPEN,
            ltout => \c0.n20_adj_2340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_659_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110111"
        )
    port map (
            in0 => \N__26254\,
            in1 => \N__28827\,
            in2 => \N__26215\,
            in3 => \N__26435\,
            lcout => \c0.n26_adj_2344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15345_2_lut_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40243\,
            in2 => \_gnd_net_\,
            in3 => \N__51938\,
            lcout => \c0.n17548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1036_2_lut_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28645\,
            in2 => \_gnd_net_\,
            in3 => \N__29050\,
            lcout => \c0.n2342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__2__2263_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26174\,
            in1 => \N__27742\,
            in2 => \_gnd_net_\,
            in3 => \N__26212\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__2__2271_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27741\,
            in1 => \N__26131\,
            in2 => \_gnd_net_\,
            in3 => \N__26175\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i84_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__31925\,
            in1 => \N__30512\,
            in2 => \N__26110\,
            in3 => \N__31113\,
            lcout => \c0.data_in_frame_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_adj_716_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__26092\,
            in1 => \N__29051\,
            in2 => \N__26077\,
            in3 => \N__30304\,
            lcout => OPEN,
            ltout => \c0.n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111011"
        )
    port map (
            in0 => \N__26581\,
            in1 => \N__26563\,
            in2 => \N__26548\,
            in3 => \N__26356\,
            lcout => \c0.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i6_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31221\,
            in1 => \N__30305\,
            in2 => \_gnd_net_\,
            in3 => \N__30434\,
            lcout => data_in_frame_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i8_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28644\,
            in1 => \_gnd_net_\,
            in2 => \N__26536\,
            in3 => \N__30435\,
            lcout => data_in_frame_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_413_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26437\,
            in2 => \_gnd_net_\,
            in3 => \N__28643\,
            lcout => \c0.n17001\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i6_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26378\,
            in1 => \N__31550\,
            in2 => \_gnd_net_\,
            in3 => \N__26401\,
            lcout => \r_Clock_Count_6_adj_2448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_417_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26781\,
            lcout => \c0.n9585\,
            ltout => \c0.n9585_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_657_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011111111"
        )
    port map (
            in0 => \N__26350\,
            in1 => \N__26335\,
            in2 => \N__26329\,
            in3 => \N__28398\,
            lcout => \c0.n27_adj_2342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111001111101"
        )
    port map (
            in0 => \N__26326\,
            in1 => \N__30580\,
            in2 => \N__26308\,
            in3 => \N__30556\,
            lcout => \c0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i83_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31115\,
            in1 => \N__31933\,
            in2 => \N__26941\,
            in3 => \N__26793\,
            lcout => \c0.data_in_frame_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_702_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26860\,
            in1 => \N__26824\,
            in2 => \N__26794\,
            in3 => \N__26782\,
            lcout => \c0.n15930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15216_3_lut_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__27471\,
            in1 => \N__27073\,
            in2 => \_gnd_net_\,
            in3 => \N__27193\,
            lcout => \c0.n17460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__26749\,
            in1 => \N__43039\,
            in2 => \N__35617\,
            in3 => \N__35511\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14798_2_lut_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26733\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26704\,
            lcout => \c0.n17236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_2_lut_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38106\,
            in2 => \_gnd_net_\,
            in3 => \N__42403\,
            lcout => \c0.n9530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i150_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41470\,
            in1 => \N__30897\,
            in2 => \_gnd_net_\,
            in3 => \N__51271\,
            lcout => data_out_frame2_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_581_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__26674\,
            in1 => \N__26645\,
            in2 => \N__26614\,
            in3 => \N__26602\,
            lcout => \c0.n23_adj_2309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i5_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__27147\,
            in1 => \N__35763\,
            in2 => \N__27052\,
            in3 => \N__26595\,
            lcout => \c0.byte_transmit_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14816_3_lut_4_lut_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__27309\,
            in1 => \N__27347\,
            in2 => \N__46399\,
            in3 => \N__27172\,
            lcout => \c0.n17254\,
            ltout => \c0.n17254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14852_3_lut_4_lut_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26958\,
            in1 => \N__27027\,
            in2 => \N__27067\,
            in3 => \N__27040\,
            lcout => \c0.n17290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i2_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__35762\,
            in1 => \N__27348\,
            in2 => \N__52437\,
            in3 => \N__27146\,
            lcout => byte_transmit_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_610_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27048\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27117\,
            lcout => \c0.n5_adj_2319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i6_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__27028\,
            in1 => \N__27013\,
            in2 => \N__35772\,
            in3 => \N__27148\,
            lcout => \c0.byte_transmit_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__6__2238_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__32055\,
            in1 => \N__42644\,
            in2 => \N__46149\,
            in3 => \N__46321\,
            lcout => \c0.data_out_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_582_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__27001\,
            in1 => \N__26995\,
            in2 => \N__31608\,
            in3 => \N__26986\,
            lcout => \c0.n16839\,
            ltout => \c0.n16839_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i0_LC_7_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__35767\,
            in1 => \N__26974\,
            in2 => \N__26962\,
            in3 => \N__51972\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i4_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__35490\,
            in1 => \N__26959\,
            in2 => \N__35760\,
            in3 => \N__27143\,
            lcout => byte_transmit_counter_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11084_2_lut_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27168\,
            in2 => \_gnd_net_\,
            in3 => \N__27188\,
            lcout => n9357,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i3_LC_7_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__27169\,
            in1 => \N__35768\,
            in2 => \N__43139\,
            in3 => \N__27142\,
            lcout => byte_transmit_counter_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i7_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__27144\,
            in1 => \N__27106\,
            in2 => \N__35773\,
            in3 => \N__27118\,
            lcout => \c0.byte_transmit_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15393_3_lut_4_lut_LC_7_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__42646\,
            in1 => \N__46306\,
            in2 => \N__45928\,
            in3 => \N__27577\,
            lcout => OPEN,
            ltout => \n17834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state_i0_i0_LC_7_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__45844\,
            in1 => \N__45548\,
            in2 => \N__27094\,
            in3 => \N__27091\,
            lcout => \UART_TRANSMITTER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state_i0_i2_LC_7_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__34291\,
            in1 => \N__27079\,
            in2 => \N__42623\,
            in3 => \N__27391\,
            lcout => \UART_TRANSMITTER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50547\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_692_LC_7_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__27377\,
            in1 => \N__27353\,
            in2 => \_gnd_net_\,
            in3 => \N__27312\,
            lcout => OPEN,
            ltout => \n9358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_792_LC_7_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__27574\,
            in1 => \N__31601\,
            in2 => \N__27085\,
            in3 => \N__27426\,
            lcout => OPEN,
            ltout => \n41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_4_lut_LC_7_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__45905\,
            in1 => \N__46299\,
            in2 => \N__27082\,
            in3 => \N__34317\,
            lcout => n35,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15262_4_lut_LC_7_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__27575\,
            in1 => \N__27378\,
            in2 => \N__27475\,
            in3 => \N__27425\,
            lcout => OPEN,
            ltout => \n17479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i57_4_lut_LC_7_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__45906\,
            in1 => \N__46300\,
            in2 => \N__27412\,
            in3 => \N__27409\,
            lcout => n38,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_690_LC_7_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__27352\,
            in1 => \N__27311\,
            in2 => \N__42622\,
            in3 => \N__27376\,
            lcout => \c0.n44_adj_2163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15277_3_lut_4_lut_LC_7_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__27379\,
            in1 => \N__46298\,
            in2 => \N__27358\,
            in3 => \N__27313\,
            lcout => \c0.n17475\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15437_2_lut_3_lut_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__27268\,
            in1 => \N__30604\,
            in2 => \_gnd_net_\,
            in3 => \N__27230\,
            lcout => \c0.tx2_transmit_N_1997\,
            ltout => \c0.tx2_transmit_N_1997_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_2249_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011101110"
        )
    port map (
            in0 => \N__32317\,
            in1 => \N__33516\,
            in2 => \N__27271\,
            in3 => \N__34275\,
            lcout => \c0.r_SM_Main_2_N_2036_0_adj_2261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50412\,
            ce => 'H',
            sr => \N__33580\
        );

    \c0.tx2.i3_4_lut_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32203\,
            in1 => \N__34756\,
            in2 => \N__34735\,
            in3 => \N__34708\,
            lcout => \c0.tx2.n113\,
            ltout => \c0.tx2.n113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_3_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30603\,
            in2 => \N__27262\,
            in3 => \N__27229\,
            lcout => n491,
            ltout => \n491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33515\,
            in2 => \N__27196\,
            in3 => \N__27939\,
            lcout => n17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i20_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27981\,
            in2 => \_gnd_net_\,
            in3 => \N__34648\,
            lcout => \c0.FRAME_MATCHER_state_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50428\,
            ce => 'H',
            sr => \N__28012\
        );

    \c0.FRAME_MATCHER_state_i24_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29473\,
            in2 => \_gnd_net_\,
            in3 => \N__34613\,
            lcout => \c0.FRAME_MATCHER_state_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50436\,
            ce => 'H',
            sr => \N__29434\
        );

    \c0.FRAME_MATCHER_state_i18_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34645\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27878\,
            lcout => \c0.FRAME_MATCHER_state_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50442\,
            ce => 'H',
            sr => \N__27841\
        );

    \c0.i6_3_lut_4_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28000\,
            in1 => \N__27982\,
            in2 => \N__30088\,
            in3 => \N__27864\,
            lcout => n9460,
            ltout => \n9460_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_519_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27910\,
            in3 => \N__33535\,
            lcout => n9462,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i64_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51224\,
            in1 => \N__44944\,
            in2 => \_gnd_net_\,
            in3 => \N__41318\,
            lcout => data_out_frame2_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50454\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_736_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29954\,
            lcout => \c0.n16343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__6__2267_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27835\,
            in1 => \N__27596\,
            in2 => \_gnd_net_\,
            in3 => \N__27790\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50454\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3112_3_lut_4_lut_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33320\,
            in1 => \N__33352\,
            in2 => \N__28342\,
            in3 => \N__32318\,
            lcout => \c0.n5543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28321\,
            in1 => \N__28291\,
            in2 => \N__28258\,
            in3 => \N__28169\,
            lcout => \c0.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i10_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33276\,
            in1 => \N__32918\,
            in2 => \_gnd_net_\,
            in3 => \N__28204\,
            lcout => \c0.FRAME_MATCHER_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50464\,
            ce => 'H',
            sr => \N__28156\
        );

    \c0.i1_2_lut_4_lut_adj_665_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40905\,
            in1 => \N__35232\,
            in2 => \N__43909\,
            in3 => \N__48882\,
            lcout => \c0.n6_adj_2293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_520_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__48883\,
            in1 => \_gnd_net_\,
            in2 => \N__35239\,
            in3 => \N__43906\,
            lcout => OPEN,
            ltout => \c0.n9819_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_449_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37021\,
            in1 => \N__49633\,
            in2 => \N__28144\,
            in3 => \N__43585\,
            lcout => \c0.n17_adj_2193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15294_2_lut_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40904\,
            in2 => \_gnd_net_\,
            in3 => \N__48211\,
            lcout => \c0.n17560\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i25_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34646\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28132\,
            lcout => \c0.FRAME_MATCHER_state_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50476\,
            ce => 'H',
            sr => \N__28102\
        );

    \c0.FRAME_MATCHER_i_i17_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33277\,
            in1 => \N__32988\,
            in2 => \_gnd_net_\,
            in3 => \N__28093\,
            lcout => \c0.FRAME_MATCHER_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50489\,
            ce => 'H',
            sr => \N__28666\
        );

    \c0.i7_4_lut_adj_656_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001101111"
        )
    port map (
            in0 => \N__29132\,
            in1 => \N__28654\,
            in2 => \N__28615\,
            in3 => \N__30192\,
            lcout => OPEN,
            ltout => \c0.n23_adj_2341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_660_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__28579\,
            in1 => \N__28540\,
            in2 => \N__28528\,
            in3 => \N__28525\,
            lcout => \c0.n30_adj_2345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_452_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111101111"
        )
    port map (
            in0 => \N__28495\,
            in1 => \N__29005\,
            in2 => \N__28486\,
            in3 => \N__28471\,
            lcout => \c0.n27_adj_2196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14914_3_lut_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__40900\,
            in1 => \N__37478\,
            in2 => \_gnd_net_\,
            in3 => \N__35018\,
            lcout => OPEN,
            ltout => \c0.n17352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i1_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__37479\,
            in1 => \N__34956\,
            in2 => \N__28453\,
            in3 => \N__37548\,
            lcout => \c0.data_out_frame2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_460_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28420\,
            in1 => \N__29062\,
            in2 => \N__28450\,
            in3 => \N__28441\,
            lcout => \c0.n15846\,
            ltout => \c0.n15846_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14903_3_lut_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37472\,
            in2 => \N__28432\,
            in3 => \N__37382\,
            lcout => \c0.n17769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_442_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111011"
        )
    port map (
            in0 => \N__28938\,
            in1 => \N__28429\,
            in2 => \N__31057\,
            in3 => \N__28960\,
            lcout => \c0.n26_adj_2184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_431_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__28414\,
            in1 => \N__28402\,
            in2 => \N__28363\,
            in3 => \N__29137\,
            lcout => OPEN,
            ltout => \c0.n23_adj_2156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111011"
        )
    port map (
            in0 => \N__28815\,
            in1 => \N__29101\,
            in2 => \N__29089\,
            in3 => \N__29086\,
            lcout => \c0.n28_adj_2183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1034_2_lut_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29056\,
            in2 => \_gnd_net_\,
            in3 => \N__30316\,
            lcout => \c0.n2340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_434_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__28704\,
            in1 => \N__28833\,
            in2 => \N__28996\,
            in3 => \N__28978\,
            lcout => \c0.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_409_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__28954\,
            in1 => \N__28939\,
            in2 => \N__28918\,
            in3 => \N__28894\,
            lcout => OPEN,
            ltout => \c0.n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110111"
        )
    port map (
            in0 => \N__28876\,
            in1 => \N__28858\,
            in2 => \N__28837\,
            in3 => \N__28834\,
            lcout => \c0.n26_adj_2147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i74_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__30679\,
            in1 => \N__28816\,
            in2 => \N__28804\,
            in3 => \N__31133\,
            lcout => \c0.data_in_frame_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i78_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31134\,
            in1 => \N__28795\,
            in2 => \N__31231\,
            in3 => \N__28705\,
            lcout => \c0.data_in_frame_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_45_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28677\,
            in1 => \N__31545\,
            in2 => \_gnd_net_\,
            in3 => \N__29275\,
            lcout => tx2_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14905_3_lut_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__35853\,
            in1 => \_gnd_net_\,
            in2 => \N__37483\,
            in3 => \N__35004\,
            lcout => \c0.n17343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i1_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001000000000"
        )
    port map (
            in0 => \N__35343\,
            in1 => \N__29184\,
            in2 => \N__35391\,
            in3 => \N__29193\,
            lcout => \r_Bit_Index_1_adj_2456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i2_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101000000000"
        )
    port map (
            in0 => \N__29256\,
            in1 => \N__29185\,
            in2 => \N__29266\,
            in3 => \N__29194\,
            lcout => \r_Bit_Index_2_adj_2455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n17903_bdd_4_lut_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__35101\,
            in1 => \N__35381\,
            in2 => \N__51484\,
            in3 => \N__35314\,
            lcout => \c0.tx2.n17906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__36793\,
            in1 => \N__35342\,
            in2 => \N__35390\,
            in3 => \N__32509\,
            lcout => OPEN,
            ltout => \c0.tx2.n18113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n18113_bdd_4_lut_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__34822\,
            in1 => \N__33949\,
            in2 => \N__29197\,
            in3 => \N__35380\,
            lcout => \c0.tx2.n18116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i14834_3_lut_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__29232\,
            in1 => \N__31027\,
            in2 => \_gnd_net_\,
            in3 => \N__29182\,
            lcout => n10398,
            ltout => \n10398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i0_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__29183\,
            in1 => \_gnd_net_\,
            in2 => \N__29155\,
            in3 => \N__35349\,
            lcout => \r_Bit_Index_0_adj_2457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i11207211_i1_3_lut_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29152\,
            in1 => \N__29146\,
            in2 => \_gnd_net_\,
            in3 => \N__29255\,
            lcout => OPEN,
            ltout => \c0.tx2.o_Tx_Serial_N_2064_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31026\,
            in2 => \N__29347\,
            in3 => \N__29340\,
            lcout => n3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2595_2_lut_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35386\,
            lcout => n5029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_3_lut_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__35385\,
            in1 => \_gnd_net_\,
            in2 => \N__29257\,
            in3 => \N__35347\,
            lcout => \c0.tx2.n13281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42968\,
            in1 => \N__47138\,
            in2 => \_gnd_net_\,
            in3 => \N__52043\,
            lcout => \c0.n8_adj_2160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52044\,
            in1 => \N__34075\,
            in2 => \_gnd_net_\,
            in3 => \N__33976\,
            lcout => OPEN,
            ltout => \c0.n2_adj_2266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18095_bdd_4_lut_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__41911\,
            in1 => \N__52150\,
            in2 => \N__29221\,
            in3 => \N__52408\,
            lcout => OPEN,
            ltout => \c0.n18098_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__52409\,
            in1 => \N__31564\,
            in2 => \N__29218\,
            in3 => \N__43150\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2139_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__29428\,
            in1 => \N__35604\,
            in2 => \N__29215\,
            in3 => \N__35518\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29212\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14956_3_lut_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29391\,
            in1 => \N__29427\,
            in2 => \_gnd_net_\,
            in3 => \N__31379\,
            lcout => n17394,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__7__2213_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__45515\,
            in1 => \N__32098\,
            in2 => \N__45929\,
            in3 => \N__46422\,
            lcout => data_out_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__29407\,
            in1 => \N__52232\,
            in2 => \N__47101\,
            in3 => \N__51970\,
            lcout => n10_adj_2426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i30_4_lut_LC_9_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51971\,
            in1 => \N__35653\,
            in2 => \N__52264\,
            in3 => \N__46756\,
            lcout => OPEN,
            ltout => \c0.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i31_4_lut_LC_9_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__32158\,
            in1 => \N__43120\,
            in2 => \N__29398\,
            in3 => \N__52460\,
            lcout => OPEN,
            ltout => \c0.n12_adj_2150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__35521\,
            in1 => \N__29392\,
            in2 => \N__29395\,
            in3 => \N__35564\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_9_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__52459\,
            in1 => \N__29557\,
            in2 => \N__29380\,
            in3 => \N__43151\,
            lcout => OPEN,
            ltout => \n10_adj_2407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_9_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__35522\,
            in1 => \N__35603\,
            in2 => \N__29371\,
            in3 => \N__29361\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15288_2_lut_LC_9_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__51997\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32478\,
            lcout => OPEN,
            ltout => \c0.n17590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18023_bdd_4_lut_LC_9_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__42898\,
            in1 => \N__32017\,
            in2 => \N__29560\,
            in3 => \N__52458\,
            lcout => n18026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15348_2_lut_LC_9_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42383\,
            in2 => \_gnd_net_\,
            in3 => \N__51996\,
            lcout => \c0.n17547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i16_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32396\,
            in2 => \_gnd_net_\,
            in3 => \N__34650\,
            lcout => \c0.FRAME_MATCHER_state_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50422\,
            ce => 'H',
            sr => \N__29551\
        );

    \c0.FRAME_MATCHER_state_i17_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30057\,
            in2 => \_gnd_net_\,
            in3 => \N__34649\,
            lcout => \c0.FRAME_MATCHER_state_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50430\,
            ce => 'H',
            sr => \N__30034\
        );

    \c0.i3_4_lut_adj_495_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32192\,
            in1 => \N__30055\,
            in2 => \N__29476\,
            in3 => \N__29503\,
            lcout => \c0.n16761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i28_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34641\,
            lcout => \c0.FRAME_MATCHER_state_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50437\,
            ce => 'H',
            sr => \N__29485\
        );

    \c0.i1_2_lut_adj_758_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29983\,
            in3 => \N__29504\,
            lcout => \c0.n16353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32193\,
            in2 => \_gnd_net_\,
            in3 => \N__29972\,
            lcout => \c0.n16377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_749_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__29472\,
            in1 => \_gnd_net_\,
            in2 => \N__29982\,
            in3 => \_gnd_net_\,
            lcout => \c0.n16361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_734_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30056\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29974\,
            lcout => \c0.n16345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_705_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30026\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29973\,
            lcout => \c0.n16339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i12_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32610\,
            in2 => \_gnd_net_\,
            in3 => \N__34647\,
            lcout => \c0.FRAME_MATCHER_state_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50443\,
            ce => 'H',
            sr => \N__32542\
        );

    \c0.data_out_frame2_0___i147_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36442\,
            in1 => \N__32529\,
            in2 => \_gnd_net_\,
            in3 => \N__51250\,
            lcout => data_out_frame2_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50455\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_640_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30133\,
            in1 => \N__29823\,
            in2 => \N__29788\,
            in3 => \N__29776\,
            lcout => \c0.n13464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48194\,
            in1 => \N__33556\,
            in2 => \_gnd_net_\,
            in3 => \N__34913\,
            lcout => \c0.n5_adj_2322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14911_3_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__37109\,
            in1 => \N__37434\,
            in2 => \_gnd_net_\,
            in3 => \N__35037\,
            lcout => OPEN,
            ltout => \c0.n17349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i2_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__37435\,
            in1 => \N__37538\,
            in2 => \N__29752\,
            in3 => \N__34978\,
            lcout => \c0.data_out_frame2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50455\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_238_Select_0_i3_2_lut_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29743\,
            in2 => \_gnd_net_\,
            in3 => \N__29581\,
            lcout => \c0.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__48209\,
            in1 => \N__30148\,
            in2 => \N__35071\,
            in3 => \N__48541\,
            lcout => \c0.n6_adj_2187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38607\,
            in1 => \N__48208\,
            in2 => \_gnd_net_\,
            in3 => \N__41521\,
            lcout => OPEN,
            ltout => \c0.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__48210\,
            in1 => \N__48542\,
            in2 => \N__30139\,
            in3 => \N__39021\,
            lcout => \c0.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14890_3_lut_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__37431\,
            in1 => \N__49525\,
            in2 => \_gnd_net_\,
            in3 => \N__35036\,
            lcout => OPEN,
            ltout => \c0.n17328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i8_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__37539\,
            in1 => \N__37432\,
            in2 => \N__30136\,
            in3 => \N__34977\,
            lcout => \c0.data_out_frame2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_596_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34912\,
            in2 => \_gnd_net_\,
            in3 => \N__38524\,
            lcout => \c0.n9758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__30129\,
            in1 => \N__34276\,
            in2 => \_gnd_net_\,
            in3 => \N__32397\,
            lcout => \c0.n16905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_adj_699_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__41703\,
            in1 => \_gnd_net_\,
            in2 => \N__33568\,
            in3 => \N__36073\,
            lcout => \c0.n16_adj_2197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i124_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36074\,
            in1 => \N__48839\,
            in2 => \_gnd_net_\,
            in3 => \N__51273\,
            lcout => data_out_frame2_15_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14899_3_lut_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__35809\,
            in1 => \N__37433\,
            in2 => \_gnd_net_\,
            in3 => \N__35035\,
            lcout => OPEN,
            ltout => \c0.n17337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i5_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37541\,
            in2 => \N__30349\,
            in3 => \N__31294\,
            lcout => \c0.data_out_frame2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i91_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36622\,
            in1 => \N__40861\,
            in2 => \_gnd_net_\,
            in3 => \N__51274\,
            lcout => data_out_frame2_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i4_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__32494\,
            in1 => \N__37540\,
            in2 => \_gnd_net_\,
            in3 => \N__31293\,
            lcout => \c0.data_out_frame2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1032_2_lut_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30346\,
            in2 => \_gnd_net_\,
            in3 => \N__30315\,
            lcout => \c0.n2338\,
            ltout => \c0.n2338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_661_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__30244\,
            in1 => \N__30223\,
            in2 => \N__30199\,
            in3 => \N__30196\,
            lcout => OPEN,
            ltout => \c0.n17_adj_2346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_662_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30172\,
            in1 => \N__30538\,
            in2 => \N__30160\,
            in3 => \N__30157\,
            lcout => n31,
            ltout => \n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_653_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__33356\,
            in1 => \N__33322\,
            in2 => \N__30151\,
            in3 => \N__34282\,
            lcout => \c0.n5_adj_2339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i127_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51279\,
            in1 => \N__49102\,
            in2 => \_gnd_net_\,
            in3 => \N__44378\,
            lcout => data_out_frame2_15_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i84_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36731\,
            in1 => \N__41815\,
            in2 => \_gnd_net_\,
            in3 => \N__51280\,
            lcout => data_out_frame2_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15387_3_lut_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__48227\,
            in1 => \N__38707\,
            in2 => \_gnd_net_\,
            in3 => \N__48667\,
            lcout => \c0.n17571\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_47_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__31039\,
            in1 => \N__30597\,
            in2 => \_gnd_net_\,
            in3 => \N__30910\,
            lcout => \c0.tx2.tx2_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14896_3_lut_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010001110100"
        )
    port map (
            in0 => \N__35017\,
            in1 => \N__37476\,
            in2 => \N__38717\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n17334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i6_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__37477\,
            in1 => \N__37553\,
            in2 => \N__30583\,
            in3 => \N__34957\,
            lcout => \c0.data_out_frame2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__43963\,
            in1 => \N__48665\,
            in2 => \N__41287\,
            in3 => \N__48226\,
            lcout => \c0.n6_adj_2278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_658_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001111011"
        )
    port map (
            in0 => \N__30579\,
            in1 => \N__30619\,
            in2 => \N__31759\,
            in3 => \N__30555\,
            lcout => \c0.n18_adj_2343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i4_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30524\,
            in1 => \N__30371\,
            in2 => \_gnd_net_\,
            in3 => \N__30442\,
            lcout => data_in_frame_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i77_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39210\,
            in1 => \N__35215\,
            in2 => \_gnd_net_\,
            in3 => \N__51180\,
            lcout => data_out_frame2_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17915_bdd_4_lut_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__41594\,
            in1 => \N__48666\,
            in2 => \N__49603\,
            in3 => \N__33655\,
            lcout => OPEN,
            ltout => \c0.n17918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15636_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__41662\,
            in1 => \N__51644\,
            in2 => \N__31303\,
            in3 => \N__47711\,
            lcout => \c0.n18107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i3_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__37554\,
            in1 => \N__31300\,
            in2 => \_gnd_net_\,
            in3 => \N__31284\,
            lcout => \c0.data_out_frame2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31273\,
            in1 => \N__31261\,
            in2 => \N__31249\,
            in3 => \N__31240\,
            lcout => \c0.n16148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i86_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__31936\,
            in1 => \N__31053\,
            in2 => \N__31230\,
            in3 => \N__31136\,
            lcout => \c0.data_in_frame_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__31552\,
            in1 => \N__31038\,
            in2 => \N__30943\,
            in3 => \N__30925\,
            lcout => \c0.tx2.n10101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15533_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__30901\,
            in1 => \N__48641\,
            in2 => \N__35986\,
            in3 => \N__48186\,
            lcout => \c0.n17981\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100010000"
        )
    port map (
            in0 => \N__30883\,
            in1 => \N__30802\,
            in2 => \N__30787\,
            in3 => \N__33661\,
            lcout => \r_SM_Main_0_adj_2441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i18_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__31934\,
            in1 => \N__30618\,
            in2 => \N__30694\,
            in3 => \N__32007\,
            lcout => \c0.data_in_frame_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i21_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32008\,
            in1 => \N__31935\,
            in2 => \N__31834\,
            in3 => \N__31758\,
            lcout => \c0.data_in_frame_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34020\,
            in1 => \N__34035\,
            in2 => \_gnd_net_\,
            in3 => \N__51993\,
            lcout => \c0.n2_adj_2298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14792_2_lut_3_lut_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__45920\,
            in1 => \N__31741\,
            in2 => \_gnd_net_\,
            in3 => \N__31671\,
            lcout => n17230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__7__2229_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011011100"
        )
    port map (
            in0 => \N__45544\,
            in1 => \N__31573\,
            in2 => \N__45982\,
            in3 => \N__46449\,
            lcout => data_out_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15355_2_lut_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__51994\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31572\,
            lcout => \c0.n17585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__33904\,
            in1 => \N__52257\,
            in2 => \N__39787\,
            in3 => \N__51995\,
            lcout => \c0.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i0_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31551\,
            in1 => \N__31420\,
            in2 => \_gnd_net_\,
            in3 => \N__31403\,
            lcout => \r_Clock_Count_0_adj_2454\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14960_3_lut_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32169\,
            in1 => \N__31377\,
            in2 => \_gnd_net_\,
            in3 => \N__32067\,
            lcout => n17398,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__0__2180_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__46855\,
            in1 => \N__46567\,
            in2 => \_gnd_net_\,
            in3 => \N__36271\,
            lcout => data_out_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i52_4_lut_LC_10_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__32038\,
            in1 => \N__43149\,
            in2 => \N__34114\,
            in3 => \N__52457\,
            lcout => OPEN,
            ltout => \c0.n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__35605\,
            in1 => \N__32082\,
            in2 => \N__32086\,
            in3 => \N__35520\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__35519\,
            in1 => \N__32068\,
            in2 => \N__35616\,
            in3 => \N__34093\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15210_3_lut_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__42701\,
            in1 => \N__40478\,
            in2 => \_gnd_net_\,
            in3 => \N__42467\,
            lcout => \c0.n17518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33987\,
            in1 => \N__32059\,
            in2 => \_gnd_net_\,
            in3 => \N__52062\,
            lcout => \c0.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10915_2_lut_LC_10_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39915\,
            in2 => \_gnd_net_\,
            in3 => \N__52042\,
            lcout => OPEN,
            ltout => \c0.n9_adj_2143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i50_4_lut_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__43147\,
            in1 => \N__32107\,
            in2 => \N__32041\,
            in3 => \N__52296\,
            lcout => \c0.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36820\,
            in1 => \N__39817\,
            in2 => \_gnd_net_\,
            in3 => \N__52040\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15562_LC_10_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__32032\,
            in1 => \N__52415\,
            in2 => \N__32020\,
            in3 => \N__52294\,
            lcout => \c0.n18023\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_10_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__32170\,
            in1 => \N__32128\,
            in2 => \N__35524\,
            in3 => \N__35615\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__52295\,
            in1 => \N__40000\,
            in2 => \N__38128\,
            in3 => \N__52041\,
            lcout => n10_adj_2423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15344_2_lut_LC_10_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__52039\,
            in1 => \N__35290\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n17592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__1__2243_LC_10_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111010"
        )
    port map (
            in0 => \N__32121\,
            in1 => \N__46421\,
            in2 => \N__45951\,
            in3 => \N__45536\,
            lcout => data_out_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18011_bdd_4_lut_LC_10_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__35260\,
            in1 => \N__34153\,
            in2 => \N__38146\,
            in3 => \N__52455\,
            lcout => \c0.n18014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18041_bdd_4_lut_LC_10_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__52454\,
            in1 => \N__32485\,
            in2 => \N__32152\,
            in3 => \N__34168\,
            lcout => OPEN,
            ltout => \n18044_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_773_LC_10_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__32137\,
            in1 => \N__43119\,
            in2 => \N__32131\,
            in3 => \N__52456\,
            lcout => n10_adj_2414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15336_3_lut_4_lut_LC_10_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42603\,
            in1 => \N__40341\,
            in2 => \N__40195\,
            in3 => \N__40242\,
            lcout => \c0.n17445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18077_bdd_4_lut_LC_10_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__43146\,
            in1 => \N__35419\,
            in2 => \N__32122\,
            in3 => \N__40366\,
            lcout => \c0.n18080\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_10_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32097\,
            in1 => \N__38380\,
            in2 => \_gnd_net_\,
            in3 => \N__52060\,
            lcout => \c0.n2_adj_2137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__4__2232_LC_10_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000100"
        )
    port map (
            in0 => \N__46437\,
            in1 => \N__46139\,
            in2 => \N__42660\,
            in3 => \N__32479\,
            lcout => \c0.data_out_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i0_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111111001111"
        )
    port map (
            in0 => \N__34248\,
            in1 => \N__32467\,
            in2 => \N__32458\,
            in3 => \N__32419\,
            lcout => \FRAME_MATCHER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_418_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__32190\,
            in1 => \N__34246\,
            in2 => \_gnd_net_\,
            in3 => \N__32389\,
            lcout => \c0.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_405_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__32191\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32325\,
            lcout => \c0.n6_adj_2140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_654_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32326\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33425\,
            lcout => OPEN,
            ltout => \c0.n16814_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_663_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__33533\,
            in1 => \N__32218\,
            in2 => \N__32206\,
            in3 => \N__34247\,
            lcout => \c0.n10052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_3_lut_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__51701\,
            in1 => \N__51535\,
            in2 => \_gnd_net_\,
            in3 => \N__47578\,
            lcout => \c0.tx2.n89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i31_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32194\,
            in2 => \_gnd_net_\,
            in3 => \N__34662\,
            lcout => \c0.FRAME_MATCHER_state_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50438\,
            ce => 'H',
            sr => \N__33292\
        );

    \c0.FRAME_MATCHER_i_i0_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33208\,
            in1 => \N__32959\,
            in2 => \_gnd_net_\,
            in3 => \N__32725\,
            lcout => \c0.FRAME_MATCHER_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50444\,
            ce => 'H',
            sr => \N__32626\
        );

    \c0.i15337_2_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35089\,
            in2 => \_gnd_net_\,
            in3 => \N__52080\,
            lcout => \c0.n17589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_717_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32588\,
            lcout => \c0.n16455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_723_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32609\,
            in2 => \_gnd_net_\,
            in3 => \N__32589\,
            lcout => \c0.n16449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15485_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__48456\,
            in1 => \N__38848\,
            in2 => \N__32530\,
            in3 => \N__48207\,
            lcout => \c0.n17927\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15641_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__34849\,
            in1 => \N__51631\,
            in2 => \N__34369\,
            in3 => \N__47642\,
            lcout => OPEN,
            ltout => \c0.n18119_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18119_bdd_4_lut_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__51632\,
            in1 => \N__35830\,
            in2 => \N__32515\,
            in3 => \N__34855\,
            lcout => OPEN,
            ltout => \c0.n18122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i2_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__34375\,
            in1 => \N__51763\,
            in2 => \N__32512\,
            in3 => \N__51633\,
            lcout => \c0.tx2.r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50456\,
            ce => \N__51451\,
            sr => \_gnd_net_\
        );

    \c0.i14902_3_lut_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__40147\,
            in1 => \N__37430\,
            in2 => \_gnd_net_\,
            in3 => \N__35034\,
            lcout => \c0.n17340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11148_2_lut_3_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111110"
        )
    port map (
            in0 => \N__33358\,
            in1 => \N__33321\,
            in2 => \N__33433\,
            in3 => \_gnd_net_\,
            lcout => \c0.n13496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_685_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35810\,
            in1 => \N__35869\,
            in2 => \N__37116\,
            in3 => \N__40146\,
            lcout => \c0.n9919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i60_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51147\,
            in2 => \N__33564\,
            in3 => \N__48844\,
            lcout => data_out_frame2_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_535_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33557\,
            in2 => \_gnd_net_\,
            in3 => \N__36076\,
            lcout => \c0.n9916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i52_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36736\,
            in1 => \N__34915\,
            in2 => \_gnd_net_\,
            in3 => \N__51277\,
            lcout => data_out_frame2_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15309_3_lut_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__48489\,
            in1 => \N__48065\,
            in2 => \_gnd_net_\,
            in3 => \N__37105\,
            lcout => \c0.n17579\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i98_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36249\,
            in1 => \N__41570\,
            in2 => \_gnd_net_\,
            in3 => \N__51278\,
            lcout => data_out_frame2_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_652_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33532\,
            in2 => \_gnd_net_\,
            in3 => \N__33429\,
            lcout => OPEN,
            ltout => \c0.n2_adj_2330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_636_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33357\,
            in1 => \N__33319\,
            in2 => \N__33295\,
            in3 => \N__34280\,
            lcout => \c0.n5545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_527_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35873\,
            in2 => \_gnd_net_\,
            in3 => \N__40152\,
            lcout => \c0.n16946\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_641_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41569\,
            in2 => \_gnd_net_\,
            in3 => \N__47371\,
            lcout => \c0.n16963\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_488_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49011\,
            in1 => \N__49743\,
            in2 => \N__43728\,
            in3 => \N__33586\,
            lcout => \c0.n17073\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_564_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45362\,
            lcout => \c0.n9754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15505_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__47231\,
            in1 => \N__48043\,
            in2 => \N__48564\,
            in3 => \N__36069\,
            lcout => \c0.n17951\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i130_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36245\,
            in1 => \N__39127\,
            in2 => \_gnd_net_\,
            in3 => \N__51276\,
            lcout => data_out_frame2_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i112_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51275\,
            in1 => \N__44012\,
            in2 => \_gnd_net_\,
            in3 => \N__43724\,
            lcout => data_out_frame2_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_694_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35237\,
            in1 => \N__44345\,
            in2 => \_gnd_net_\,
            in3 => \N__41345\,
            lcout => \c0.n17091\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15465_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__48044\,
            in1 => \N__38779\,
            in2 => \N__49744\,
            in3 => \N__48465\,
            lcout => \c0.n17891\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_637_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35238\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44346\,
            lcout => \c0.n16936\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i145_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__34806\,
            in1 => \_gnd_net_\,
            in2 => \N__39547\,
            in3 => \N__51213\,
            lcout => data_out_frame2_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17987_bdd_4_lut_4_lut_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011000"
        )
    port map (
            in0 => \N__39301\,
            in1 => \N__48224\,
            in2 => \N__35814\,
            in3 => \N__47712\,
            lcout => \c0.n17990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15475_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__48578\,
            in1 => \N__48223\,
            in2 => \N__49469\,
            in3 => \N__47181\,
            lcout => \c0.n17915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i97_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39545\,
            in1 => \N__47360\,
            in2 => \_gnd_net_\,
            in3 => \N__51214\,
            lcout => data_out_frame2_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i146_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51212\,
            in2 => \N__33643\,
            in3 => \N__36250\,
            lcout => data_out_frame2_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15470_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__48225\,
            in1 => \N__33639\,
            in2 => \N__49216\,
            in3 => \N__48579\,
            lcout => OPEN,
            ltout => \c0.n17909_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17909_bdd_4_lut_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__39126\,
            in1 => \N__37867\,
            in2 => \N__33631\,
            in3 => \N__48493\,
            lcout => \c0.n17912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18107_bdd_4_lut_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__33628\,
            in1 => \N__33619\,
            in2 => \N__33613\,
            in3 => \N__51645\,
            lcout => \c0.n18110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__47815\,
            in1 => \N__33601\,
            in2 => \N__35908\,
            in3 => \N__47713\,
            lcout => OPEN,
            ltout => \c0.n22_adj_2359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i1_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__51646\,
            in1 => \N__33595\,
            in2 => \N__33589\,
            in3 => \N__51762\,
            lcout => \c0.tx2.r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50512\,
            ce => \N__51404\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15567_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__52451\,
            in1 => \N__33937\,
            in2 => \N__33895\,
            in3 => \N__52290\,
            lcout => OPEN,
            ltout => \c0.n18029_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18029_bdd_4_lut_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__33925\,
            in1 => \N__33916\,
            in2 => \N__33907\,
            in3 => \N__52452\,
            lcout => n18032,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40508\,
            in1 => \N__46856\,
            in2 => \_gnd_net_\,
            in3 => \N__52064\,
            lcout => \c0.n8_adj_2138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_15528_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010110000"
        )
    port map (
            in0 => \N__35143\,
            in1 => \N__47660\,
            in2 => \N__48629\,
            in3 => \N__36028\,
            lcout => \c0.n17897\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34141\,
            in1 => \N__46201\,
            in2 => \_gnd_net_\,
            in3 => \N__52063\,
            lcout => \c0.n5_adj_2299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__0__2172_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39760\,
            in1 => \N__40087\,
            in2 => \_gnd_net_\,
            in3 => \N__37993\,
            lcout => \c0.data_out_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50530\,
            ce => \N__46589\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__4__2160_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38034\,
            in1 => \N__33958\,
            in2 => \_gnd_net_\,
            in3 => \N__35305\,
            lcout => \c0.data_out_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50530\,
            ce => \N__46589\,
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__33834\,
            in1 => \N__33790\,
            in2 => \_gnd_net_\,
            in3 => \N__33731\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__2__2226_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__46485\,
            in1 => \N__35272\,
            in2 => \N__45990\,
            in3 => \N__45547\,
            lcout => data_out_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__5__2215_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__45545\,
            in1 => \N__34036\,
            in2 => \N__45976\,
            in3 => \N__46487\,
            lcout => data_out_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__5__2223_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111110000"
        )
    port map (
            in0 => \N__46486\,
            in1 => \N__45546\,
            in2 => \N__34024\,
            in3 => \N__45911\,
            lcout => data_out_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_501_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46654\,
            in1 => \N__40504\,
            in2 => \N__34009\,
            in3 => \N__36827\,
            lcout => \c0.n10_adj_2276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_664_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34196\,
            in1 => \N__46853\,
            in2 => \N__39706\,
            in3 => \N__40408\,
            lcout => \c0.n16990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__5__2183_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__36514\,
            in1 => \N__34355\,
            in2 => \N__34140\,
            in3 => \N__42798\,
            lcout => \c0.data_out_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__6__2230_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__46447\,
            in1 => \N__45943\,
            in2 => \N__33991\,
            in3 => \N__45487\,
            lcout => data_out_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__0__2228_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011011100"
        )
    port map (
            in0 => \N__45486\,
            in1 => \N__33972\,
            in2 => \N__45989\,
            in3 => \N__46448\,
            lcout => data_out_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_550_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46854\,
            in1 => \N__34198\,
            in2 => \_gnd_net_\,
            in3 => \N__40414\,
            lcout => \c0.n9509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__2__2170_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__38097\,
            in1 => \N__37972\,
            in2 => \N__42761\,
            in3 => \N__42822\,
            lcout => data_out_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_544_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38025\,
            in1 => \N__34197\,
            in2 => \_gnd_net_\,
            in3 => \N__34133\,
            lcout => \c0.n9505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i53_4_lut_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__45191\,
            in1 => \N__52289\,
            in2 => \N__34087\,
            in3 => \N__52061\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__4__2184_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__42864\,
            in1 => \N__34348\,
            in2 => \N__36828\,
            in3 => \N__36535\,
            lcout => \c0.data_out_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_769_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__34102\,
            in1 => \N__43148\,
            in2 => \N__39970\,
            in3 => \N__52405\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__40550\,
            in1 => \N__39705\,
            in2 => \N__52097\,
            in3 => \_gnd_net_\,
            lcout => \c0.n5_adj_2142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__0__2220_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__45492\,
            in1 => \N__42131\,
            in2 => \N__45988\,
            in3 => \N__34074\,
            lcout => data_out_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15297_2_lut_LC_11_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__52076\,
            in1 => \N__34060\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n17588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15417_2_lut_3_lut_4_lut_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__45491\,
            in1 => \N__42680\,
            in2 => \N__45987\,
            in3 => \N__46466\,
            lcout => \c0.n10054\,
            ltout => \c0.n10054_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__6__2182_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__42865\,
            in1 => \N__36493\,
            in2 => \N__34039\,
            in3 => \N__38029\,
            lcout => \c0.data_out_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52054\,
            in2 => \N__47049\,
            in3 => \N__46689\,
            lcout => \c0.n5_adj_2208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__7__2181_LC_11_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__36472\,
            in1 => \N__34195\,
            in2 => \N__34356\,
            in3 => \N__42863\,
            lcout => \c0.data_out_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34194\,
            in1 => \N__52056\,
            in2 => \_gnd_net_\,
            in3 => \N__40270\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15616_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__35668\,
            in1 => \N__52465\,
            in2 => \N__34171\,
            in3 => \N__52231\,
            lcout => \c0.n18041\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_522_LC_11_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__47045\,
            in1 => \N__42937\,
            in2 => \_gnd_net_\,
            in3 => \N__40241\,
            lcout => \c0.n16981\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15370_2_lut_LC_11_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52055\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40474\,
            lcout => OPEN,
            ltout => \c0.n17543_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15552_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__52230\,
            in1 => \N__34162\,
            in2 => \N__34156\,
            in3 => \N__52453\,
            lcout => \c0.n18011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__1__2187_LC_11_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__46434\,
            in1 => \N__45956\,
            in2 => \N__36319\,
            in3 => \N__34147\,
            lcout => \c0.data_out_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50577\,
            ce => \N__34357\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__2__2186_LC_11_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__42725\,
            in1 => \N__40335\,
            in2 => \N__45640\,
            in3 => \N__46435\,
            lcout => \c0.data_out_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50577\,
            ce => \N__34357\,
            sr => \_gnd_net_\
        );

    \c0.i15208_2_lut_LC_11_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36562\,
            in2 => \_gnd_net_\,
            in3 => \N__45954\,
            lcout => OPEN,
            ltout => \c0.n17456_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__3__2185_LC_11_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__42726\,
            in1 => \N__45069\,
            in2 => \N__34360\,
            in3 => \N__46436\,
            lcout => \c0.data_out_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50577\,
            ce => \N__34357\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__0__2188_LC_11_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__46433\,
            in1 => \N__45955\,
            in2 => \N__36346\,
            in3 => \N__40162\,
            lcout => \c0.data_out_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50577\,
            ce => \N__34357\,
            sr => \_gnd_net_\
        );

    \i14716_2_lut_3_lut_LC_11_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__45953\,
            in1 => \N__46432\,
            in2 => \_gnd_net_\,
            in3 => \N__34321\,
            lcout => n17154,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i139_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36620\,
            in1 => \N__34392\,
            in2 => \_gnd_net_\,
            in3 => \N__51223\,
            lcout => data_out_frame2_17_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7942_2_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34683\,
            in2 => \_gnd_net_\,
            in3 => \N__34262\,
            lcout => \c0.n10297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2353__i0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34219\,
            in2 => \N__48096\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter2_0\,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \c0.n15615\,
            clk => \N__50446\,
            ce => \N__34690\,
            sr => \N__34672\
        );

    \c0.byte_transmit_counter2_2353__i1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48354\,
            in2 => \_gnd_net_\,
            in3 => \N__34207\,
            lcout => \c0.byte_transmit_counter2_1\,
            ltout => OPEN,
            carryin => \c0.n15615\,
            carryout => \c0.n15616\,
            clk => \N__50446\,
            ce => \N__34690\,
            sr => \N__34672\
        );

    \c0.byte_transmit_counter2_2353__i2_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47658\,
            in2 => \_gnd_net_\,
            in3 => \N__34204\,
            lcout => \c0.byte_transmit_counter2_2\,
            ltout => OPEN,
            carryin => \c0.n15616\,
            carryout => \c0.n15617\,
            clk => \N__50446\,
            ce => \N__34690\,
            sr => \N__34672\
        );

    \c0.byte_transmit_counter2_2353__i3_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51576\,
            in2 => \_gnd_net_\,
            in3 => \N__34201\,
            lcout => \c0.byte_transmit_counter2_3\,
            ltout => OPEN,
            carryin => \c0.n15617\,
            carryout => \c0.n15618\,
            clk => \N__50446\,
            ce => \N__34690\,
            sr => \N__34672\
        );

    \c0.byte_transmit_counter2_2353__i4_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51714\,
            in2 => \_gnd_net_\,
            in3 => \N__34759\,
            lcout => \c0.byte_transmit_counter2_4\,
            ltout => OPEN,
            carryin => \c0.n15618\,
            carryout => \c0.n15619\,
            clk => \N__50446\,
            ce => \N__34690\,
            sr => \N__34672\
        );

    \c0.byte_transmit_counter2_2353__i5_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34752\,
            in2 => \_gnd_net_\,
            in3 => \N__34738\,
            lcout => \c0.byte_transmit_counter2_5\,
            ltout => OPEN,
            carryin => \c0.n15619\,
            carryout => \c0.n15620\,
            clk => \N__50446\,
            ce => \N__34690\,
            sr => \N__34672\
        );

    \c0.byte_transmit_counter2_2353__i6_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34728\,
            in2 => \_gnd_net_\,
            in3 => \N__34714\,
            lcout => \c0.byte_transmit_counter2_6\,
            ltout => OPEN,
            carryin => \c0.n15620\,
            carryout => \c0.n15621\,
            clk => \N__50446\,
            ce => \N__34690\,
            sr => \N__34672\
        );

    \c0.byte_transmit_counter2_2353__i7_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34704\,
            in2 => \_gnd_net_\,
            in3 => \N__34711\,
            lcout => \c0.byte_transmit_counter2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50446\,
            ce => \N__34690\,
            sr => \N__34672\
        );

    \c0.FRAME_MATCHER_state_i9_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34431\,
            in2 => \_gnd_net_\,
            in3 => \N__34651\,
            lcout => \c0.FRAME_MATCHER_state_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50457\,
            ce => 'H',
            sr => \N__34411\
        );

    \c0.n17927_bdd_4_lut_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__48459\,
            in1 => \N__34405\,
            in2 => \N__34399\,
            in3 => \N__37043\,
            lcout => OPEN,
            ltout => \c0.n17930_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__47817\,
            in1 => \N__36919\,
            in2 => \N__34378\,
            in3 => \N__47645\,
            lcout => \c0.n22_adj_2358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17933_bdd_4_lut_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__48458\,
            in1 => \N__43380\,
            in2 => \N__49283\,
            in3 => \N__35971\,
            lcout => \c0.n17936\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_551_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44646\,
            in1 => \N__36987\,
            in2 => \N__41968\,
            in3 => \N__39049\,
            lcout => \c0.n28_adj_2294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__35959\,
            in1 => \N__48460\,
            in2 => \N__37672\,
            in3 => \N__48066\,
            lcout => \c0.n6_adj_2201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17939_bdd_4_lut_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__48457\,
            in1 => \N__34924\,
            in2 => \N__43908\,
            in3 => \N__38514\,
            lcout => \c0.n17942\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14863_4_lut_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__48492\,
            in1 => \N__35779\,
            in2 => \N__34843\,
            in3 => \N__47643\,
            lcout => OPEN,
            ltout => \c0.n17301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14865_3_lut_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39229\,
            in2 => \N__34828\,
            in3 => \N__51617\,
            lcout => OPEN,
            ltout => \c0.n17303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i0_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__51618\,
            in1 => \N__34765\,
            in2 => \N__34825\,
            in3 => \N__51739\,
            lcout => \c0.tx2.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50479\,
            ce => \N__51452\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__34807\,
            in1 => \N__48490\,
            in2 => \N__36943\,
            in3 => \N__48052\,
            lcout => OPEN,
            ltout => \c0.n18101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18101_bdd_4_lut_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48491\,
            in1 => \N__34792\,
            in2 => \N__34771\,
            in3 => \N__43847\,
            lcout => OPEN,
            ltout => \c0.n18104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__47644\,
            in1 => \N__35884\,
            in2 => \N__34768\,
            in3 => \N__47816\,
            lcout => \c0.n22_adj_2337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_642_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43690\,
            lcout => \c0.n17106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15495_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__48051\,
            in1 => \N__40871\,
            in2 => \N__48580\,
            in3 => \N__35166\,
            lcout => \c0.n17939\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_4_lut_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41344\,
            in1 => \N__40979\,
            in2 => \N__36756\,
            in3 => \N__39598\,
            lcout => \c0.n18_adj_2251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_595_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38522\,
            in1 => \N__34914\,
            in2 => \_gnd_net_\,
            in3 => \N__38580\,
            lcout => \c0.n17118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_626_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43771\,
            in1 => \N__45367\,
            in2 => \N__37738\,
            in3 => \N__35062\,
            lcout => \c0.n17061\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_453_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37304\,
            in1 => \N__41017\,
            in2 => \N__34891\,
            in3 => \N__34876\,
            lcout => \c0.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_451_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41343\,
            in1 => \N__47224\,
            in2 => \N__44806\,
            in3 => \N__38752\,
            lcout => \c0.n22_adj_2194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_532_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__37303\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44282\,
            lcout => \c0.n9901\,
            ltout => \c0.n9901_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_473_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34867\,
            in1 => \N__35874\,
            in2 => \N__34858\,
            in3 => \N__41704\,
            lcout => \c0.n19_adj_2254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i122_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51196\,
            in1 => \N__37911\,
            in2 => \_gnd_net_\,
            in3 => \N__47188\,
            lcout => data_out_frame2_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i44_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37953\,
            in1 => \N__35064\,
            in2 => \_gnd_net_\,
            in3 => \N__51198\,
            lcout => data_out_frame2_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_526_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47313\,
            in1 => \N__41238\,
            in2 => \N__38724\,
            in3 => \N__37606\,
            lcout => \c0.n9692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_605_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35159\,
            in2 => \_gnd_net_\,
            in3 => \N__43573\,
            lcout => \c0.n9707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i58_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51197\,
            in1 => \N__37912\,
            in2 => \_gnd_net_\,
            in3 => \N__38600\,
            lcout => data_out_frame2_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14893_3_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__48694\,
            in1 => \N__37454\,
            in2 => \_gnd_net_\,
            in3 => \N__35038\,
            lcout => OPEN,
            ltout => \c0.n17331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i7_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__37455\,
            in1 => \N__37552\,
            in2 => \N__34981\,
            in3 => \N__34976\,
            lcout => \c0.data_out_frame2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17891_bdd_4_lut_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__34930\,
            in1 => \N__37731\,
            in2 => \N__45256\,
            in3 => \N__48391\,
            lcout => \c0.n17894\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i129_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51073\,
            in2 => \N__39533\,
            in3 => \N__43831\,
            lcout => data_out_frame2_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i125_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37767\,
            in1 => \N__44160\,
            in2 => \_gnd_net_\,
            in3 => \N__51211\,
            lcout => data_out_frame2_15_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i83_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51210\,
            in1 => \N__44487\,
            in2 => \_gnd_net_\,
            in3 => \N__35165\,
            lcout => data_out_frame2_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37580\,
            in1 => \N__47962\,
            in2 => \_gnd_net_\,
            in3 => \N__37756\,
            lcout => \c0.n12_adj_2305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11219217_i1_3_lut_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35134\,
            in1 => \N__35404\,
            in2 => \_gnd_net_\,
            in3 => \N__51613\,
            lcout => \c0.n15_adj_2356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15538_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__47963\,
            in1 => \N__48392\,
            in2 => \N__38570\,
            in3 => \N__41140\,
            lcout => OPEN,
            ltout => \c0.n17993_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17993_bdd_4_lut_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48393\,
            in1 => \N__41868\,
            in2 => \N__35128\,
            in3 => \N__44854\,
            lcout => OPEN,
            ltout => \c0.n17393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15606_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__35125\,
            in1 => \N__51614\,
            in2 => \N__35119\,
            in3 => \N__47631\,
            lcout => OPEN,
            ltout => \c0.n17963_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17963_bdd_4_lut_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__51615\,
            in1 => \N__35116\,
            in2 => \N__35107\,
            in3 => \N__44581\,
            lcout => OPEN,
            ltout => \c0.n17966_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i5_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__51761\,
            in1 => \N__51616\,
            in2 => \N__35104\,
            in3 => \N__36115\,
            lcout => \c0.tx2.r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50521\,
            ce => \N__51411\,
            sr => \_gnd_net_\
        );

    \c0.data_out_0__5__2239_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__42156\,
            in1 => \N__45978\,
            in2 => \N__45537\,
            in3 => \N__35085\,
            lcout => data_out_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i66_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36231\,
            in1 => \N__47270\,
            in2 => \_gnd_net_\,
            in3 => \N__51178\,
            lcout => data_out_frame2_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i86_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40619\,
            in1 => \N__38569\,
            in2 => \_gnd_net_\,
            in3 => \N__51179\,
            lcout => data_out_frame2_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37838\,
            in1 => \N__48107\,
            in2 => \_gnd_net_\,
            in3 => \N__42072\,
            lcout => \c0.n9_adj_2347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__3__2241_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011011100"
        )
    port map (
            in0 => \N__45510\,
            in1 => \N__35286\,
            in2 => \N__45999\,
            in3 => \N__46492\,
            lcout => data_out_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i149_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37348\,
            in1 => \N__37236\,
            in2 => \_gnd_net_\,
            in3 => \N__51177\,
            lcout => data_out_frame2_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35247\,
            in1 => \N__52065\,
            in2 => \_gnd_net_\,
            in3 => \N__35271\,
            lcout => \c0.n2_adj_2291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15249_3_lut_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__45206\,
            in1 => \N__42752\,
            in2 => \_gnd_net_\,
            in3 => \N__40480\,
            lcout => \c0.n17514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__2__2218_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__35248\,
            in1 => \N__45977\,
            in2 => \N__42155\,
            in3 => \N__45514\,
            lcout => data_out_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50542\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48121\,
            in1 => \N__35236\,
            in2 => \_gnd_net_\,
            in3 => \N__49343\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17897_bdd_4_lut_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__35185\,
            in1 => \N__35173\,
            in2 => \N__35407\,
            in3 => \N__47632\,
            lcout => \c0.n17900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4030_2_lut_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45936\,
            in2 => \_gnd_net_\,
            in3 => \N__46481\,
            lcout => n2547,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_667_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47139\,
            in1 => \N__52511\,
            in2 => \N__46702\,
            in3 => \N__39786\,
            lcout => \c0.n16975\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_15631_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__47530\,
            in1 => \N__45565\,
            in2 => \N__35392\,
            in3 => \N__35350\,
            lcout => \c0.tx2.n17903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_643_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43011\,
            in1 => \N__39877\,
            in2 => \_gnd_net_\,
            in3 => \N__40412\,
            lcout => \c0.n32_adj_2297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__3__2177_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__42753\,
            in1 => \N__36390\,
            in2 => \N__42861\,
            in3 => \N__43012\,
            lcout => \c0.data_out_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_683_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__42284\,
            in1 => \N__38101\,
            in2 => \_gnd_net_\,
            in3 => \N__42400\,
            lcout => \c0.n17055\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_539_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38102\,
            in1 => \N__46804\,
            in2 => \_gnd_net_\,
            in3 => \N__46898\,
            lcout => OPEN,
            ltout => \c0.n16978_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_507_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35304\,
            in1 => \N__35659\,
            in2 => \N__35293\,
            in3 => \N__46719\,
            lcout => \c0.n20_adj_2282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__4__2176_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__36372\,
            in1 => \N__42843\,
            in2 => \N__42762\,
            in3 => \N__42958\,
            lcout => data_out_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_689_LC_12_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35701\,
            in2 => \_gnd_net_\,
            in3 => \N__42957\,
            lcout => \c0.n9728\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_499_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45114\,
            in1 => \N__42469\,
            in2 => \N__40524\,
            in3 => \N__42936\,
            lcout => \c0.n16969\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_513_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40336\,
            in2 => \_gnd_net_\,
            in3 => \N__45070\,
            lcout => \c0.n16912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_3_lut_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__38096\,
            in1 => \N__39871\,
            in2 => \N__52098\,
            in3 => \_gnd_net_\,
            lcout => \c0.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18035_bdd_4_lut_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__35641\,
            in1 => \N__35677\,
            in2 => \N__35635\,
            in3 => \N__52406\,
            lcout => OPEN,
            ltout => \n18038_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_771_LC_12_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__52407\,
            in1 => \N__38191\,
            in2 => \N__35620\,
            in3 => \N__43153\,
            lcout => OPEN,
            ltout => \n10_adj_2413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__35602\,
            in1 => \N__35433\,
            in2 => \N__35527\,
            in3 => \N__35523\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__1__2203_LC_12_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46403\,
            in1 => \N__45785\,
            in2 => \N__42751\,
            in3 => \N__36645\,
            lcout => \c0.data_out_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50578\,
            ce => \N__46131\,
            sr => \_gnd_net_\
        );

    \c0.data_out_1__1__2235_LC_12_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__46402\,
            in1 => \N__45784\,
            in2 => \N__42750\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50578\,
            ce => \N__46131\,
            sr => \_gnd_net_\
        );

    \c0.mux_1210_i1_3_lut_LC_12_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45782\,
            in1 => \N__42712\,
            in2 => \_gnd_net_\,
            in3 => \N__46401\,
            lcout => n2652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_LC_12_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__45781\,
            in1 => \N__42711\,
            in2 => \_gnd_net_\,
            in3 => \N__46400\,
            lcout => \c0.n10181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__6__2190_LC_12_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__45783\,
            in1 => \N__36669\,
            in2 => \N__37789\,
            in3 => \N__46404\,
            lcout => \c0.data_out_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50578\,
            ce => \N__46131\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_12_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38033\,
            in1 => \N__35700\,
            in2 => \_gnd_net_\,
            in3 => \N__52071\,
            lcout => \c0.n5_adj_2300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15362_2_lut_LC_12_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52072\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40322\,
            lcout => OPEN,
            ltout => \c0.n17555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15572_LC_12_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__35686\,
            in1 => \N__52464\,
            in2 => \N__35680\,
            in3 => \N__52303\,
            lcout => \c0.n18035\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__6__2198_LC_12_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36870\,
            in2 => \_gnd_net_\,
            in3 => \N__45997\,
            lcout => \c0.data_out_7__2__N_447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50584\,
            ce => \N__46137\,
            sr => \N__41896\
        );

    \c0.data_out_5__7__2197_LC_12_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36849\,
            in2 => \_gnd_net_\,
            in3 => \N__45998\,
            lcout => \c0.data_out_7__3__N_441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50584\,
            ce => \N__46137\,
            sr => \N__41896\
        );

    \c0.i15281_2_lut_LC_12_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45057\,
            in2 => \_gnd_net_\,
            in3 => \N__52070\,
            lcout => \c0.n17569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_645_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36961\,
            in1 => \N__40875\,
            in2 => \N__35941\,
            in3 => \N__43584\,
            lcout => \c0.n20_adj_2333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15324_2_lut_3_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__35875\,
            in1 => \N__48353\,
            in2 => \_gnd_net_\,
            in3 => \N__48009\,
            lcout => \c0.n17578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_470_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40978\,
            in2 => \_gnd_net_\,
            in3 => \N__39597\,
            lcout => \c0.n17121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_572_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43651\,
            in2 => \_gnd_net_\,
            in3 => \N__40803\,
            lcout => \c0.n9810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_630_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43464\,
            in2 => \_gnd_net_\,
            in3 => \N__37148\,
            lcout => \c0.n9859\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i67_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36441\,
            in1 => \N__38518\,
            in2 => \_gnd_net_\,
            in3 => \N__51183\,
            lcout => data_out_frame2_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_450_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35818\,
            in1 => \N__37587\,
            in2 => \_gnd_net_\,
            in3 => \N__37771\,
            lcout => \c0.n17124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i131_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36439\,
            in1 => \N__37053\,
            in2 => \_gnd_net_\,
            in3 => \N__51136\,
            lcout => data_out_frame2_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i99_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51135\,
            in1 => \N__36440\,
            in2 => \_gnd_net_\,
            in3 => \N__49272\,
            lcout => data_out_frame2_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__47961\,
            in1 => \N__48513\,
            in2 => \N__37126\,
            in3 => \N__44737\,
            lcout => \c0.n6_adj_2335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40977\,
            in1 => \N__47960\,
            in2 => \_gnd_net_\,
            in3 => \N__44442\,
            lcout => \c0.n5_adj_2317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i49_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41755\,
            in1 => \N__37150\,
            in2 => \_gnd_net_\,
            in3 => \N__51137\,
            lcout => data_out_frame2_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_486_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49702\,
            in1 => \N__43902\,
            in2 => \N__38470\,
            in3 => \N__35950\,
            lcout => \c0.n15_adj_2269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i76_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37957\,
            in1 => \N__37302\,
            in2 => \_gnd_net_\,
            in3 => \N__51138\,
            lcout => data_out_frame2_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_624_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37847\,
            in1 => \N__49271\,
            in2 => \N__37668\,
            in3 => \N__43646\,
            lcout => \c0.n16957\,
            ltout => \c0.n16957_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_570_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35937\,
            in1 => \N__35892\,
            in2 => \N__35917\,
            in3 => \N__37693\,
            lcout => \c0.n21_adj_2304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i162_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35914\,
            in1 => \N__41938\,
            in2 => \N__36892\,
            in3 => \N__37060\,
            lcout => \c0.data_out_frame2_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50492\,
            ce => \N__51184\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i161_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__35893\,
            in1 => \N__38683\,
            in2 => \_gnd_net_\,
            in3 => \N__40828\,
            lcout => \c0.data_out_frame2_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50492\,
            ce => \N__51184\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_562_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37664\,
            in2 => \_gnd_net_\,
            in3 => \N__37848\,
            lcout => \c0.n9886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_448_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43477\,
            in1 => \N__49431\,
            in2 => \N__41067\,
            in3 => \N__36016\,
            lcout => OPEN,
            ltout => \c0.n16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i167_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36007\,
            in1 => \N__37081\,
            in2 => \N__35995\,
            in3 => \N__36967\,
            lcout => \c0.data_out_frame2_20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50503\,
            ce => \N__50965\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_696_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44284\,
            in1 => \N__37736\,
            in2 => \_gnd_net_\,
            in3 => \N__49007\,
            lcout => \c0.n17112\,
            ltout => \c0.n17112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_580_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38664\,
            in1 => \N__38455\,
            in2 => \N__35992\,
            in3 => \N__39403\,
            lcout => OPEN,
            ltout => \c0.n14_adj_2308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i158_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__38545\,
            in1 => \N__37165\,
            in2 => \N__35989\,
            in3 => \N__47415\,
            lcout => \c0.data_out_frame2_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50503\,
            ce => \N__50965\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_620_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37652\,
            in1 => \N__43647\,
            in2 => \_gnd_net_\,
            in3 => \N__40782\,
            lcout => \c0.n17067\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i63_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50939\,
            in1 => \N__49106\,
            in2 => \_gnd_net_\,
            in3 => \N__44354\,
            lcout => data_out_frame2_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15490_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__48584\,
            in1 => \N__48042\,
            in2 => \N__39159\,
            in3 => \N__39589\,
            lcout => \c0.n17933\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i116_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50937\,
            in1 => \_gnd_net_\,
            in2 => \N__36735\,
            in3 => \N__47237\,
            lcout => data_out_frame2_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i111_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48935\,
            in1 => \N__49651\,
            in2 => \_gnd_net_\,
            in3 => \N__50941\,
            lcout => data_out_frame2_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_518_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39334\,
            in1 => \N__37594\,
            in2 => \N__49658\,
            in3 => \N__37206\,
            lcout => \c0.n17133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_588_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40717\,
            in1 => \N__36075\,
            in2 => \N__44736\,
            in3 => \N__39014\,
            lcout => \c0.n9865\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i59_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50938\,
            in1 => \_gnd_net_\,
            in2 => \N__36621\,
            in3 => \N__40983\,
            lcout => data_out_frame2_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i109_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39203\,
            in1 => \N__36043\,
            in2 => \_gnd_net_\,
            in3 => \N__50940\,
            lcout => data_out_frame2_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_589_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39151\,
            in2 => \_gnd_net_\,
            in3 => \N__36042\,
            lcout => \c0.n9814\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36041\,
            in1 => \N__38439\,
            in2 => \_gnd_net_\,
            in3 => \N__48030\,
            lcout => \c0.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i101_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__38440\,
            in1 => \_gnd_net_\,
            in2 => \N__37353\,
            in3 => \N__50923\,
            lcout => data_out_frame2_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i133_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50921\,
            in1 => \N__37344\,
            in2 => \_gnd_net_\,
            in3 => \N__40781\,
            lcout => data_out_frame2_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i123_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36619\,
            in1 => \N__39152\,
            in2 => \_gnd_net_\,
            in3 => \N__50924\,
            lcout => data_out_frame2_15_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17981_bdd_4_lut_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__36130\,
            in1 => \N__48586\,
            in2 => \N__36108\,
            in3 => \N__41406\,
            lcout => OPEN,
            ltout => \c0.n17984_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__38905\,
            in1 => \N__47804\,
            in2 => \N__36118\,
            in3 => \N__47706\,
            lcout => \c0.n22_adj_2354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i142_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50922\,
            in1 => \_gnd_net_\,
            in2 => \N__36109\,
            in3 => \N__44557\,
            lcout => data_out_frame2_17_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i0_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39522\,
            in2 => \_gnd_net_\,
            in3 => \N__36094\,
            lcout => rand_data_0,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => n15528,
            clk => \N__50532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i1_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36224\,
            in2 => \_gnd_net_\,
            in3 => \N__36091\,
            lcout => rand_data_1,
            ltout => OPEN,
            carryin => n15528,
            carryout => n15529,
            clk => \N__50532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i2_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36418\,
            in2 => \_gnd_net_\,
            in3 => \N__36088\,
            lcout => rand_data_2,
            ltout => OPEN,
            carryin => n15529,
            carryout => n15530,
            clk => \N__50532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i3_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49780\,
            in2 => \_gnd_net_\,
            in3 => \N__36085\,
            lcout => rand_data_3,
            ltout => OPEN,
            carryin => n15530,
            carryout => n15531,
            clk => \N__50532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i4_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37343\,
            in2 => \_gnd_net_\,
            in3 => \N__36082\,
            lcout => rand_data_4,
            ltout => OPEN,
            carryin => n15531,
            carryout => n15532,
            clk => \N__50532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i5_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41444\,
            in2 => \_gnd_net_\,
            in3 => \N__36079\,
            lcout => rand_data_5,
            ltout => OPEN,
            carryin => n15532,
            carryout => n15533,
            clk => \N__50532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i6_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49878\,
            in2 => \_gnd_net_\,
            in3 => \N__36160\,
            lcout => rand_data_6,
            ltout => OPEN,
            carryin => n15533,
            carryout => n15534,
            clk => \N__50532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i7_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51304\,
            in2 => \_gnd_net_\,
            in3 => \N__36157\,
            lcout => rand_data_7,
            ltout => OPEN,
            carryin => n15534,
            carryout => n15535,
            clk => \N__50532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i8_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48732\,
            in2 => \_gnd_net_\,
            in3 => \N__36154\,
            lcout => rand_data_8,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => n15536,
            clk => \N__50543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i9_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37896\,
            in2 => \_gnd_net_\,
            in3 => \N__36151\,
            lcout => rand_data_9,
            ltout => OPEN,
            carryin => n15536,
            carryout => n15537,
            clk => \N__50543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i10_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36596\,
            in2 => \_gnd_net_\,
            in3 => \N__36148\,
            lcout => rand_data_10,
            ltout => OPEN,
            carryin => n15537,
            carryout => n15538,
            clk => \N__50543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i11_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48815\,
            in2 => \_gnd_net_\,
            in3 => \N__36145\,
            lcout => rand_data_11,
            ltout => OPEN,
            carryin => n15538,
            carryout => n15539,
            clk => \N__50543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i12_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44139\,
            in2 => \_gnd_net_\,
            in3 => \N__36142\,
            lcout => rand_data_12,
            ltout => OPEN,
            carryin => n15539,
            carryout => n15540,
            clk => \N__50543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i13_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44547\,
            in2 => \_gnd_net_\,
            in3 => \N__36139\,
            lcout => rand_data_13,
            ltout => OPEN,
            carryin => n15540,
            carryout => n15541,
            clk => \N__50543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i14_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49073\,
            in2 => \_gnd_net_\,
            in3 => \N__36136\,
            lcout => rand_data_14,
            ltout => OPEN,
            carryin => n15541,
            carryout => n15542,
            clk => \N__50543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i15_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44918\,
            in2 => \_gnd_net_\,
            in3 => \N__36133\,
            lcout => rand_data_15,
            ltout => OPEN,
            carryin => n15542,
            carryout => n15543,
            clk => \N__50543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i16_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41733\,
            in2 => \_gnd_net_\,
            in3 => \N__36187\,
            lcout => rand_data_16,
            ltout => OPEN,
            carryin => \bfn_13_27_0_\,
            carryout => n15544,
            clk => \N__50551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i17_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39358\,
            in2 => \_gnd_net_\,
            in3 => \N__36184\,
            lcout => rand_data_17,
            ltout => OPEN,
            carryin => n15544,
            carryout => n15545,
            clk => \N__50551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i18_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44462\,
            in2 => \_gnd_net_\,
            in3 => \N__36181\,
            lcout => rand_data_18,
            ltout => OPEN,
            carryin => n15545,
            carryout => n15546,
            clk => \N__50551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i19_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36708\,
            in2 => \_gnd_net_\,
            in3 => \N__36178\,
            lcout => rand_data_19,
            ltout => OPEN,
            carryin => n15546,
            carryout => n15547,
            clk => \N__50551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i20_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39073\,
            in2 => \_gnd_net_\,
            in3 => \N__36175\,
            lcout => rand_data_20,
            ltout => OPEN,
            carryin => n15547,
            carryout => n15548,
            clk => \N__50551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i21_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40618\,
            in2 => \_gnd_net_\,
            in3 => \N__36172\,
            lcout => rand_data_21,
            ltout => OPEN,
            carryin => n15548,
            carryout => n15549,
            clk => \N__50551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i22_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41185\,
            in2 => \_gnd_net_\,
            in3 => \N__36169\,
            lcout => rand_data_22,
            ltout => OPEN,
            carryin => n15549,
            carryout => n15550,
            clk => \N__50551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i23_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44068\,
            in2 => \_gnd_net_\,
            in3 => \N__36166\,
            lcout => rand_data_23,
            ltout => OPEN,
            carryin => n15550,
            carryout => n15551,
            clk => \N__50551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i24_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44761\,
            in2 => \_gnd_net_\,
            in3 => \N__36163\,
            lcout => rand_data_24,
            ltout => OPEN,
            carryin => \bfn_13_28_0_\,
            carryout => n15552,
            clk => \N__50561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i25_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44666\,
            in2 => \_gnd_net_\,
            in3 => \N__36292\,
            lcout => rand_data_25,
            ltout => OPEN,
            carryin => n15552,
            carryout => n15553,
            clk => \N__50561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i26_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39622\,
            in2 => \_gnd_net_\,
            in3 => \N__36289\,
            lcout => rand_data_26,
            ltout => OPEN,
            carryin => n15553,
            carryout => n15554,
            clk => \N__50561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i27_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37936\,
            in2 => \_gnd_net_\,
            in3 => \N__36286\,
            lcout => rand_data_27,
            ltout => OPEN,
            carryin => n15554,
            carryout => n15555,
            clk => \N__50561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i28_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39198\,
            in2 => \_gnd_net_\,
            in3 => \N__36283\,
            lcout => rand_data_28,
            ltout => OPEN,
            carryin => n15555,
            carryout => n15556,
            clk => \N__50561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i29_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45279\,
            in2 => \_gnd_net_\,
            in3 => \N__36280\,
            lcout => rand_data_29,
            ltout => OPEN,
            carryin => n15556,
            carryout => n15557,
            clk => \N__50561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i30_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48912\,
            in2 => \_gnd_net_\,
            in3 => \N__36277\,
            lcout => rand_data_30,
            ltout => OPEN,
            carryin => n15557,
            carryout => n15558,
            clk => \N__50561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2350__i31_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43990\,
            in2 => \_gnd_net_\,
            in3 => \N__36274\,
            lcout => rand_data_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i0_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39532\,
            in2 => \N__36267\,
            in3 => \_gnd_net_\,
            lcout => rand_setpoint_0,
            ltout => OPEN,
            carryin => \bfn_13_29_0_\,
            carryout => n15559,
            clk => \N__50571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i1_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36232\,
            in2 => \N__40569\,
            in3 => \N__36190\,
            lcout => rand_setpoint_1,
            ltout => OPEN,
            carryin => n15559,
            carryout => n15560,
            clk => \N__50571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i2_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36424\,
            in2 => \N__38163\,
            in3 => \N__36394\,
            lcout => rand_setpoint_2,
            ltout => OPEN,
            carryin => n15560,
            carryout => n15561,
            clk => \N__50571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i3_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49784\,
            in2 => \N__36391\,
            in3 => \N__36376\,
            lcout => rand_setpoint_3,
            ltout => OPEN,
            carryin => n15561,
            carryout => n15562,
            clk => \N__50571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i4_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37354\,
            in2 => \N__36373\,
            in3 => \N__36358\,
            lcout => rand_setpoint_4,
            ltout => OPEN,
            carryin => n15562,
            carryout => n15563,
            clk => \N__50571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i5_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41465\,
            in2 => \N__40104\,
            in3 => \N__36355\,
            lcout => rand_setpoint_5,
            ltout => OPEN,
            carryin => n15563,
            carryout => n15564,
            clk => \N__50571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i6_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49897\,
            in2 => \N__40044\,
            in3 => \N__36352\,
            lcout => rand_setpoint_6,
            ltout => OPEN,
            carryin => n15564,
            carryout => n15565,
            clk => \N__50571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i7_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38205\,
            in2 => \N__51327\,
            in3 => \N__36349\,
            lcout => rand_setpoint_7,
            ltout => OPEN,
            carryin => n15565,
            carryout => n15566,
            clk => \N__50571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i8_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48744\,
            in2 => \N__36339\,
            in3 => \N__36322\,
            lcout => rand_setpoint_8,
            ltout => OPEN,
            carryin => \bfn_13_30_0_\,
            carryout => n15567,
            clk => \N__50579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i9_LC_13_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37901\,
            in2 => \N__36312\,
            in3 => \N__36295\,
            lcout => rand_setpoint_9,
            ltout => OPEN,
            carryin => n15567,
            carryout => n15568,
            clk => \N__50579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i10_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36609\,
            in2 => \N__46017\,
            in3 => \N__36565\,
            lcout => rand_setpoint_10,
            ltout => OPEN,
            carryin => n15568,
            carryout => n15569,
            clk => \N__50579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i11_LC_13_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48828\,
            in2 => \N__36555\,
            in3 => \N__36538\,
            lcout => rand_setpoint_11,
            ltout => OPEN,
            carryin => n15569,
            carryout => n15570,
            clk => \N__50579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i12_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36528\,
            in2 => \N__44164\,
            in3 => \N__36517\,
            lcout => rand_setpoint_12,
            ltout => OPEN,
            carryin => n15570,
            carryout => n15571,
            clk => \N__50579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i13_LC_13_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36507\,
            in2 => \N__44566\,
            in3 => \N__36496\,
            lcout => rand_setpoint_13,
            ltout => OPEN,
            carryin => n15571,
            carryout => n15572,
            clk => \N__50579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i14_LC_13_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49095\,
            in2 => \N__36492\,
            in3 => \N__36475\,
            lcout => rand_setpoint_14,
            ltout => OPEN,
            carryin => n15572,
            carryout => n15573,
            clk => \N__50579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i15_LC_13_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36465\,
            in2 => \N__44943\,
            in3 => \N__36454\,
            lcout => rand_setpoint_15,
            ltout => OPEN,
            carryin => n15573,
            carryout => n15574,
            clk => \N__50579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i16_LC_13_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41752\,
            in2 => \N__42882\,
            in3 => \N__36451\,
            lcout => rand_setpoint_16,
            ltout => OPEN,
            carryin => \bfn_13_31_0_\,
            carryout => n15575,
            clk => \N__50585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i17_LC_13_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39374\,
            in2 => \N__38272\,
            in3 => \N__36448\,
            lcout => rand_setpoint_17,
            ltout => OPEN,
            carryin => n15575,
            carryout => n15576,
            clk => \N__50585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i18_LC_13_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44470\,
            in2 => \N__38299\,
            in3 => \N__36445\,
            lcout => rand_setpoint_18,
            ltout => OPEN,
            carryin => n15576,
            carryout => n15577,
            clk => \N__50585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i19_LC_13_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36718\,
            in2 => \N__38332\,
            in3 => \N__36679\,
            lcout => rand_setpoint_19,
            ltout => OPEN,
            carryin => n15577,
            carryout => n15578,
            clk => \N__50585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i20_LC_13_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39082\,
            in2 => \N__38362\,
            in3 => \N__36676\,
            lcout => rand_setpoint_20,
            ltout => OPEN,
            carryin => n15578,
            carryout => n15579,
            clk => \N__50585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i21_LC_13_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40634\,
            in2 => \N__46518\,
            in3 => \N__36673\,
            lcout => rand_setpoint_21,
            ltout => OPEN,
            carryin => n15579,
            carryout => n15580,
            clk => \N__50585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i22_LC_13_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41203\,
            in2 => \N__36670\,
            in3 => \N__36655\,
            lcout => rand_setpoint_22,
            ltout => OPEN,
            carryin => n15580,
            carryout => n15581,
            clk => \N__50585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i23_LC_13_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44081\,
            in2 => \N__40290\,
            in3 => \N__36652\,
            lcout => rand_setpoint_23,
            ltout => OPEN,
            carryin => n15581,
            carryout => n15582,
            clk => \N__50585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i24_LC_13_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44782\,
            in2 => \N__38224\,
            in3 => \N__36649\,
            lcout => rand_setpoint_24,
            ltout => OPEN,
            carryin => \bfn_13_32_0_\,
            carryout => n15583,
            clk => \N__50589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i25_LC_13_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44686\,
            in2 => \N__36646\,
            in3 => \N__36631\,
            lcout => rand_setpoint_25,
            ltout => OPEN,
            carryin => n15583,
            carryout => n15584,
            clk => \N__50589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i26_LC_13_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38253\,
            in2 => \N__39636\,
            in3 => \N__36628\,
            lcout => rand_setpoint_26,
            ltout => OPEN,
            carryin => n15584,
            carryout => n15585,
            clk => \N__50589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i27_LC_13_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37945\,
            in2 => \N__38641\,
            in3 => \N__36625\,
            lcout => rand_setpoint_27,
            ltout => OPEN,
            carryin => n15585,
            carryout => n15586,
            clk => \N__50589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i28_LC_13_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39202\,
            in2 => \N__38626\,
            in3 => \N__36877\,
            lcout => rand_setpoint_28,
            ltout => OPEN,
            carryin => n15586,
            carryout => n15587,
            clk => \N__50589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i29_LC_13_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45292\,
            in2 => \N__38241\,
            in3 => \N__36874\,
            lcout => rand_setpoint_29,
            ltout => OPEN,
            carryin => n15587,
            carryout => n15588,
            clk => \N__50589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i30_LC_13_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48934\,
            in2 => \N__36871\,
            in3 => \N__36856\,
            lcout => rand_setpoint_30,
            ltout => OPEN,
            carryin => n15588,
            carryout => n15589,
            clk => \N__50589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2351__i31_LC_13_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44002\,
            in1 => \N__36850\,
            in2 => \_gnd_net_\,
            in3 => \N__36853\,
            lcout => rand_setpoint_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_537_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52513\,
            in1 => \N__40351\,
            in2 => \_gnd_net_\,
            in3 => \N__36838\,
            lcout => \c0.n17064\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__47821\,
            in1 => \N__48955\,
            in2 => \N__38791\,
            in3 => \N__47659\,
            lcout => OPEN,
            ltout => \c0.n22_adj_2357_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i3_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__51609\,
            in1 => \N__36769\,
            in2 => \N__36796\,
            in3 => \N__51738\,
            lcout => \c0.tx2.r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50468\,
            ce => \N__51447\,
            sr => \_gnd_net_\
        );

    \c0.n18125_bdd_4_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__38386\,
            in1 => \N__36781\,
            in2 => \N__40744\,
            in3 => \N__51608\,
            lcout => \c0.n18128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_644_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40799\,
            in1 => \N__49198\,
            in2 => \N__36763\,
            in3 => \N__41242\,
            lcout => \c0.n18_adj_2331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_573_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49557\,
            in1 => \N__43465\,
            in2 => \_gnd_net_\,
            in3 => \N__37149\,
            lcout => \c0.n17100\,
            ltout => \c0.n17100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36955\,
            in3 => \N__41934\,
            lcout => OPEN,
            ltout => \c0.n16_adj_2332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i153_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38419\,
            in1 => \N__37195\,
            in2 => \N__36952\,
            in3 => \N__36949\,
            lcout => \c0.data_out_frame2_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50481\,
            ce => \N__51185\,
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_481_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39670\,
            in1 => \N__43189\,
            in2 => \N__42010\,
            in3 => \N__39496\,
            lcout => OPEN,
            ltout => \c0.n12_adj_2263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i163_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36928\,
            in1 => \N__41068\,
            in2 => \N__36922\,
            in3 => \N__38833\,
            lcout => \c0.data_out_frame2_20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50493\,
            ce => \N__51182\,
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_590_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39435\,
            in1 => \N__37588\,
            in2 => \N__37054\,
            in3 => \N__37624\,
            lcout => OPEN,
            ltout => \c0.n16_adj_2312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i157_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36907\,
            in1 => \N__36888\,
            in2 => \N__36895\,
            in3 => \N__38401\,
            lcout => \c0.data_out_frame2_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50493\,
            ce => \N__51182\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_584_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43309\,
            in2 => \_gnd_net_\,
            in3 => \N__39669\,
            lcout => \c0.n17097\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39668\,
            in1 => \N__48092\,
            in2 => \_gnd_net_\,
            in3 => \N__37147\,
            lcout => \c0.n5_adj_2334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_480_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37117\,
            in1 => \N__38541\,
            in2 => \N__49476\,
            in3 => \N__38976\,
            lcout => \c0.n17052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37737\,
            in1 => \N__40148\,
            in2 => \N__37077\,
            in3 => \N__49015\,
            lcout => \c0.n20_adj_2202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_593_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__37042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38462\,
            lcout => \c0.n9839\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41110\,
            in1 => \N__43524\,
            in2 => \_gnd_net_\,
            in3 => \N__38679\,
            lcout => \c0.n14_adj_2264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17957_bdd_4_lut_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__48512\,
            in1 => \N__37156\,
            in2 => \N__37305\,
            in3 => \N__40725\,
            lcout => \c0.n17960\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_490_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37041\,
            in2 => \_gnd_net_\,
            in3 => \N__44434\,
            lcout => \c0.n17031\,
            ltout => \c0.n17031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_493_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37003\,
            in1 => \N__37692\,
            in2 => \N__36991\,
            in3 => \N__37264\,
            lcout => \c0.n26_adj_2273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_447_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38773\,
            in1 => \N__45628\,
            in2 => \_gnd_net_\,
            in3 => \N__36988\,
            lcout => \c0.n17085\,
            ltout => \c0.n17085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_445_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37309\,
            in1 => \N__44307\,
            in2 => \N__37267\,
            in3 => \N__37263\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15523_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__37243\,
            in1 => \N__48142\,
            in2 => \N__48583\,
            in3 => \N__37222\,
            lcout => \c0.n17969\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_607_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37849\,
            in1 => \N__37174\,
            in2 => \_gnd_net_\,
            in3 => \N__37213\,
            lcout => \c0.n17088\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_606_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45363\,
            in1 => \N__37191\,
            in2 => \N__49290\,
            in3 => \N__41160\,
            lcout => \c0.n9579\,
            ltout => \c0.n9579_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_579_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38774\,
            in2 => \N__37168\,
            in3 => \_gnd_net_\,
            lcout => \c0.n10_adj_2307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15621_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__38892\,
            in1 => \N__48141\,
            in2 => \N__48582\,
            in3 => \N__41159\,
            lcout => \c0.n18071\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15514_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__48140\,
            in1 => \N__41831\,
            in2 => \N__48581\,
            in3 => \N__41263\,
            lcout => \c0.n17957\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i90_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41535\,
            in1 => \N__50936\,
            in2 => \_gnd_net_\,
            in3 => \N__37910\,
            lcout => data_out_frame2_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i68_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50932\,
            in1 => \N__49802\,
            in2 => \_gnd_net_\,
            in3 => \N__40724\,
            lcout => data_out_frame2_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i81_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41753\,
            in1 => \N__50935\,
            in2 => \_gnd_net_\,
            in3 => \N__43572\,
            lcout => data_out_frame2_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_525_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41534\,
            in2 => \_gnd_net_\,
            in3 => \N__40860\,
            lcout => \c0.n16908\,
            ltout => \c0.n16908_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_475_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49698\,
            in1 => \N__38890\,
            in2 => \N__37597\,
            in3 => \N__41264\,
            lcout => \c0.n17022\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_684_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39275\,
            in1 => \N__39128\,
            in2 => \_gnd_net_\,
            in3 => \N__49423\,
            lcout => \c0.n6_adj_2286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i104_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__51328\,
            in1 => \N__50934\,
            in2 => \_gnd_net_\,
            in3 => \N__43756\,
            lcout => data_out_frame2_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i92_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50933\,
            in1 => \_gnd_net_\,
            in2 => \N__41269\,
            in3 => \N__48829\,
            lcout => data_out_frame2_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i117_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39090\,
            in1 => \N__37579\,
            in2 => \_gnd_net_\,
            in3 => \N__51104\,
            lcout => data_out_frame2_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15414_3_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__37555\,
            in1 => \N__37453\,
            in2 => \_gnd_net_\,
            in3 => \N__37383\,
            lcout => n10197,
            ltout => \n10197_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i69_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__37349\,
            in1 => \_gnd_net_\,
            in2 => \N__37312\,
            in3 => \N__49324\,
            lcout => data_out_frame2_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i82_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51102\,
            in1 => \N__39368\,
            in2 => \_gnd_net_\,
            in3 => \N__47409\,
            lcout => data_out_frame2_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i119_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41204\,
            in1 => \N__43678\,
            in2 => \_gnd_net_\,
            in3 => \N__51105\,
            lcout => data_out_frame2_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_575_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__49323\,
            in1 => \N__37766\,
            in2 => \N__39495\,
            in3 => \_gnd_net_\,
            lcout => \c0.n9749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i102_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37732\,
            in1 => \N__41454\,
            in2 => \_gnd_net_\,
            in3 => \N__51103\,
            lcout => data_out_frame2_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_629_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40774\,
            in1 => \N__41859\,
            in2 => \N__43267\,
            in3 => \N__41689\,
            lcout => \c0.n17049\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i75_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39635\,
            in1 => \N__43884\,
            in2 => \_gnd_net_\,
            in3 => \N__50927\,
            lcout => data_out_frame2_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15224_3_lut_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__48165\,
            in1 => \N__49536\,
            in2 => \_gnd_net_\,
            in3 => \N__48585\,
            lcout => \c0.n17561\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_631_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49535\,
            in2 => \_gnd_net_\,
            in3 => \N__48705\,
            lcout => \c0.n9589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i43_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50925\,
            in1 => \N__39634\,
            in2 => \_gnd_net_\,
            in3 => \N__37651\,
            lcout => data_out_frame2_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_576_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37623\,
            in2 => \_gnd_net_\,
            in3 => \N__39038\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_577_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38893\,
            in1 => \N__45248\,
            in2 => \N__37960\,
            in3 => \N__49503\,
            lcout => \c0.n16987\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i42_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44687\,
            in1 => \N__39013\,
            in2 => \_gnd_net_\,
            in3 => \N__50926\,
            lcout => data_out_frame2_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i108_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__37946\,
            in1 => \N__39274\,
            in2 => \N__51246\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_444_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43682\,
            in2 => \_gnd_net_\,
            in3 => \N__48706\,
            lcout => \c0.n10_adj_2191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i138_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__37897\,
            in1 => \N__37863\,
            in2 => \N__51247\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_17_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i85_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51161\,
            in2 => \N__39083\,
            in3 => \N__37837\,
            lcout => data_out_frame2_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i168_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41608\,
            in1 => \N__43766\,
            in2 => \N__37807\,
            in3 => \N__37798\,
            lcout => \c0.data_out_frame2_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50562\,
            ce => \N__51181\,
            sr => \_gnd_net_\
        );

    \c0.i15256_3_lut_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__42396\,
            in1 => \N__42754\,
            in2 => \_gnd_net_\,
            in3 => \N__40228\,
            lcout => \c0.n17528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15245_3_lut_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__45205\,
            in1 => \_gnd_net_\,
            in2 => \N__42763\,
            in3 => \N__52140\,
            lcout => \c0.n17507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__2__2162_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38107\,
            in1 => \N__46803\,
            in2 => \N__38065\,
            in3 => \N__46911\,
            lcout => \c0.data_out_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50572\,
            ce => \N__46620\,
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_533_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39957\,
            in1 => \N__39721\,
            in2 => \N__38064\,
            in3 => \N__42464\,
            lcout => OPEN,
            ltout => \c0.n12_adj_2289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__1__2163_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46697\,
            in1 => \N__47140\,
            in2 => \N__38041\,
            in3 => \N__39730\,
            lcout => \c0.data_out_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50572\,
            ce => \N__46620\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__0__2164_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38038\,
            in1 => \N__42288\,
            in2 => \N__42217\,
            in3 => \N__39729\,
            lcout => \c0.data_out_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50572\,
            ce => \N__46620\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_524_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39832\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39898\,
            lcout => \c0.n9496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_494_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40479\,
            in2 => \_gnd_net_\,
            in3 => \N__40025\,
            lcout => \c0.n6_adj_2274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40024\,
            in1 => \N__40077\,
            in2 => \_gnd_net_\,
            in3 => \N__52136\,
            lcout => \c0.n9716\,
            ltout => \c0.n9716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_693_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46739\,
            in1 => \N__52544\,
            in2 => \N__37996\,
            in3 => \N__37989\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46646\,
            in1 => \N__45201\,
            in2 => \N__37975\,
            in3 => \N__45106\,
            lcout => \data_out_9__2__N_367\,
            ltout => \data_out_9__2__N_367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_686_LC_14_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__39899\,
            in1 => \_gnd_net_\,
            in2 => \N__37963\,
            in3 => \N__39833\,
            lcout => \c0.n17094\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_648_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39813\,
            in1 => \N__40057\,
            in2 => \N__40413\,
            in3 => \N__46863\,
            lcout => \c0.n16998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__7__2173_LC_14_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__45107\,
            in1 => \N__42745\,
            in2 => \N__38209\,
            in3 => \N__42838\,
            lcout => data_out_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52091\,
            in1 => \N__46798\,
            in2 => \_gnd_net_\,
            in3 => \N__40023\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2169_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__52301\,
            in1 => \N__46647\,
            in2 => \N__38194\,
            in3 => \N__52092\,
            lcout => n10_adj_2427,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_484_LC_14_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46200\,
            in1 => \N__38179\,
            in2 => \N__38173\,
            in3 => \N__40269\,
            lcout => \c0.n10_adj_2268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__2__2178_LC_14_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__42847\,
            in1 => \N__42760\,
            in2 => \N__38164\,
            in3 => \N__39875\,
            lcout => \c0.data_out_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15347_2_lut_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52090\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38115\,
            lcout => \c0.n17594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_14_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45099\,
            in1 => \N__46969\,
            in2 => \_gnd_net_\,
            in3 => \N__52089\,
            lcout => \c0.n8_adj_2176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__2__2234_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__46488\,
            in1 => \N__38116\,
            in2 => \N__46138\,
            in3 => \N__42727\,
            lcout => \c0.data_out_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__7__2221_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011011100"
        )
    port map (
            in0 => \N__45455\,
            in1 => \N__38379\,
            in2 => \N__46000\,
            in3 => \N__46489\,
            lcout => data_out_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__4__2192_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38361\,
            in1 => \N__45803\,
            in2 => \N__38347\,
            in3 => \N__46420\,
            lcout => \c0.data_out_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50590\,
            ce => \N__46130\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__3__2193_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46417\,
            in1 => \N__38331\,
            in2 => \N__38317\,
            in3 => \N__45874\,
            lcout => \c0.data_out_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50590\,
            ce => \N__46130\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__2__2194_LC_14_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38298\,
            in1 => \N__45802\,
            in2 => \N__38284\,
            in3 => \N__46419\,
            lcout => \c0.data_out_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50590\,
            ce => \N__46130\,
            sr => \_gnd_net_\
        );

    \c0.i15246_2_lut_LC_14_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45801\,
            in1 => \N__38271\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n17506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__1__2195_LC_14_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111010001"
        )
    port map (
            in0 => \N__42758\,
            in1 => \N__46418\,
            in2 => \N__38257\,
            in3 => \N__52135\,
            lcout => \c0.data_out_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50590\,
            ce => \N__46130\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__2__2202_LC_14_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45994\,
            in1 => \N__38254\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50595\,
            ce => \N__46129\,
            sr => \N__41889\
        );

    \c0.data_out_5__5__2199_LC_14_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38242\,
            in3 => \N__45992\,
            lcout => \c0.data_out_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50595\,
            ce => \N__46129\,
            sr => \N__41889\
        );

    \c0.data_out_5__0__2204_LC_14_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45993\,
            in1 => \N__38223\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_6__1__N_537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50595\,
            ce => \N__46129\,
            sr => \N__41889\
        );

    \c0.data_out_5__3__2201_LC_14_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45991\,
            in2 => \_gnd_net_\,
            in3 => \N__38640\,
            lcout => \c0.data_out_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50595\,
            ce => \N__46129\,
            sr => \N__41889\
        );

    \c0.data_out_5__4__2200_LC_14_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45995\,
            in1 => \N__38625\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50595\,
            ce => \N__46129\,
            sr => \N__41889\
        );

    \c0.i1_2_lut_adj_574_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38611\,
            in2 => \_gnd_net_\,
            in3 => \N__38581\,
            lcout => \c0.n9763\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_639_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39333\,
            in2 => \_gnd_net_\,
            in3 => \N__38523\,
            lcout => \c0.n17037\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_541_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39442\,
            in1 => \N__38485\,
            in2 => \N__40692\,
            in3 => \N__43523\,
            lcout => \c0.n17040\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_586_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42331\,
            in2 => \_gnd_net_\,
            in3 => \N__38469\,
            lcout => \c0.n16933\,
            ltout => \c0.n16933_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_591_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38415\,
            in1 => \N__38862\,
            in2 => \N__38404\,
            in3 => \N__44242\,
            lcout => \c0.n17_adj_2313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__38395\,
            in1 => \N__51643\,
            in2 => \N__39244\,
            in3 => \N__47674\,
            lcout => \c0.n18125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_611_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43216\,
            in1 => \N__44441\,
            in2 => \N__38986\,
            in3 => \N__39593\,
            lcout => OPEN,
            ltout => \c0.n15_adj_2320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i155_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__38839\,
            in1 => \N__38935\,
            in2 => \N__38866\,
            in3 => \N__38863\,
            lcout => \c0.data_out_frame2_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50504\,
            ce => \N__51168\,
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_674_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43463\,
            in1 => \N__47200\,
            in2 => \N__47320\,
            in3 => \N__49345\,
            lcout => \c0.n14_adj_2323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_474_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38832\,
            in1 => \N__47505\,
            in2 => \N__38821\,
            in3 => \N__40654\,
            lcout => OPEN,
            ltout => \c0.n21_adj_2255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i164_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__38806\,
            in1 => \_gnd_net_\,
            in2 => \N__38794\,
            in3 => \N__41788\,
            lcout => \c0.data_out_frame2_20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50504\,
            ce => \N__51168\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i118_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40641\,
            in1 => \N__38775\,
            in2 => \_gnd_net_\,
            in3 => \N__51001\,
            lcout => data_out_frame2_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50515\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_478_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42327\,
            in2 => \_gnd_net_\,
            in3 => \N__38751\,
            lcout => \c0.n9555\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_503_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38734\,
            in1 => \N__43318\,
            in2 => \N__38728\,
            in3 => \N__39385\,
            lcout => \c0.n17103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38668\,
            in1 => \N__41487\,
            in2 => \N__47484\,
            in3 => \N__38650\,
            lcout => \c0.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_569_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39048\,
            in1 => \N__39022\,
            in2 => \N__41413\,
            in3 => \N__47376\,
            lcout => \c0.n19_adj_2303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_609_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41872\,
            in2 => \_gnd_net_\,
            in3 => \N__43278\,
            lcout => \c0.n9776\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_465_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43411\,
            in1 => \N__38977\,
            in2 => \N__43795\,
            in3 => \N__39494\,
            lcout => OPEN,
            ltout => \c0.n22_adj_2207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i165_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41379\,
            in1 => \N__38965\,
            in2 => \N__38953\,
            in3 => \N__38950\,
            lcout => \c0.data_out_frame2_20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50524\,
            ce => \N__50995\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_603_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41135\,
            in2 => \_gnd_net_\,
            in3 => \N__42073\,
            lcout => \c0.n9892\,
            ltout => \c0.n9892_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_682_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39133\,
            in1 => \N__49427\,
            in2 => \N__38938\,
            in3 => \N__44241\,
            lcout => \c0.n17079\,
            ltout => \c0.n17079_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i166_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__38926\,
            in1 => \N__41488\,
            in2 => \N__38917\,
            in3 => \N__38914\,
            lcout => \c0.data_out_frame2_20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50524\,
            ce => \N__50995\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i94_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50944\,
            in1 => \N__44568\,
            in2 => \_gnd_net_\,
            in3 => \N__41136\,
            lcout => data_out_frame2_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i88_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44092\,
            in1 => \N__38891\,
            in2 => \_gnd_net_\,
            in3 => \N__50947\,
            lcout => data_out_frame2_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i45_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50942\,
            in1 => \N__39214\,
            in2 => \_gnd_net_\,
            in3 => \N__43519\,
            lcout => data_out_frame2_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i79_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48936\,
            in1 => \N__43472\,
            in2 => \_gnd_net_\,
            in3 => \N__50946\,
            lcout => data_out_frame2_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_597_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39163\,
            in1 => \N__39277\,
            in2 => \_gnd_net_\,
            in3 => \N__39132\,
            lcout => \c0.n17082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i96_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44946\,
            in1 => \N__41161\,
            in2 => \_gnd_net_\,
            in3 => \N__50948\,
            lcout => data_out_frame2_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i55_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50943\,
            in1 => \_gnd_net_\,
            in2 => \N__41217\,
            in3 => \N__43266\,
            lcout => data_out_frame2_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i126_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44567\,
            in1 => \N__49735\,
            in2 => \_gnd_net_\,
            in3 => \N__50945\,
            lcout => data_out_frame2_15_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i50_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39376\,
            in1 => \N__50930\,
            in2 => \_gnd_net_\,
            in3 => \N__41514\,
            lcout => data_out_frame2_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i53_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50928\,
            in1 => \_gnd_net_\,
            in2 => \N__39094\,
            in3 => \N__39326\,
            lcout => data_out_frame2_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i61_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__41041\,
            in1 => \N__50931\,
            in2 => \N__44173\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_498_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39434\,
            in1 => \N__39396\,
            in2 => \N__47312\,
            in3 => \N__49227\,
            lcout => \c0.n25_adj_2275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i114_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39375\,
            in1 => \N__50929\,
            in2 => \_gnd_net_\,
            in3 => \N__49459\,
            lcout => data_out_frame2_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48120\,
            in1 => \N__41040\,
            in2 => \_gnd_net_\,
            in3 => \N__39325\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_15582_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__48630\,
            in1 => \N__43489\,
            in2 => \N__39304\,
            in3 => \N__47705\,
            lcout => \c0.n17987\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17951_bdd_4_lut_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__48568\,
            in1 => \N__39289\,
            in2 => \N__45361\,
            in3 => \N__39276\,
            lcout => \c0.n17954\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i70_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41464\,
            in1 => \N__41867\,
            in2 => \_gnd_net_\,
            in3 => \N__50952\,
            lcout => data_out_frame2_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i74_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50950\,
            in1 => \_gnd_net_\,
            in2 => \N__44694\,
            in3 => \N__41696\,
            lcout => data_out_frame2_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14884_3_lut_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41956\,
            in1 => \N__48187\,
            in2 => \_gnd_net_\,
            in3 => \N__47372\,
            lcout => \c0.n17322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18053_bdd_4_lut_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47715\,
            in1 => \N__39646\,
            in2 => \N__41764\,
            in3 => \N__43537\,
            lcout => \c0.n18056\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i57_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50949\,
            in1 => \N__48768\,
            in2 => \_gnd_net_\,
            in3 => \N__39660\,
            lcout => data_out_frame2_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i105_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41957\,
            in1 => \N__44784\,
            in2 => \_gnd_net_\,
            in3 => \N__50951\,
            lcout => data_out_frame2_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14908_3_lut_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48164\,
            in1 => \N__49415\,
            in2 => \_gnd_net_\,
            in3 => \N__39477\,
            lcout => \c0.n17346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i107_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39637\,
            in1 => \N__43372\,
            in2 => \_gnd_net_\,
            in3 => \N__51192\,
            lcout => data_out_frame2_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_558_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42205\,
            in2 => \_gnd_net_\,
            in3 => \N__46199\,
            lcout => \c0.n16918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i115_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44480\,
            in1 => \N__39576\,
            in2 => \_gnd_net_\,
            in3 => \N__51193\,
            lcout => data_out_frame2_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i65_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49416\,
            in1 => \N__39546\,
            in2 => \_gnd_net_\,
            in3 => \N__51194\,
            lcout => data_out_frame2_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i73_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51191\,
            in1 => \N__44783\,
            in2 => \_gnd_net_\,
            in3 => \N__39478\,
            lcout => data_out_frame2_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i78_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45293\,
            in1 => \N__44842\,
            in2 => \_gnd_net_\,
            in3 => \N__51195\,
            lcout => data_out_frame2_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__7__2157_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47023\,
            in1 => \N__46968\,
            in2 => \N__42982\,
            in3 => \N__39454\,
            lcout => \c0.data_out_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50573\,
            ce => \N__46616\,
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_523_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47096\,
            in1 => \N__39812\,
            in2 => \N__39782\,
            in3 => \N__40056\,
            lcout => \c0.n16966\,
            ltout => \c0.n16966_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_530_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46967\,
            in1 => \N__45000\,
            in2 => \N__39745\,
            in3 => \N__46791\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_531_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39742\,
            in1 => \N__45144\,
            in2 => \N__39733\,
            in3 => \N__47004\,
            lcout => \c0.n17109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_552_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39720\,
            in2 => \_gnd_net_\,
            in3 => \N__39934\,
            lcout => \c0.n17070\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52066\,
            in1 => \N__45022\,
            in2 => \_gnd_net_\,
            in3 => \N__43020\,
            lcout => \c0.n8_adj_2153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_545_LC_15_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39704\,
            in2 => \_gnd_net_\,
            in3 => \N__46966\,
            lcout => \c0.n17007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_688_LC_15_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40079\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40026\,
            lcout => \c0.n16949\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39932\,
            in1 => \N__40078\,
            in2 => \_gnd_net_\,
            in3 => \N__52082\,
            lcout => \c0.n8_adj_2166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__45930\,
            in1 => \N__42647\,
            in2 => \_gnd_net_\,
            in3 => \N__46475\,
            lcout => n4445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__5__2175_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__42648\,
            in1 => \N__40105\,
            in2 => \N__42860\,
            in3 => \N__40080\,
            lcout => data_out_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_509_LC_15_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42402\,
            in1 => \N__39933\,
            in2 => \N__40429\,
            in3 => \N__42466\,
            lcout => \c0.n19_adj_2283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_557_LC_15_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39858\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43013\,
            lcout => \c0.n28_adj_2287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__6__2174_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__40045\,
            in1 => \N__42842\,
            in2 => \N__42708\,
            in3 => \N__40027\,
            lcout => data_out_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_529_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46822\,
            in1 => \N__39993\,
            in2 => \_gnd_net_\,
            in3 => \N__40425\,
            lcout => \c0.n17043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__52088\,
            in1 => \N__39976\,
            in2 => \N__39838\,
            in3 => \N__52288\,
            lcout => n10_adj_2425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__5__2167_LC_15_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39837\,
            in1 => \N__39958\,
            in2 => \N__44973\,
            in3 => \N__40552\,
            lcout => \c0.data_out_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50591\,
            ce => \N__46606\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__5__2159_LC_15_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42253\,
            in1 => \N__42202\,
            in2 => \N__39916\,
            in3 => \N__39876\,
            lcout => \c0.data_out_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50591\,
            ce => \N__46606\,
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_553_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42228\,
            in1 => \N__40455\,
            in2 => \N__45214\,
            in3 => \N__52131\,
            lcout => \c0.n17025\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__1__2179_LC_15_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__40385\,
            in1 => \N__40573\,
            in2 => \N__42862\,
            in3 => \N__42759\,
            lcout => data_out_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_521_LC_15_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40551\,
            in1 => \N__40259\,
            in2 => \N__40525\,
            in3 => \N__40454\,
            lcout => \c0.n9522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__40384\,
            in1 => \N__43112\,
            in2 => \N__52081\,
            in3 => \N__42921\,
            lcout => \c0.n18077\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15213_3_lut_4_lut_LC_15_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__42653\,
            in1 => \N__40340\,
            in2 => \N__40188\,
            in3 => \N__45075\,
            lcout => OPEN,
            ltout => \c0.n17532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__7__2189_LC_15_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__40294\,
            in1 => \N__45996\,
            in2 => \N__40273\,
            in3 => \N__46490\,
            lcout => \c0.data_out_6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50599\,
            ce => \N__46128\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_538_LC_15_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42439\,
            in2 => \_gnd_net_\,
            in3 => \N__42371\,
            lcout => \c0.n9737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15255_3_lut_4_lut_LC_15_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__42652\,
            in1 => \N__40219\,
            in2 => \N__40187\,
            in3 => \N__45074\,
            lcout => \c0.n17534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15543_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__40669\,
            in1 => \N__48535\,
            in2 => \N__40924\,
            in3 => \N__48105\,
            lcout => \c0.n17999\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15284_3_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__40153\,
            in1 => \N__48624\,
            in2 => \_gnd_net_\,
            in3 => \N__48106\,
            lcout => \c0.n17576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_628_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41347\,
            in1 => \N__44200\,
            in2 => \_gnd_net_\,
            in3 => \N__40729\,
            lcout => \c0.n9826\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_608_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43848\,
            in1 => \N__43373\,
            in2 => \N__49855\,
            in3 => \N__49379\,
            lcout => \c0.n17016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_601_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43231\,
            in1 => \N__44044\,
            in2 => \N__40696\,
            in3 => \N__44887\,
            lcout => \c0.n25_adj_2316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i151_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__49917\,
            in1 => \N__40668\,
            in2 => \N__51248\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_621_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41832\,
            in2 => \_gnd_net_\,
            in3 => \N__44632\,
            lcout => \c0.n9843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_516_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43959\,
            lcout => \c0.n16994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i54_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51170\,
            in2 => \N__44642\,
            in3 => \N__40645\,
            lcout => data_out_frame2_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_3_lut_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44308\,
            in1 => \N__40594\,
            in2 => \_gnd_net_\,
            in3 => \N__43336\,
            lcout => OPEN,
            ltout => \c0.n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i160_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41353\,
            in1 => \N__41005\,
            in2 => \N__40582\,
            in3 => \N__40579\,
            lcout => \c0.data_out_frame2_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50525\,
            ce => \N__51169\,
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_559_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44735\,
            in1 => \N__43279\,
            in2 => \N__44443\,
            in3 => \N__49003\,
            lcout => \c0.n29_adj_2296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_598_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41596\,
            in2 => \_gnd_net_\,
            in3 => \N__44734\,
            lcout => \c0.n16915\,
            ltout => \c0.n16915_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_568_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40999\,
            in1 => \N__49629\,
            in2 => \N__40987\,
            in3 => \N__40984\,
            lcout => OPEN,
            ltout => \c0.n20_adj_2302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i159_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40942\,
            in2 => \N__40936\,
            in3 => \N__40933\,
            lcout => \c0.data_out_frame2_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50525\,
            ce => \N__51169\,
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_673_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49576\,
            in1 => \N__41074\,
            in2 => \N__44614\,
            in3 => \N__41049\,
            lcout => \c0.n16972\,
            ltout => \c0.n16972_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_505_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40912\,
            in1 => \N__49380\,
            in2 => \N__40879\,
            in3 => \N__40876\,
            lcout => \c0.n10_adj_2281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17969_bdd_4_lut_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__40813\,
            in1 => \N__40804\,
            in2 => \N__44110\,
            in3 => \N__48625\,
            lcout => OPEN,
            ltout => \c0.n17972_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__47761\,
            in1 => \N__40753\,
            in2 => \N__40747\,
            in3 => \N__47710\,
            lcout => \c0.n22_adj_2355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_555_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41380\,
            in1 => \N__43182\,
            in2 => \N__41623\,
            in3 => \N__41359\,
            lcout => \c0.n30_adj_2295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41346\,
            in1 => \N__48167\,
            in2 => \_gnd_net_\,
            in3 => \N__44040\,
            lcout => \c0.n5_adj_2351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_638_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41268\,
            in1 => \N__42068\,
            in2 => \_gnd_net_\,
            in3 => \N__47451\,
            lcout => \c0.n9695\,
            ltout => \c0.n9695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_617_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41221\,
            in3 => \N__41509\,
            lcout => \c0.n6_adj_2325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i87_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51199\,
            in1 => \N__41218\,
            in2 => \_gnd_net_\,
            in3 => \N__42316\,
            lcout => data_out_frame2_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_634_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41158\,
            in1 => \N__41131\,
            in2 => \_gnd_net_\,
            in3 => \N__44221\,
            lcout => \c0.n17019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_542_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41109\,
            in1 => \N__41086\,
            in2 => \N__41995\,
            in3 => \N__42315\,
            lcout => \c0.n10_adj_2292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6319_2_lut_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__48614\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48190\,
            lcout => \c0.n8621\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_534_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44605\,
            lcout => \c0.n9913\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i103_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49906\,
            in1 => \N__43636\,
            in2 => \_gnd_net_\,
            in3 => \N__51200\,
            lcout => data_out_frame2_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i80_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51202\,
            in1 => \N__44013\,
            in2 => \_gnd_net_\,
            in3 => \N__44878\,
            lcout => data_out_frame2_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44877\,
            in1 => \N__47410\,
            in2 => \N__44852\,
            in3 => \N__47361\,
            lcout => \c0.n17034\,
            ltout => \c0.n17034_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_615_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41611\,
            in3 => \N__41398\,
            lcout => \c0.n9688\,
            ltout => \c0.n9688_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_618_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43832\,
            in1 => \N__41595\,
            in2 => \N__41551\,
            in3 => \N__41548\,
            lcout => \c0.n17010\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i46_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51201\,
            in1 => \N__45301\,
            in2 => \_gnd_net_\,
            in3 => \N__44610\,
            lcout => data_out_frame2_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15480_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__48171\,
            in1 => \N__41542\,
            in2 => \N__48653\,
            in3 => \N__47411\,
            lcout => \c0.n17921\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_514_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41513\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45252\,
            lcout => \c0.n17115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i134_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41399\,
            in1 => \N__41469\,
            in2 => \_gnd_net_\,
            in3 => \N__51203\,
            lcout => data_out_frame2_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_600_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45348\,
            in1 => \N__41866\,
            in2 => \N__50644\,
            in3 => \N__41833\,
            lcout => \c0.n24_adj_2315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_472_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45596\,
            in1 => \N__44841\,
            in2 => \N__49156\,
            in3 => \N__42066\,
            lcout => \c0.n20_adj_2252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14885_3_lut_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49365\,
            in1 => \N__42023\,
            in2 => \_gnd_net_\,
            in3 => \N__48188\,
            lcout => OPEN,
            ltout => \c0.n17323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__48655\,
            in1 => \N__41773\,
            in2 => \N__41767\,
            in3 => \N__47714\,
            lcout => \c0.n18053\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i121_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48766\,
            in2 => \N__49378\,
            in3 => \N__51186\,
            lcout => data_out_frame2_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i113_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42024\,
            in1 => \N__41754\,
            in2 => \_gnd_net_\,
            in3 => \N__51190\,
            lcout => data_out_frame2_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17921_bdd_4_lut_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__41690\,
            in1 => \N__48654\,
            in2 => \N__47302\,
            in3 => \N__41668\,
            lcout => \c0.n17924\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i152_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51187\,
            in1 => \N__51339\,
            in2 => \_gnd_net_\,
            in3 => \N__41647\,
            lcout => data_out_frame2_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15592_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__41646\,
            in1 => \N__48651\,
            in2 => \N__41638\,
            in3 => \N__48189\,
            lcout => OPEN,
            ltout => \c0.n18059_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18059_bdd_4_lut_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48652\,
            in1 => \N__42033\,
            in2 => \N__42094\,
            in3 => \N__50637\,
            lcout => OPEN,
            ltout => \c0.n18062_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__42091\,
            in1 => \N__47787\,
            in2 => \N__42076\,
            in3 => \N__47716\,
            lcout => \c0.n22_adj_2352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i93_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51188\,
            in1 => \N__44165\,
            in2 => \_gnd_net_\,
            in3 => \N__42067\,
            lcout => data_out_frame2_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i144_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42034\,
            in1 => \N__44945\,
            in2 => \_gnd_net_\,
            in3 => \N__51189\,
            lcout => data_out_frame2_17_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_632_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42025\,
            in2 => \_gnd_net_\,
            in3 => \N__44395\,
            lcout => \c0.n9853\,
            ltout => \c0.n9853_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_633_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41994\,
            in1 => \N__49854\,
            in2 => \N__41971\,
            in3 => \N__41958\,
            lcout => \c0.n17046\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15331_2_lut_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45378\,
            in2 => \_gnd_net_\,
            in3 => \N__52096\,
            lcout => \c0.n17581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15411_2_lut_3_lut_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45931\,
            in1 => \N__45435\,
            in2 => \_gnd_net_\,
            in3 => \N__46480\,
            lcout => \c0.n10259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_16_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42289\,
            in1 => \N__42203\,
            in2 => \_gnd_net_\,
            in3 => \N__52084\,
            lcout => \c0.n5_adj_2350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_16_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__52085\,
            in1 => \N__42259\,
            in2 => \N__52300\,
            in3 => \N__46821\,
            lcout => \c0.n10_adj_2154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_515_LC_16_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42249\,
            in1 => \N__42340\,
            in2 => \N__42238\,
            in3 => \N__46878\,
            lcout => \c0.n12_adj_2285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_647_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__42204\,
            in1 => \N__46820\,
            in2 => \_gnd_net_\,
            in3 => \N__46192\,
            lcout => \c0.n17028\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__3__2225_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__42172\,
            in1 => \N__42710\,
            in2 => \N__46133\,
            in3 => \N__46479\,
            lcout => \c0.data_out_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15290_2_lut_LC_16_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52086\,
            in2 => \_gnd_net_\,
            in3 => \N__42171\,
            lcout => \c0.n17593\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__4__2216_LC_16_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__45935\,
            in1 => \N__42910\,
            in2 => \N__42163\,
            in3 => \N__45454\,
            lcout => data_out_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15261_2_lut_LC_16_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__52087\,
            in1 => \N__42465\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n17546_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15557_LC_16_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__42118\,
            in1 => \N__52461\,
            in2 => \N__42112\,
            in3 => \N__52302\,
            lcout => OPEN,
            ltout => \c0.n18017_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18017_bdd_4_lut_LC_16_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52462\,
            in1 => \N__42109\,
            in2 => \N__43171\,
            in3 => \N__43168\,
            lcout => OPEN,
            ltout => \c0.n18020_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_adj_426_LC_16_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__43162\,
            in1 => \N__52463\,
            in2 => \N__43156\,
            in3 => \N__43152\,
            lcout => \c0.n10_adj_2155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__1__2171_LC_16_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43030\,
            in1 => \N__43021\,
            in2 => \_gnd_net_\,
            in3 => \N__42981\,
            lcout => \c0.data_out_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50597\,
            ce => \N__46621\,
            sr => \_gnd_net_\
        );

    \c0.i15289_2_lut_LC_16_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42909\,
            in2 => \_gnd_net_\,
            in3 => \N__52083\,
            lcout => \c0.n17591\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__0__2196_LC_16_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__42883\,
            in1 => \N__52498\,
            in2 => \N__46132\,
            in3 => \N__42851\,
            lcout => data_out_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15211_3_lut_LC_16_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__42709\,
            in1 => \N__42468\,
            in2 => \_gnd_net_\,
            in3 => \N__42401\,
            lcout => \c0.n17522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_547_LC_16_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52497\,
            in2 => \_gnd_net_\,
            in3 => \N__46690\,
            lcout => \c0.n9783\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15423_4_lut_LC_16_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45875\,
            in2 => \_gnd_net_\,
            in3 => \N__45456\,
            lcout => n10055,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15587_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__42326\,
            in1 => \N__48104\,
            in2 => \N__48636\,
            in3 => \N__44231\,
            lcout => \c0.n18047\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15368_2_lut_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43525\,
            in2 => \_gnd_net_\,
            in3 => \N__48097\,
            lcout => \c0.n17495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_594_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__43300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49273\,
            lcout => \c0.n9671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18047_bdd_4_lut_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__43473\,
            in1 => \N__48595\,
            in2 => \N__43305\,
            in3 => \N__43417\,
            lcout => \c0.n18050\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_502_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43410\,
            in1 => \N__43915\,
            in2 => \N__43387\,
            in3 => \N__43335\,
            lcout => \c0.n27_adj_2277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i71_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43304\,
            in1 => \N__49918\,
            in2 => \_gnd_net_\,
            in3 => \N__51207\,
            lcout => data_out_frame2_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44355\,
            in1 => \N__43277\,
            in2 => \_gnd_net_\,
            in3 => \N__48221\,
            lcout => \c0.n5_adj_2321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15611_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__43237\,
            in1 => \N__51620\,
            in2 => \N__43597\,
            in3 => \N__47708\,
            lcout => \c0.n18083\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_548_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43227\,
            in1 => \N__43215\,
            in2 => \N__45601\,
            in3 => \N__43204\,
            lcout => \c0.n16960\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_492_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48865\,
            in1 => \N__44039\,
            in2 => \N__43958\,
            in3 => \N__45597\,
            lcout => \c0.n24_adj_2272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_463_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43907\,
            in1 => \N__43849\,
            in2 => \N__47248\,
            in3 => \N__43804\,
            lcout => \c0.n20_adj_2205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18071_bdd_4_lut_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__48594\,
            in1 => \N__43783\,
            in2 => \N__44283\,
            in3 => \N__44886\,
            lcout => OPEN,
            ltout => \c0.n18074_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15626_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__43696\,
            in1 => \N__51619\,
            in2 => \N__43774\,
            in3 => \N__47709\,
            lcout => \c0.n18089\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15597_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__49194\,
            in1 => \N__44196\,
            in2 => \N__48637\,
            in3 => \N__48215\,
            lcout => OPEN,
            ltout => \c0.n18065_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18065_bdd_4_lut_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__43767\,
            in1 => \N__43732\,
            in2 => \N__43699\,
            in3 => \N__48593\,
            lcout => \c0.n18068\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15577_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__44393\,
            in1 => \N__43686\,
            in2 => \N__48649\,
            in3 => \N__48214\,
            lcout => OPEN,
            ltout => \c0.n18005_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18005_bdd_4_lut_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__49659\,
            in1 => \N__43626\,
            in2 => \N__43600\,
            in3 => \N__48623\,
            lcout => \c0.n18008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14909_3_lut_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49684\,
            in1 => \N__48213\,
            in2 => \_gnd_net_\,
            in3 => \N__43574\,
            lcout => \c0.n17347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i132_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49813\,
            in1 => \N__48993\,
            in2 => \_gnd_net_\,
            in3 => \N__51205\,
            lcout => data_out_frame2_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i51_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51204\,
            in1 => \N__44488\,
            in2 => \_gnd_net_\,
            in3 => \N__44421\,
            lcout => data_out_frame2_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_687_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44394\,
            in1 => \N__44347\,
            in2 => \_gnd_net_\,
            in3 => \N__43947\,
            lcout => \c0.n17127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i72_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__51338\,
            in1 => \N__44272\,
            in2 => \_gnd_net_\,
            in3 => \N__51206\,
            lcout => data_out_frame2_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i95_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__51128\,
            in1 => \_gnd_net_\,
            in2 => \N__49111\,
            in3 => \N__44230\,
            lcout => data_out_frame2_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i120_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44090\,
            in1 => \N__51129\,
            in2 => \_gnd_net_\,
            in3 => \N__44195\,
            lcout => data_out_frame2_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i141_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51126\,
            in1 => \N__44172\,
            in2 => \_gnd_net_\,
            in3 => \N__44106\,
            lcout => data_out_frame2_17_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i56_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44091\,
            in1 => \N__51131\,
            in2 => \_gnd_net_\,
            in3 => \N__44038\,
            lcout => data_out_frame2_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i48_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51127\,
            in1 => \N__44014\,
            in2 => \_gnd_net_\,
            in3 => \N__43948\,
            lcout => data_out_frame2_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i128_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44950\,
            in1 => \N__51130\,
            in2 => \_gnd_net_\,
            in3 => \N__49187\,
            lcout => data_out_frame2_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_613_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44882\,
            in2 => \_gnd_net_\,
            in3 => \N__44853\,
            lcout => \c0.n16926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i41_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51243\,
            in1 => \N__44788\,
            in2 => \_gnd_net_\,
            in3 => \N__44716\,
            lcout => data_out_frame2_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i106_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44695\,
            in1 => \N__49596\,
            in2 => \_gnd_net_\,
            in3 => \N__51245\,
            lcout => data_out_frame2_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45617\,
            in1 => \N__48228\,
            in2 => \_gnd_net_\,
            in3 => \N__44647\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__48229\,
            in1 => \N__44606\,
            in2 => \N__44584\,
            in3 => \N__48650\,
            lcout => \c0.n6_adj_2280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i62_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51244\,
            in1 => \_gnd_net_\,
            in2 => \N__45624\,
            in3 => \N__44569\,
            lcout => data_out_frame2_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18089_bdd_4_lut_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__44518\,
            in1 => \N__44509\,
            in2 => \N__44500\,
            in3 => \N__51621\,
            lcout => \c0.n18092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_510_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45616\,
            in2 => \_gnd_net_\,
            in3 => \N__47198\,
            lcout => \c0.n9678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i7_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__45577\,
            in1 => \N__51622\,
            in2 => \N__51775\,
            in3 => \N__45571\,
            lcout => \c0.tx2.r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50581\,
            ce => \N__51446\,
            sr => \_gnd_net_\
        );

    \c0.data_out_0__0__2244_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__45986\,
            in1 => \N__45516\,
            in2 => \N__45382\,
            in3 => \N__46491\,
            lcout => data_out_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i100_LC_17_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49809\,
            in1 => \N__45336\,
            in2 => \_gnd_net_\,
            in3 => \N__51209\,
            lcout => data_out_frame2_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i110_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51208\,
            in1 => \N__45300\,
            in2 => \_gnd_net_\,
            in3 => \N__45238\,
            lcout => data_out_frame2_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__3__2169_LC_17_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__45213\,
            in1 => \N__45151\,
            in2 => \N__45133\,
            in3 => \N__45118\,
            lcout => \c0.data_out_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50593\,
            ce => \N__46623\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_543_LC_17_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45020\,
            in2 => \_gnd_net_\,
            in3 => \N__45079\,
            lcout => \c0.n17076\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__6__2166_LC_17_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__45034\,
            in1 => \N__45021\,
            in2 => \_gnd_net_\,
            in3 => \N__45004\,
            lcout => \c0.data_out_9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50593\,
            ce => \N__46623\,
            sr => \_gnd_net_\
        );

    \c0.data_out_9__4__2168_LC_17_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__44977\,
            in1 => \N__47029\,
            in2 => \N__47152\,
            in3 => \N__52549\,
            lcout => \c0.data_out_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50598\,
            ce => \N__46624\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_506_LC_17_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47097\,
            in2 => \_gnd_net_\,
            in3 => \N__47056\,
            lcout => \c0.n17058\,
            ltout => \c0.n17058_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_511_LC_17_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47022\,
            in1 => \N__46926\,
            in2 => \N__47011\,
            in3 => \N__47008\,
            lcout => OPEN,
            ltout => \c0.n21_adj_2284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__7__2165_LC_17_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__46993\,
            in1 => \_gnd_net_\,
            in2 => \N__46984\,
            in3 => \N__46981\,
            lcout => \c0.data_out_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50598\,
            ce => \N__46624\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__3__2161_LC_17_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46927\,
            in1 => \N__46912\,
            in2 => \N__46882\,
            in3 => \N__46867\,
            lcout => \c0.data_out_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50598\,
            ce => \N__46624\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__6__2158_LC_17_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46799\,
            in1 => \N__46755\,
            in2 => \N__46726\,
            in3 => \N__46701\,
            lcout => \c0.data_out_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50601\,
            ce => \N__46622\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__5__2191_LC_17_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__46519\,
            in1 => \N__45879\,
            in2 => \N__46501\,
            in3 => \N__46423\,
            lcout => \c0.data_out_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50602\,
            ce => \N__46106\,
            sr => \_gnd_net_\
        );

    \c0.i15206_2_lut_LC_17_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__46024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45947\,
            lcout => \c0.n17450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17999_bdd_4_lut_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__49847\,
            in1 => \N__47830\,
            in2 => \N__49042\,
            in3 => \N__48461\,
            lcout => \c0.n18002\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__47814\,
            in1 => \N__47740\,
            in2 => \N__47734\,
            in3 => \N__47707\,
            lcout => \c0.n22_adj_2353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i6_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__47422\,
            in1 => \N__51651\,
            in2 => \N__51774\,
            in3 => \N__47536\,
            lcout => \c0.tx2.r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50536\,
            ce => \N__51462\,
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_599_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47518\,
            in1 => \N__47509\,
            in2 => \N__47488\,
            in3 => \N__47458\,
            lcout => \c0.n26_adj_2314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__48166\,
            in1 => \N__48876\,
            in2 => \N__47440\,
            in3 => \N__48604\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18083_bdd_4_lut_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__47839\,
            in1 => \N__47431\,
            in2 => \N__47425\,
            in3 => \N__51647\,
            lcout => \c0.n18086\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_614_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47416\,
            in2 => \_gnd_net_\,
            in3 => \N__47377\,
            lcout => OPEN,
            ltout => \c0.n9895_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47301\,
            in1 => \N__47247\,
            in2 => \N__47203\,
            in3 => \N__47199\,
            lcout => OPEN,
            ltout => \c0.n23_adj_2318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i156_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__49144\,
            in1 => \N__49138\,
            in2 => \N__49126\,
            in3 => \N__49123\,
            lcout => \c0.data_out_frame2_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50556\,
            ce => \N__51216\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i143_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49110\,
            in1 => \N__49038\,
            in2 => \_gnd_net_\,
            in3 => \N__51217\,
            lcout => data_out_frame2_17_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15500_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__49755\,
            in1 => \N__48638\,
            in2 => \N__48222\,
            in3 => \N__49024\,
            lcout => OPEN,
            ltout => \c0.n17945_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n17945_bdd_4_lut_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48639\,
            in1 => \N__48780\,
            in2 => \N__49018\,
            in3 => \N__48989\,
            lcout => \c0.n17948\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i47_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48940\,
            in1 => \N__48872\,
            in2 => \_gnd_net_\,
            in3 => \N__51218\,
            lcout => data_out_frame2_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i140_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51219\,
            in1 => \N__48840\,
            in2 => \_gnd_net_\,
            in3 => \N__48781\,
            lcout => data_out_frame2_17_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50576\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i89_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48767\,
            in1 => \N__49686\,
            in2 => \_gnd_net_\,
            in3 => \N__51222\,
            lcout => data_out_frame2_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50576\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15313_3_lut_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__48701\,
            in1 => \N__48640\,
            in2 => \_gnd_net_\,
            in3 => \N__48212\,
            lcout => \c0.n17563\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i135_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49916\,
            in1 => \N__49843\,
            in2 => \_gnd_net_\,
            in3 => \N__51220\,
            lcout => data_out_frame2_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50576\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i148_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49801\,
            in1 => \N__49756\,
            in2 => \_gnd_net_\,
            in3 => \N__51221\,
            lcout => data_out_frame2_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50576\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_563_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49742\,
            in1 => \N__49685\,
            in2 => \_gnd_net_\,
            in3 => \N__49663\,
            lcout => \c0.n16923\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_578_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50635\,
            in1 => \N__49595\,
            in2 => \_gnd_net_\,
            in3 => \N__49182\,
            lcout => \c0.n9910\,
            ltout => \c0.n9910_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_622_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49564\,
            in1 => \N__49540\,
            in2 => \N__49507\,
            in3 => \N__49504\,
            lcout => \c0.n16_adj_2327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_623_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49477\,
            in1 => \N__49432\,
            in2 => \N__49384\,
            in3 => \N__49344\,
            lcout => OPEN,
            ltout => \c0.n17_adj_2328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i154_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49300\,
            in1 => \N__49294\,
            in2 => \N__49237\,
            in3 => \N__49234\,
            lcout => \c0.data_out_frame2_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50582\,
            ce => \N__51215\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_619_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__49183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50636\,
            lcout => \c0.n16940\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_18_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52548\,
            in1 => \N__52512\,
            in2 => \_gnd_net_\,
            in3 => \N__52099\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__51781\,
            in1 => \N__52404\,
            in2 => \N__52306\,
            in3 => \N__52265\,
            lcout => \c0.n18095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15367_2_lut_LC_18_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52141\,
            in2 => \_gnd_net_\,
            in3 => \N__52038\,
            lcout => \c0.n17632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i4_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__51770\,
            in1 => \N__51670\,
            in2 => \N__51655\,
            in3 => \N__51496\,
            lcout => \c0.tx2.r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50583\,
            ce => \N__51463\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i136_LC_19_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__51346\,
            in1 => \N__50634\,
            in2 => \_gnd_net_\,
            in3 => \N__51272\,
            lcout => data_out_frame2_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50594\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
