// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Aug 25 2019 21:15:49

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    output PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    input PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    output PIN_1;
    output LED;
    input CLK;

    wire N__20080;
    wire N__20079;
    wire N__20078;
    wire N__20069;
    wire N__20068;
    wire N__20067;
    wire N__20060;
    wire N__20059;
    wire N__20058;
    wire N__20051;
    wire N__20050;
    wire N__20049;
    wire N__20042;
    wire N__20041;
    wire N__20040;
    wire N__20033;
    wire N__20032;
    wire N__20031;
    wire N__20014;
    wire N__20013;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19983;
    wire N__19978;
    wire N__19977;
    wire N__19974;
    wire N__19973;
    wire N__19970;
    wire N__19969;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19952;
    wire N__19947;
    wire N__19946;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19922;
    wire N__19915;
    wire N__19914;
    wire N__19913;
    wire N__19912;
    wire N__19909;
    wire N__19904;
    wire N__19903;
    wire N__19900;
    wire N__19899;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19883;
    wire N__19876;
    wire N__19875;
    wire N__19872;
    wire N__19871;
    wire N__19870;
    wire N__19867;
    wire N__19862;
    wire N__19861;
    wire N__19860;
    wire N__19859;
    wire N__19858;
    wire N__19857;
    wire N__19856;
    wire N__19853;
    wire N__19848;
    wire N__19841;
    wire N__19834;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19818;
    wire N__19817;
    wire N__19816;
    wire N__19815;
    wire N__19812;
    wire N__19811;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19780;
    wire N__19779;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19764;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19747;
    wire N__19746;
    wire N__19745;
    wire N__19742;
    wire N__19741;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19723;
    wire N__19722;
    wire N__19721;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19677;
    wire N__19676;
    wire N__19675;
    wire N__19674;
    wire N__19673;
    wire N__19672;
    wire N__19671;
    wire N__19670;
    wire N__19669;
    wire N__19668;
    wire N__19667;
    wire N__19666;
    wire N__19665;
    wire N__19664;
    wire N__19663;
    wire N__19662;
    wire N__19661;
    wire N__19660;
    wire N__19659;
    wire N__19658;
    wire N__19657;
    wire N__19656;
    wire N__19655;
    wire N__19654;
    wire N__19653;
    wire N__19652;
    wire N__19651;
    wire N__19650;
    wire N__19649;
    wire N__19648;
    wire N__19647;
    wire N__19646;
    wire N__19645;
    wire N__19644;
    wire N__19643;
    wire N__19642;
    wire N__19641;
    wire N__19640;
    wire N__19639;
    wire N__19638;
    wire N__19637;
    wire N__19636;
    wire N__19635;
    wire N__19634;
    wire N__19633;
    wire N__19632;
    wire N__19631;
    wire N__19630;
    wire N__19629;
    wire N__19628;
    wire N__19627;
    wire N__19626;
    wire N__19625;
    wire N__19624;
    wire N__19623;
    wire N__19622;
    wire N__19621;
    wire N__19620;
    wire N__19619;
    wire N__19618;
    wire N__19617;
    wire N__19616;
    wire N__19615;
    wire N__19614;
    wire N__19613;
    wire N__19612;
    wire N__19611;
    wire N__19610;
    wire N__19609;
    wire N__19608;
    wire N__19607;
    wire N__19606;
    wire N__19605;
    wire N__19604;
    wire N__19603;
    wire N__19602;
    wire N__19601;
    wire N__19600;
    wire N__19599;
    wire N__19598;
    wire N__19597;
    wire N__19596;
    wire N__19595;
    wire N__19594;
    wire N__19593;
    wire N__19592;
    wire N__19591;
    wire N__19590;
    wire N__19589;
    wire N__19588;
    wire N__19587;
    wire N__19586;
    wire N__19585;
    wire N__19584;
    wire N__19583;
    wire N__19582;
    wire N__19581;
    wire N__19580;
    wire N__19579;
    wire N__19578;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19354;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19342;
    wire N__19341;
    wire N__19340;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19300;
    wire N__19291;
    wire N__19288;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19248;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19240;
    wire N__19237;
    wire N__19232;
    wire N__19225;
    wire N__19222;
    wire N__19221;
    wire N__19220;
    wire N__19219;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19205;
    wire N__19198;
    wire N__19195;
    wire N__19194;
    wire N__19193;
    wire N__19192;
    wire N__19191;
    wire N__19186;
    wire N__19183;
    wire N__19178;
    wire N__19171;
    wire N__19168;
    wire N__19167;
    wire N__19166;
    wire N__19165;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19151;
    wire N__19144;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19138;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19127;
    wire N__19122;
    wire N__19115;
    wire N__19108;
    wire N__19107;
    wire N__19106;
    wire N__19105;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19078;
    wire N__19077;
    wire N__19074;
    wire N__19071;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19056;
    wire N__19051;
    wire N__19048;
    wire N__19047;
    wire N__19046;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19024;
    wire N__19021;
    wire N__19020;
    wire N__19019;
    wire N__19014;
    wire N__19011;
    wire N__19006;
    wire N__19003;
    wire N__19002;
    wire N__19001;
    wire N__18996;
    wire N__18993;
    wire N__18988;
    wire N__18987;
    wire N__18984;
    wire N__18983;
    wire N__18978;
    wire N__18975;
    wire N__18970;
    wire N__18969;
    wire N__18968;
    wire N__18963;
    wire N__18960;
    wire N__18955;
    wire N__18954;
    wire N__18949;
    wire N__18948;
    wire N__18947;
    wire N__18944;
    wire N__18939;
    wire N__18934;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18869;
    wire N__18864;
    wire N__18861;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18849;
    wire N__18848;
    wire N__18847;
    wire N__18844;
    wire N__18839;
    wire N__18836;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18819;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18804;
    wire N__18799;
    wire N__18798;
    wire N__18797;
    wire N__18796;
    wire N__18795;
    wire N__18792;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18784;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18768;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18762;
    wire N__18759;
    wire N__18754;
    wire N__18749;
    wire N__18746;
    wire N__18741;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18720;
    wire N__18719;
    wire N__18718;
    wire N__18717;
    wire N__18716;
    wire N__18715;
    wire N__18714;
    wire N__18713;
    wire N__18712;
    wire N__18711;
    wire N__18710;
    wire N__18709;
    wire N__18708;
    wire N__18705;
    wire N__18700;
    wire N__18697;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18674;
    wire N__18671;
    wire N__18666;
    wire N__18663;
    wire N__18658;
    wire N__18657;
    wire N__18656;
    wire N__18655;
    wire N__18654;
    wire N__18649;
    wire N__18646;
    wire N__18641;
    wire N__18636;
    wire N__18633;
    wire N__18626;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18594;
    wire N__18593;
    wire N__18592;
    wire N__18591;
    wire N__18590;
    wire N__18589;
    wire N__18588;
    wire N__18587;
    wire N__18586;
    wire N__18583;
    wire N__18582;
    wire N__18579;
    wire N__18578;
    wire N__18577;
    wire N__18576;
    wire N__18573;
    wire N__18572;
    wire N__18571;
    wire N__18570;
    wire N__18569;
    wire N__18568;
    wire N__18567;
    wire N__18566;
    wire N__18565;
    wire N__18562;
    wire N__18555;
    wire N__18550;
    wire N__18543;
    wire N__18536;
    wire N__18533;
    wire N__18532;
    wire N__18531;
    wire N__18528;
    wire N__18527;
    wire N__18526;
    wire N__18521;
    wire N__18520;
    wire N__18519;
    wire N__18518;
    wire N__18515;
    wire N__18514;
    wire N__18513;
    wire N__18510;
    wire N__18501;
    wire N__18496;
    wire N__18493;
    wire N__18490;
    wire N__18485;
    wire N__18484;
    wire N__18483;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18468;
    wire N__18465;
    wire N__18458;
    wire N__18453;
    wire N__18450;
    wire N__18443;
    wire N__18436;
    wire N__18429;
    wire N__18406;
    wire N__18403;
    wire N__18402;
    wire N__18401;
    wire N__18400;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18385;
    wire N__18376;
    wire N__18375;
    wire N__18374;
    wire N__18373;
    wire N__18372;
    wire N__18371;
    wire N__18370;
    wire N__18369;
    wire N__18366;
    wire N__18365;
    wire N__18362;
    wire N__18361;
    wire N__18358;
    wire N__18357;
    wire N__18356;
    wire N__18355;
    wire N__18354;
    wire N__18353;
    wire N__18352;
    wire N__18349;
    wire N__18348;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18334;
    wire N__18333;
    wire N__18332;
    wire N__18331;
    wire N__18330;
    wire N__18329;
    wire N__18324;
    wire N__18319;
    wire N__18312;
    wire N__18309;
    wire N__18306;
    wire N__18305;
    wire N__18304;
    wire N__18303;
    wire N__18302;
    wire N__18301;
    wire N__18298;
    wire N__18293;
    wire N__18286;
    wire N__18283;
    wire N__18282;
    wire N__18279;
    wire N__18278;
    wire N__18275;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18253;
    wire N__18248;
    wire N__18237;
    wire N__18232;
    wire N__18229;
    wire N__18224;
    wire N__18215;
    wire N__18208;
    wire N__18199;
    wire N__18194;
    wire N__18181;
    wire N__18178;
    wire N__18175;
    wire N__18174;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18096;
    wire N__18095;
    wire N__18094;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18082;
    wire N__18073;
    wire N__18070;
    wire N__18067;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18036;
    wire N__18035;
    wire N__18034;
    wire N__18031;
    wire N__18026;
    wire N__18023;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17993;
    wire N__17988;
    wire N__17985;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17968;
    wire N__17965;
    wire N__17964;
    wire N__17961;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17922;
    wire N__17919;
    wire N__17916;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17904;
    wire N__17901;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17863;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17851;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17839;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17827;
    wire N__17824;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17791;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17781;
    wire N__17776;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17761;
    wire N__17758;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17746;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17727;
    wire N__17726;
    wire N__17725;
    wire N__17724;
    wire N__17723;
    wire N__17722;
    wire N__17721;
    wire N__17720;
    wire N__17719;
    wire N__17718;
    wire N__17717;
    wire N__17716;
    wire N__17715;
    wire N__17712;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17649;
    wire N__17648;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17620;
    wire N__17619;
    wire N__17618;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17583;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17485;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17465;
    wire N__17460;
    wire N__17457;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17391;
    wire N__17388;
    wire N__17385;
    wire N__17382;
    wire N__17379;
    wire N__17374;
    wire N__17371;
    wire N__17370;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17346;
    wire N__17341;
    wire N__17338;
    wire N__17337;
    wire N__17334;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17316;
    wire N__17311;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17292;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17275;
    wire N__17272;
    wire N__17271;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17251;
    wire N__17248;
    wire N__17247;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17217;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17187;
    wire N__17186;
    wire N__17185;
    wire N__17184;
    wire N__17183;
    wire N__17182;
    wire N__17181;
    wire N__17180;
    wire N__17179;
    wire N__17178;
    wire N__17177;
    wire N__17176;
    wire N__17175;
    wire N__17174;
    wire N__17173;
    wire N__17172;
    wire N__17171;
    wire N__17170;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17115;
    wire N__17114;
    wire N__17113;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17105;
    wire N__17104;
    wire N__17103;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17093;
    wire N__17092;
    wire N__17091;
    wire N__17090;
    wire N__17089;
    wire N__17088;
    wire N__17087;
    wire N__17086;
    wire N__17085;
    wire N__17076;
    wire N__17075;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17061;
    wire N__17060;
    wire N__17057;
    wire N__17056;
    wire N__17053;
    wire N__17040;
    wire N__17037;
    wire N__17032;
    wire N__17029;
    wire N__17024;
    wire N__17021;
    wire N__17020;
    wire N__17019;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17011;
    wire N__17010;
    wire N__17009;
    wire N__17008;
    wire N__17007;
    wire N__17006;
    wire N__17001;
    wire N__16996;
    wire N__16991;
    wire N__16988;
    wire N__16981;
    wire N__16976;
    wire N__16967;
    wire N__16962;
    wire N__16961;
    wire N__16960;
    wire N__16959;
    wire N__16958;
    wire N__16957;
    wire N__16956;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16942;
    wire N__16935;
    wire N__16920;
    wire N__16909;
    wire N__16906;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16882;
    wire N__16881;
    wire N__16880;
    wire N__16879;
    wire N__16878;
    wire N__16877;
    wire N__16876;
    wire N__16875;
    wire N__16874;
    wire N__16873;
    wire N__16872;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16839;
    wire N__16838;
    wire N__16837;
    wire N__16836;
    wire N__16835;
    wire N__16834;
    wire N__16833;
    wire N__16832;
    wire N__16831;
    wire N__16830;
    wire N__16829;
    wire N__16828;
    wire N__16827;
    wire N__16826;
    wire N__16825;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16791;
    wire N__16738;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16674;
    wire N__16671;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16656;
    wire N__16651;
    wire N__16648;
    wire N__16647;
    wire N__16646;
    wire N__16643;
    wire N__16638;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16594;
    wire N__16591;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16545;
    wire N__16544;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16516;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16505;
    wire N__16502;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16464;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16437;
    wire N__16436;
    wire N__16435;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16405;
    wire N__16404;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16371;
    wire N__16368;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16336;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16328;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16306;
    wire N__16303;
    wire N__16302;
    wire N__16301;
    wire N__16298;
    wire N__16295;
    wire N__16292;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16272;
    wire N__16269;
    wire N__16268;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16246;
    wire N__16245;
    wire N__16244;
    wire N__16243;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16229;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16184;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16171;
    wire N__16162;
    wire N__16161;
    wire N__16158;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16102;
    wire N__16099;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16069;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16051;
    wire N__16050;
    wire N__16047;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16015;
    wire N__16012;
    wire N__16011;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15985;
    wire N__15982;
    wire N__15981;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15966;
    wire N__15963;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15933;
    wire N__15930;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15918;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15906;
    wire N__15905;
    wire N__15902;
    wire N__15897;
    wire N__15892;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15870;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15853;
    wire N__15850;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15826;
    wire N__15823;
    wire N__15820;
    wire N__15819;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15772;
    wire N__15769;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15750;
    wire N__15747;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15717;
    wire N__15714;
    wire N__15711;
    wire N__15706;
    wire N__15705;
    wire N__15704;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15657;
    wire N__15656;
    wire N__15653;
    wire N__15652;
    wire N__15651;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15633;
    wire N__15632;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15611;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15596;
    wire N__15593;
    wire N__15586;
    wire N__15583;
    wire N__15568;
    wire N__15567;
    wire N__15566;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15558;
    wire N__15557;
    wire N__15556;
    wire N__15555;
    wire N__15550;
    wire N__15541;
    wire N__15540;
    wire N__15539;
    wire N__15538;
    wire N__15537;
    wire N__15536;
    wire N__15535;
    wire N__15534;
    wire N__15533;
    wire N__15532;
    wire N__15531;
    wire N__15530;
    wire N__15529;
    wire N__15528;
    wire N__15523;
    wire N__15518;
    wire N__15517;
    wire N__15516;
    wire N__15515;
    wire N__15512;
    wire N__15511;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15503;
    wire N__15502;
    wire N__15501;
    wire N__15500;
    wire N__15489;
    wire N__15482;
    wire N__15479;
    wire N__15478;
    wire N__15475;
    wire N__15474;
    wire N__15473;
    wire N__15472;
    wire N__15471;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15451;
    wire N__15438;
    wire N__15435;
    wire N__15430;
    wire N__15429;
    wire N__15426;
    wire N__15421;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15397;
    wire N__15394;
    wire N__15379;
    wire N__15376;
    wire N__15375;
    wire N__15374;
    wire N__15373;
    wire N__15372;
    wire N__15371;
    wire N__15370;
    wire N__15369;
    wire N__15368;
    wire N__15367;
    wire N__15366;
    wire N__15365;
    wire N__15364;
    wire N__15361;
    wire N__15356;
    wire N__15347;
    wire N__15346;
    wire N__15345;
    wire N__15344;
    wire N__15343;
    wire N__15342;
    wire N__15341;
    wire N__15340;
    wire N__15339;
    wire N__15338;
    wire N__15337;
    wire N__15336;
    wire N__15335;
    wire N__15334;
    wire N__15333;
    wire N__15332;
    wire N__15321;
    wire N__15318;
    wire N__15311;
    wire N__15304;
    wire N__15295;
    wire N__15290;
    wire N__15289;
    wire N__15288;
    wire N__15287;
    wire N__15286;
    wire N__15285;
    wire N__15284;
    wire N__15283;
    wire N__15282;
    wire N__15279;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15251;
    wire N__15238;
    wire N__15233;
    wire N__15214;
    wire N__15213;
    wire N__15212;
    wire N__15211;
    wire N__15210;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15199;
    wire N__15198;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15187;
    wire N__15186;
    wire N__15183;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15167;
    wire N__15166;
    wire N__15165;
    wire N__15164;
    wire N__15163;
    wire N__15156;
    wire N__15153;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15120;
    wire N__15111;
    wire N__15110;
    wire N__15107;
    wire N__15102;
    wire N__15099;
    wire N__15096;
    wire N__15093;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15075;
    wire N__15072;
    wire N__15069;
    wire N__15064;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15030;
    wire N__15027;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15001;
    wire N__14998;
    wire N__14997;
    wire N__14994;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14959;
    wire N__14958;
    wire N__14957;
    wire N__14954;
    wire N__14949;
    wire N__14946;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14934;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14907;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14895;
    wire N__14894;
    wire N__14891;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14875;
    wire N__14874;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14830;
    wire N__14829;
    wire N__14826;
    wire N__14823;
    wire N__14820;
    wire N__14819;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14807;
    wire N__14804;
    wire N__14799;
    wire N__14794;
    wire N__14793;
    wire N__14790;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14776;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14760;
    wire N__14749;
    wire N__14748;
    wire N__14747;
    wire N__14744;
    wire N__14743;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14713;
    wire N__14710;
    wire N__14709;
    wire N__14706;
    wire N__14705;
    wire N__14704;
    wire N__14701;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14667;
    wire N__14666;
    wire N__14665;
    wire N__14662;
    wire N__14657;
    wire N__14654;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14629;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14617;
    wire N__14614;
    wire N__14613;
    wire N__14612;
    wire N__14611;
    wire N__14608;
    wire N__14603;
    wire N__14600;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14579;
    wire N__14574;
    wire N__14571;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14502;
    wire N__14499;
    wire N__14498;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14475;
    wire N__14470;
    wire N__14467;
    wire N__14466;
    wire N__14465;
    wire N__14464;
    wire N__14461;
    wire N__14456;
    wire N__14453;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14410;
    wire N__14409;
    wire N__14406;
    wire N__14403;
    wire N__14398;
    wire N__14395;
    wire N__14394;
    wire N__14391;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14379;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14361;
    wire N__14360;
    wire N__14357;
    wire N__14352;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14283;
    wire N__14280;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14251;
    wire N__14248;
    wire N__14247;
    wire N__14246;
    wire N__14245;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14237;
    wire N__14234;
    wire N__14233;
    wire N__14228;
    wire N__14227;
    wire N__14222;
    wire N__14221;
    wire N__14218;
    wire N__14217;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14196;
    wire N__14185;
    wire N__14184;
    wire N__14181;
    wire N__14180;
    wire N__14179;
    wire N__14178;
    wire N__14177;
    wire N__14176;
    wire N__14175;
    wire N__14174;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14153;
    wire N__14150;
    wire N__14145;
    wire N__14140;
    wire N__14125;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14117;
    wire N__14116;
    wire N__14113;
    wire N__14112;
    wire N__14111;
    wire N__14110;
    wire N__14109;
    wire N__14106;
    wire N__14105;
    wire N__14104;
    wire N__14103;
    wire N__14100;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14073;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13965;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13935;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13903;
    wire N__13902;
    wire N__13901;
    wire N__13900;
    wire N__13897;
    wire N__13890;
    wire N__13885;
    wire N__13884;
    wire N__13883;
    wire N__13878;
    wire N__13875;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13834;
    wire N__13833;
    wire N__13830;
    wire N__13827;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13797;
    wire N__13794;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13777;
    wire N__13774;
    wire N__13773;
    wire N__13770;
    wire N__13767;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13750;
    wire N__13749;
    wire N__13748;
    wire N__13745;
    wire N__13740;
    wire N__13737;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13709;
    wire N__13704;
    wire N__13701;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13689;
    wire N__13688;
    wire N__13685;
    wire N__13680;
    wire N__13675;
    wire N__13672;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13642;
    wire N__13641;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13621;
    wire N__13618;
    wire N__13617;
    wire N__13614;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13594;
    wire N__13591;
    wire N__13588;
    wire N__13585;
    wire N__13584;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13558;
    wire N__13555;
    wire N__13552;
    wire N__13549;
    wire N__13548;
    wire N__13545;
    wire N__13542;
    wire N__13541;
    wire N__13536;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13507;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13494;
    wire N__13489;
    wire N__13486;
    wire N__13485;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13467;
    wire N__13464;
    wire N__13459;
    wire N__13456;
    wire N__13453;
    wire N__13452;
    wire N__13449;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13441;
    wire N__13438;
    wire N__13433;
    wire N__13428;
    wire N__13423;
    wire N__13420;
    wire N__13417;
    wire N__13414;
    wire N__13411;
    wire N__13408;
    wire N__13405;
    wire N__13404;
    wire N__13401;
    wire N__13400;
    wire N__13399;
    wire N__13396;
    wire N__13395;
    wire N__13392;
    wire N__13389;
    wire N__13386;
    wire N__13383;
    wire N__13380;
    wire N__13375;
    wire N__13366;
    wire N__13365;
    wire N__13362;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13347;
    wire N__13344;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13329;
    wire N__13328;
    wire N__13327;
    wire N__13324;
    wire N__13321;
    wire N__13316;
    wire N__13313;
    wire N__13308;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13282;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13270;
    wire N__13267;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13255;
    wire N__13252;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13219;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13192;
    wire N__13189;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13140;
    wire N__13137;
    wire N__13136;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13108;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13054;
    wire N__13051;
    wire N__13050;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13039;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13021;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13013;
    wire N__13010;
    wire N__13009;
    wire N__13006;
    wire N__13003;
    wire N__13000;
    wire N__12997;
    wire N__12988;
    wire N__12985;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12942;
    wire N__12941;
    wire N__12938;
    wire N__12935;
    wire N__12934;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12921;
    wire N__12916;
    wire N__12913;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12886;
    wire N__12883;
    wire N__12880;
    wire N__12879;
    wire N__12878;
    wire N__12875;
    wire N__12870;
    wire N__12865;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12844;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12829;
    wire N__12828;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12811;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12775;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12767;
    wire N__12764;
    wire N__12759;
    wire N__12754;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12739;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12727;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12675;
    wire N__12674;
    wire N__12671;
    wire N__12666;
    wire N__12661;
    wire N__12658;
    wire N__12657;
    wire N__12656;
    wire N__12653;
    wire N__12648;
    wire N__12643;
    wire N__12642;
    wire N__12641;
    wire N__12638;
    wire N__12637;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12618;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12606;
    wire N__12603;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12538;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12508;
    wire N__12505;
    wire N__12504;
    wire N__12501;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12481;
    wire N__12480;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12472;
    wire N__12469;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12455;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12387;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12366;
    wire N__12361;
    wire N__12358;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12324;
    wire N__12323;
    wire N__12320;
    wire N__12315;
    wire N__12310;
    wire N__12307;
    wire N__12306;
    wire N__12305;
    wire N__12302;
    wire N__12297;
    wire N__12292;
    wire N__12289;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12259;
    wire N__12258;
    wire N__12255;
    wire N__12252;
    wire N__12251;
    wire N__12246;
    wire N__12243;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12199;
    wire N__12198;
    wire N__12195;
    wire N__12194;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12139;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12121;
    wire N__12120;
    wire N__12115;
    wire N__12114;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12091;
    wire N__12090;
    wire N__12087;
    wire N__12086;
    wire N__12083;
    wire N__12082;
    wire N__12079;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12049;
    wire N__12046;
    wire N__12043;
    wire N__12040;
    wire N__12037;
    wire N__12036;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12019;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__11998;
    wire N__11997;
    wire N__11996;
    wire N__11993;
    wire N__11992;
    wire N__11989;
    wire N__11986;
    wire N__11983;
    wire N__11980;
    wire N__11977;
    wire N__11974;
    wire N__11969;
    wire N__11964;
    wire N__11959;
    wire N__11956;
    wire N__11955;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11940;
    wire N__11935;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11866;
    wire N__11863;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11835;
    wire N__11832;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11824;
    wire N__11821;
    wire N__11816;
    wire N__11813;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11796;
    wire N__11791;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11779;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11762;
    wire N__11757;
    wire N__11754;
    wire N__11749;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11741;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11718;
    wire N__11713;
    wire N__11712;
    wire N__11711;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11690;
    wire N__11687;
    wire N__11684;
    wire N__11681;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11667;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11638;
    wire N__11635;
    wire N__11630;
    wire N__11627;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11518;
    wire N__11517;
    wire N__11514;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11385;
    wire N__11382;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11337;
    wire N__11336;
    wire N__11333;
    wire N__11328;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11303;
    wire N__11298;
    wire N__11295;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11278;
    wire N__11273;
    wire N__11268;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11230;
    wire N__11227;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11196;
    wire N__11195;
    wire N__11192;
    wire N__11187;
    wire N__11182;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11170;
    wire N__11167;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11131;
    wire N__11128;
    wire N__11127;
    wire N__11124;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11104;
    wire N__11101;
    wire N__11100;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11083;
    wire N__11080;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11049;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11032;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11020;
    wire N__11017;
    wire N__11014;
    wire N__11013;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__10996;
    wire N__10993;
    wire N__10992;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10957;
    wire N__10956;
    wire N__10953;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10933;
    wire N__10932;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10897;
    wire N__10896;
    wire N__10895;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10885;
    wire N__10882;
    wire N__10875;
    wire N__10870;
    wire N__10867;
    wire N__10866;
    wire N__10863;
    wire N__10860;
    wire N__10857;
    wire N__10854;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10803;
    wire N__10802;
    wire N__10799;
    wire N__10794;
    wire N__10789;
    wire N__10788;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10765;
    wire N__10762;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10750;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10678;
    wire N__10675;
    wire N__10674;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10653;
    wire N__10652;
    wire N__10651;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10642;
    wire N__10635;
    wire N__10628;
    wire N__10623;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10606;
    wire N__10605;
    wire N__10604;
    wire N__10603;
    wire N__10602;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10584;
    wire N__10579;
    wire N__10570;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10566;
    wire N__10563;
    wire N__10556;
    wire N__10553;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10539;
    wire N__10538;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10530;
    wire N__10529;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10513;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10499;
    wire N__10498;
    wire N__10495;
    wire N__10494;
    wire N__10487;
    wire N__10486;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10446;
    wire N__10441;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10402;
    wire N__10399;
    wire N__10398;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10368;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10360;
    wire N__10357;
    wire N__10356;
    wire N__10347;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10327;
    wire N__10324;
    wire N__10323;
    wire N__10320;
    wire N__10319;
    wire N__10318;
    wire N__10317;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10299;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10254;
    wire N__10251;
    wire N__10248;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10207;
    wire N__10204;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10186;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10174;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10162;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10150;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10138;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10126;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10114;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10072;
    wire N__10071;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10027;
    wire N__10024;
    wire N__10023;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10006;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9998;
    wire N__9993;
    wire N__9990;
    wire N__9985;
    wire N__9984;
    wire N__9981;
    wire N__9980;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9965;
    wire N__9958;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9940;
    wire N__9937;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9922;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9903;
    wire N__9902;
    wire N__9901;
    wire N__9898;
    wire N__9891;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9879;
    wire N__9878;
    wire N__9877;
    wire N__9876;
    wire N__9873;
    wire N__9864;
    wire N__9863;
    wire N__9858;
    wire N__9857;
    wire N__9856;
    wire N__9855;
    wire N__9854;
    wire N__9853;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9841;
    wire N__9832;
    wire N__9823;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9819;
    wire N__9818;
    wire N__9817;
    wire N__9816;
    wire N__9815;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9803;
    wire N__9796;
    wire N__9787;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9771;
    wire N__9770;
    wire N__9769;
    wire N__9768;
    wire N__9767;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9748;
    wire N__9741;
    wire N__9736;
    wire N__9735;
    wire N__9734;
    wire N__9729;
    wire N__9726;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9702;
    wire N__9701;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9577;
    wire N__9574;
    wire N__9571;
    wire N__9568;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9485;
    wire N__9480;
    wire N__9477;
    wire N__9472;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9464;
    wire N__9459;
    wire N__9456;
    wire N__9451;
    wire N__9450;
    wire N__9447;
    wire N__9442;
    wire N__9439;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9427;
    wire N__9426;
    wire N__9421;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9339;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9283;
    wire N__9282;
    wire N__9277;
    wire N__9274;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9262;
    wire N__9259;
    wire N__9258;
    wire N__9253;
    wire N__9250;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9231;
    wire N__9226;
    wire N__9223;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9144;
    wire N__9143;
    wire N__9142;
    wire N__9141;
    wire N__9140;
    wire N__9137;
    wire N__9132;
    wire N__9125;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9102;
    wire N__9097;
    wire N__9096;
    wire N__9095;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9091;
    wire N__9088;
    wire N__9081;
    wire N__9074;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9053;
    wire N__9052;
    wire N__9051;
    wire N__9050;
    wire N__9049;
    wire N__9048;
    wire N__9047;
    wire N__9046;
    wire N__9045;
    wire N__9044;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9005;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8976;
    wire N__8971;
    wire N__8970;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8950;
    wire N__8947;
    wire N__8946;
    wire N__8945;
    wire N__8944;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8930;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8898;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8886;
    wire N__8885;
    wire N__8884;
    wire N__8883;
    wire N__8882;
    wire N__8881;
    wire N__8878;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8854;
    wire N__8851;
    wire N__8850;
    wire N__8849;
    wire N__8848;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8834;
    wire N__8833;
    wire N__8832;
    wire N__8831;
    wire N__8830;
    wire N__8829;
    wire N__8826;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8810;
    wire N__8801;
    wire N__8788;
    wire N__8787;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8779;
    wire N__8776;
    wire N__8775;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8754;
    wire N__8751;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8736;
    wire N__8735;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8723;
    wire N__8720;
    wire N__8715;
    wire N__8710;
    wire N__8709;
    wire N__8708;
    wire N__8707;
    wire N__8706;
    wire N__8705;
    wire N__8700;
    wire N__8697;
    wire N__8690;
    wire N__8687;
    wire N__8682;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8669;
    wire N__8662;
    wire N__8657;
    wire N__8650;
    wire N__8649;
    wire N__8648;
    wire N__8647;
    wire N__8646;
    wire N__8645;
    wire N__8644;
    wire N__8641;
    wire N__8636;
    wire N__8635;
    wire N__8634;
    wire N__8633;
    wire N__8632;
    wire N__8627;
    wire N__8626;
    wire N__8625;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8596;
    wire N__8581;
    wire N__8580;
    wire N__8579;
    wire N__8576;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8568;
    wire N__8567;
    wire N__8566;
    wire N__8561;
    wire N__8556;
    wire N__8553;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8526;
    wire N__8525;
    wire N__8524;
    wire N__8521;
    wire N__8520;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8501;
    wire N__8494;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8422;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8410;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8395;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8365;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8353;
    wire N__8352;
    wire N__8351;
    wire N__8348;
    wire N__8343;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8272;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8260;
    wire N__8257;
    wire N__8256;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8239;
    wire N__8236;
    wire N__8235;
    wire N__8234;
    wire N__8233;
    wire N__8232;
    wire N__8231;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8216;
    wire N__8211;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7987;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7966;
    wire N__7963;
    wire N__7960;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7942;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7930;
    wire N__7927;
    wire N__7924;
    wire N__7921;
    wire N__7918;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7882;
    wire N__7879;
    wire VCCG0;
    wire PIN_2_c;
    wire \c0.rx.r_Rx_Data_RZ0 ;
    wire bfn_5_22_0_;
    wire \c0.tx.r_Clock_Count_i_1 ;
    wire \c0.tx.r_Clock_Count12_cry_0 ;
    wire \c0.tx.r_Clock_Count_i_2 ;
    wire \c0.tx.r_Clock_Count12_cry_1 ;
    wire \c0.tx.r_Clock_Count_i_3 ;
    wire \c0.tx.r_Clock_Count12_cry_2 ;
    wire \c0.tx.r_Clock_Count12 ;
    wire \c0.tx.r_Clock_Count_i_0 ;
    wire \c0.rx.r_Rx_Bytece_0_4_cascade_ ;
    wire \c0.rx.N_336_cascade_ ;
    wire \c0.rx.r_Rx_Bytece_0_1 ;
    wire \c0.rx.r_SM_Main_RNI58REZ0Z_0_cascade_ ;
    wire \c0.rx.rx_data_ready ;
    wire blink_counterZ0Z_0;
    wire bfn_6_21_0_;
    wire blink_counterZ0Z_1;
    wire blink_counter_cry_0;
    wire blink_counterZ0Z_2;
    wire blink_counter_cry_1;
    wire blink_counterZ0Z_3;
    wire blink_counter_cry_2;
    wire blink_counterZ0Z_4;
    wire blink_counter_cry_3;
    wire blink_counterZ0Z_5;
    wire blink_counter_cry_4;
    wire blink_counterZ0Z_6;
    wire blink_counter_cry_5;
    wire blink_counterZ0Z_7;
    wire blink_counter_cry_6;
    wire blink_counter_cry_7;
    wire blink_counterZ0Z_8;
    wire bfn_6_22_0_;
    wire blink_counterZ0Z_9;
    wire blink_counter_cry_8;
    wire blink_counterZ0Z_10;
    wire blink_counter_cry_9;
    wire blink_counterZ0Z_11;
    wire blink_counter_cry_10;
    wire blink_counterZ0Z_12;
    wire blink_counter_cry_11;
    wire blink_counterZ0Z_13;
    wire blink_counter_cry_12;
    wire blink_counterZ0Z_14;
    wire blink_counter_cry_13;
    wire blink_counterZ0Z_15;
    wire blink_counter_cry_14;
    wire blink_counter_cry_15;
    wire blink_counterZ0Z_16;
    wire bfn_6_23_0_;
    wire blink_counterZ0Z_17;
    wire blink_counter_cry_16;
    wire blink_counterZ0Z_18;
    wire blink_counter_cry_17;
    wire blink_counterZ0Z_19;
    wire blink_counter_cry_18;
    wire blink_counterZ0Z_20;
    wire blink_counter_cry_19;
    wire blink_counter_cry_20;
    wire blink_counter_cry_21;
    wire blink_counter_cry_22;
    wire blink_counter_cry_23;
    wire bfn_6_24_0_;
    wire blink_counter_cry_24;
    wire \c0.rx.r_Rx_Bytece_0_2_cascade_ ;
    wire \c0.rx.N_325 ;
    wire \c0.rx.N_325_cascade_ ;
    wire \c0.rx.r_Rx_Bytece_0_5_cascade_ ;
    wire \c0.rx.N_388 ;
    wire \c0.rx.r_Rx_Bytece_0_6_cascade_ ;
    wire \c0.rx.r_Rx_Byte_1_sqmuxa ;
    wire \c0.rx.r_Rx_Bytece_0_0 ;
    wire \c0.rx.r_Rx_Byte_1_sqmuxa_cascade_ ;
    wire \c0.rx.r_Clock_Count_RNO_0_0_0 ;
    wire bfn_7_19_0_;
    wire \c0.rx.r_Clock_Count_RNO_0_0_1 ;
    wire \c0.rx.un1_r_Clock_Count_5_cry_0 ;
    wire \c0.rx.un1_r_Clock_Count_5_cry_1 ;
    wire \c0.rx.un1_r_Clock_Count_5_cry_2 ;
    wire \c0.rx.r_Clock_Count_RNO_0Z0Z_4 ;
    wire \c0.rx.un1_r_Clock_Count_5_cry_3 ;
    wire \c0.rx.un1_r_Clock_Count_5_cry_4 ;
    wire \c0.rx.r_Clock_Count_RNO_0Z0Z_6 ;
    wire \c0.rx.un1_r_Clock_Count_5_cry_5 ;
    wire \c0.rx.un1_r_Clock_Count_5_cry_6 ;
    wire \c0.rx.r_Clock_Count_RNO_0Z0Z_7 ;
    wire \c0.rx.r_Clock_CountZ1Z_1 ;
    wire \c0.rx.r_Clock_CountZ1Z_0 ;
    wire \c0.rx.N_320_cascade_ ;
    wire \c0.rx.r_Clock_Count_8_f0_0_o2_0_2_cascade_ ;
    wire \c0.rx.un1_r_Clock_Count_2_sqmuxa_0_i ;
    wire \c0.rx.r_Clock_Count_8_f0_0_o2_0_2 ;
    wire \c0.rx.r_Clock_Count_RNO_0_0_2 ;
    wire \c0.rx.N_332_cascade_ ;
    wire \c0.rx.r_Clock_CountZ1Z_2 ;
    wire \c0.rx.r_Clock_CountZ1Z_6 ;
    wire \c0.rx.r_Clock_CountZ0Z_7 ;
    wire \c0.rx.r_Clock_CountZ1Z_4 ;
    wire \c0.rx.r_Clock_Count_RNO_0Z0Z_5 ;
    wire \c0.rx.r_Clock_CountZ1Z_5 ;
    wire \c0.rx.N_320 ;
    wire \c0.rx.N_317 ;
    wire \c0.rx.N_337 ;
    wire \c0.rx.N_383_cascade_ ;
    wire \c0.rx.N_138r_0_i_1_cascade_ ;
    wire \c0.rx.r_SM_MainZ0Z_0 ;
    wire \c0.rx.N_91_0_cascade_ ;
    wire \c0.rx.r_SM_Main_illegal_0 ;
    wire \c0.rx.r_SM_Main_ns_0_i_a2_0_3_cascade_ ;
    wire \c0.rx.r_SM_Main_ns_0_i_a2_1_0_2 ;
    wire \c0.rx.r_SM_Main_dup_1 ;
    wire \c0.rx.un1_r_Rx_DV7_i_0_cascade_ ;
    wire \c0.rx.r_Rx_DV_RNOZ0Z_0 ;
    wire \c0.rx.r_SM_Main_dup_2 ;
    wire \c0.rx.r_SM_Main_ns_0_i_0_0_2 ;
    wire \c0.rx.r_Rx_DataZ0 ;
    wire \c0.rx.N_383 ;
    wire \c0.rx.N_321 ;
    wire \c0.rx.r_Clock_Count_8_f0_0_a2_0_0_2_cascade_ ;
    wire \c0.rx.N_371 ;
    wire \c0.rx.N_332 ;
    wire \c0.rx.r_SM_Main_RNI58REZ0Z_0 ;
    wire \c0.rx.N_361 ;
    wire \c0.rx.r_Clock_Count_RNO_0_0_3 ;
    wire \c0.rx.r_Clock_CountZ1Z_3 ;
    wire \c0.rx.N_386 ;
    wire \c0.rx.r_SM_Main_dup_3 ;
    wire \c0.rx.N_98_dup ;
    wire \c0.rx.r_SM_Main_dup_4 ;
    wire bfn_9_19_0_;
    wire \c0.i12_0 ;
    wire \c0.i12_1 ;
    wire \c0.i12_2 ;
    wire \c0.i12_3 ;
    wire \c0.i12_4 ;
    wire \c0.i12_5 ;
    wire \c0.i12_7_and ;
    wire \c0.i12_6 ;
    wire \c0.i12 ;
    wire bfn_9_20_0_;
    wire \c0.i12_0_and ;
    wire \c0.i12_1_and ;
    wire blink_counterZ0Z_21;
    wire blink_counterZ0Z_22;
    wire blink_counterZ0Z_24;
    wire N_12;
    wire blink_counterZ0Z_25;
    wire N_8_0_cascade_;
    wire blink_counterZ0Z_23;
    wire LED_c;
    wire \c0.tx.N_90_ip_RNIVJLQZ0_cascade_ ;
    wire \c0.tx.r_SM_Main_illegal_0 ;
    wire \c0.tx.N_90_dup_cascade_ ;
    wire \c0.tx.N_83_0 ;
    wire \c0.tx.r_Clock_Count_0_sqmuxa ;
    wire \c0.tx.r_Clock_Count_RNO_0Z0Z_0 ;
    wire bfn_9_23_0_;
    wire \c0.tx.r_Clock_Count_RNO_0Z0Z_1 ;
    wire \c0.tx.un1_r_Clock_Count_cry_0 ;
    wire \c0.tx.r_Clock_Count_RNO_0Z0Z_2 ;
    wire \c0.tx.un1_r_Clock_Count_cry_1 ;
    wire \c0.tx.un1_r_Clock_Count_cry_2 ;
    wire \c0.tx.r_Clock_Count_RNO_0Z0Z_3 ;
    wire \c0.tx.r_Clock_CountZ0Z_2 ;
    wire \c0.tx.r_Clock_CountZ0Z_1 ;
    wire \c0.tx.r_Clock_CountZ0Z_3 ;
    wire \c0.tx.r_Clock_CountZ0Z_0 ;
    wire \c0.tx.r_SM_Main_RNO_0Z0Z_1 ;
    wire \c0.tx.N_171_0_cascade_ ;
    wire \c0.nextCRC16_3_0_a2_1_8_cascade_ ;
    wire \c0.data_out_6_Z0Z_0 ;
    wire \c0.N_71 ;
    wire bfn_9_27_0_;
    wire \c0.dataZ0Z_1 ;
    wire \c0.data_cry_0 ;
    wire \c0.data_cry_1 ;
    wire \c0.dataZ0Z_3 ;
    wire \c0.data_cry_2 ;
    wire \c0.data_cry_3 ;
    wire \c0.dataZ0Z_5 ;
    wire \c0.data_cry_4 ;
    wire \c0.data_cry_5 ;
    wire \c0.dataZ0Z_7 ;
    wire \c0.data_cry_6 ;
    wire \c0.data_cry_7 ;
    wire bfn_9_28_0_;
    wire \c0.dataZ0Z_9 ;
    wire \c0.data_cry_8 ;
    wire \c0.dataZ0Z_10 ;
    wire \c0.data_cry_9 ;
    wire \c0.data_cry_10 ;
    wire \c0.data_cry_11 ;
    wire \c0.dataZ0Z_13 ;
    wire \c0.data_cry_12 ;
    wire \c0.data_cry_13 ;
    wire \c0.data_cry_14 ;
    wire \c0.i12_3_and ;
    wire \c0.i12_6_and ;
    wire \c0.i12_2_and ;
    wire \c0.i12_5_and ;
    wire \c0.i12_4_and ;
    wire \c0.tx.r_Bit_Index_RNO_0Z0Z_2_cascade_ ;
    wire \c0.tx.r_Tx_Active_1_sqmuxa_cascade_ ;
    wire \c0.tx.N_90_ip_RNIVJLQZ0 ;
    wire \c0.tx_active ;
    wire \c0.tx.N_90_ip_RNI1U1EZ0_cascade_ ;
    wire \c0.tx.r_SM_Main_dup_4 ;
    wire \c0.tx_transmitZ0 ;
    wire \c0.tx.r_SM_Main_RNO_0Z0Z_0 ;
    wire \c0.tx.N_171_0 ;
    wire \c0.tx.r_SM_Main_RNO_0Z0Z_2_cascade_ ;
    wire \c0.tx.r_SM_MainZ0Z_0 ;
    wire \c0.tx.N_90_dup ;
    wire \c0.tx.r_Clock_Count12_THRU_CO ;
    wire \c0.tx.r_SM_Main_RNIVDI71Z0Z_2 ;
    wire \c0.nextCRC16_3_0_a2_6_0_15 ;
    wire \c0.nextCRC16_3_9_cascade_ ;
    wire \c0.N_106_cascade_ ;
    wire \c0.N_92 ;
    wire \c0.N_106 ;
    wire \c0.data_out_7_Z0Z_0 ;
    wire \c0.nextCRC16_3_0_a2_0_10 ;
    wire \c0.dataZ0Z_12 ;
    wire \c0.N_77 ;
    wire \c0.N_76 ;
    wire \c0.dataZ0Z_0 ;
    wire \c0.dataZ0Z_14 ;
    wire \c0.dataZ0Z_11 ;
    wire \c0.dataZ0Z_2 ;
    wire \c0.dataZ0Z_15 ;
    wire \c0.dataZ0Z_4 ;
    wire \c0.dataZ0Z_8 ;
    wire \c0.data_in_0_Z0Z_4 ;
    wire \c0.data_in_1_Z0Z_0 ;
    wire \c0.rx_data_3 ;
    wire \c0.rx_data_1 ;
    wire \c0.rx_data_0 ;
    wire \c0.tx.o_Tx_Serial_2_3_i_m2_ns_1_cascade_ ;
    wire \c0.tx.N_90_ip_RNI1U1EZ0 ;
    wire \c0.tx.o_Tx_Serial_2_6_i_m2_ns_1_cascade_ ;
    wire \c0.tx.o_Tx_Serial_RNO_3_0 ;
    wire \c0.tx.o_Tx_Serial_RNO_2_0_cascade_ ;
    wire \c0.tx.r_SM_Main_RNI522EZ0Z_4 ;
    wire \c0.tx.o_Tx_Serial_RNOZ0Z_1_cascade_ ;
    wire \c0.tx.r_SM_Main_dup_3 ;
    wire PIN_1_c;
    wire \c0.tx.N_390_i ;
    wire \c0.tx.r_SM_Main_dup_2 ;
    wire \c0.tx.r_SM_Main_recr_i_0_a2_0_2_0_1_3 ;
    wire \c0.tx.r_Bit_IndexZ0Z_1 ;
    wire \c0.tx.r_Bit_IndexZ0Z_2 ;
    wire \c0.tx.r_SM_Main_dup_1 ;
    wire \c0.tx.r_Bit_IndexZ0Z_0 ;
    wire \c0.tx.r_SM_Main_recr_i_i_a2_0_1_2 ;
    wire \c0.data_out_7_Z0Z_5 ;
    wire \c0.tx_data_RNO_3Z0Z_3_cascade_ ;
    wire \c0.d_2_19 ;
    wire \c0.tx_data_RNO_4Z0Z_3 ;
    wire \c0.nextCRC16_3_0_a2_1_2_cascade_ ;
    wire \c0.dataZ0Z_6 ;
    wire \c0.N_99_cascade_ ;
    wire \c0.nextCRC16_3_0_a2_0_0 ;
    wire \c0.nextCRC16_3_0_a2_3_0_cascade_ ;
    wire \c0.nextCRC16_3_0_a2_4_0 ;
    wire \c0.d_2_27 ;
    wire \c0.N_81_cascade_ ;
    wire \c0.N_105 ;
    wire \c0.N_105_cascade_ ;
    wire \c0.data_out_6_Z0Z_5 ;
    wire \c0.nextCRC16_3_0_a2_1_15_cascade_ ;
    wire \c0.N_99 ;
    wire \c0.nextCRC16_3_0_a2_5_15 ;
    wire \c0.nextCRC16_3_0_a2_2_15 ;
    wire \c0.N_95_cascade_ ;
    wire \c0.N_85 ;
    wire \c0.nextCRC16_3_2_1 ;
    wire \c0.d_2_3 ;
    wire \c0.N_75 ;
    wire \c0.N_75_cascade_ ;
    wire \c0.N_93 ;
    wire \c0.d_2_35 ;
    wire \c0.rx_data_7 ;
    wire \c0.data_in_2_Z0Z_5 ;
    wire \c0.data_in_2_Z0Z_3 ;
    wire \c0.data_in_0_Z0Z_7 ;
    wire \c0.data_in_2_Z0Z_7 ;
    wire \c0.data_in_6_Z0Z_0 ;
    wire \c0.data_in_2_Z0Z_4 ;
    wire \c0.data_in_4_Z0Z_2 ;
    wire \c0.data_in_4_Z0Z_5 ;
    wire \c0.data_in_0_Z0Z_0 ;
    wire \c0.data_in_1_Z0Z_3 ;
    wire \c0.data_in_1_Z0Z_7 ;
    wire \c0.data_in_3_Z0Z_0 ;
    wire \c0.data_in_3_Z0Z_5 ;
    wire \c0.data_in_4_Z0Z_1 ;
    wire \c0.data_in_4_Z0Z_7 ;
    wire \c0.data_in_5_Z0Z_3 ;
    wire \c0.N_108_cascade_ ;
    wire \c0.N_122_cascade_ ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_2_cascade_ ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_4_cascade_ ;
    wire \c0.data_in_7_Z0Z_3 ;
    wire \c0.data_in_2_Z0Z_1 ;
    wire \c0.data_in_3_Z0Z_6 ;
    wire \c0.data_in_frame_7_Z0Z_3 ;
    wire \c0.data_in_6_Z0Z_3 ;
    wire \c0.data_in_frame_6_Z0Z_3 ;
    wire \c0.d_4_17 ;
    wire \c0.tx2_data_RNO_4Z0Z_1 ;
    wire \c0.m161_ns_1_cascade_ ;
    wire \c0.tx2_data_RNO_0Z0Z_1 ;
    wire \c0.tx2_data_RNO_0Z0Z_2_cascade_ ;
    wire \c0.data_in_frame_6_Z0Z_2 ;
    wire \c0.data_in_frame_7_Z0Z_2 ;
    wire \c0.tx2_data_RNO_1Z0Z_2 ;
    wire \c0.tx_data_RNO_0Z0Z_3 ;
    wire \c0.tx_data_1_0_i_ns_1_3 ;
    wire \c0.tx.r_Tx_DataZ0Z_3 ;
    wire \c0.d_2_7 ;
    wire \c0.tx_data_RNO_3Z0Z_7_cascade_ ;
    wire \c0.tx_data_RNO_4Z0Z_7 ;
    wire \c0.tx_data_1_0_i_ns_1_7_cascade_ ;
    wire \c0.tx.r_Tx_DataZ0Z_7 ;
    wire \c0.tx.r_Tx_DataZ0Z_4 ;
    wire \c0.tx_data_RNO_1Z0Z_5 ;
    wire \c0.tx.r_Tx_DataZ0Z_5 ;
    wire \c0.N_24_0 ;
    wire \c0.un144_newcrc_2 ;
    wire \c0.un144_newcrc_5_cascade_ ;
    wire \c0.data_out_7_Z0Z_6 ;
    wire \c0.N_81 ;
    wire \c0.data_out_6_Z0Z_6 ;
    wire \c0.tx_data_RNO_3Z0Z_4_cascade_ ;
    wire \c0.tx_data_1_0_i_ns_1_4 ;
    wire \c0.d_2_20 ;
    wire \c0.tx_data_RNO_4Z0Z_4 ;
    wire \c0.N_95 ;
    wire \c0.d_2_8 ;
    wire \c0.d_2_0 ;
    wire \c0.tx_data_RNO_3Z0Z_0_cascade_ ;
    wire \c0.tx_data_RNO_4Z0Z_0 ;
    wire \c0.d_2_33 ;
    wire \c0.d_2_34 ;
    wire \c0.d_2_15 ;
    wire \c0.d_2_43 ;
    wire \c0.un105_newcrc_0_a2_0_cascade_ ;
    wire \c0.N_100 ;
    wire \c0.d_2_31 ;
    wire \c0.un105_newcrc_0_a2_3 ;
    wire \c0.d_2_32 ;
    wire \c0.d_2_24 ;
    wire \c0.nextCRC16_3_3_12 ;
    wire \c0.nextCRC16_3_4_12_cascade_ ;
    wire \c0.d_2_41 ;
    wire \c0.N_94 ;
    wire \c0.N_94_cascade_ ;
    wire \c0.d_2_23 ;
    wire \c0.d_2_40 ;
    wire \c0.nextCRC16_3_0_a2_1_11 ;
    wire \c0.data_out_6_Z0Z_4 ;
    wire \c0.data_out_7_Z0Z_4 ;
    wire \c0.tx_data_RNO_1Z0Z_4 ;
    wire \c0.data_in_5_Z0Z_5 ;
    wire \c0.rx_data_4 ;
    wire \c0.rx_data_2 ;
    wire \c0.d_4_34 ;
    wire \c0.un1_data_in_7__7_0_a2_0_a2_2_cascade_ ;
    wire \c0.un1_data_in_6__0_0_a2_5_a2_2 ;
    wire \c0.un1_data_in_7__7_i_cascade_ ;
    wire \c0.data_in_5_Z0Z_7 ;
    wire \c0.data_in_4_Z0Z_3 ;
    wire \c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_ ;
    wire \c0.data_in_3_Z0Z_4 ;
    wire \c0.data_in_1_Z0Z_5 ;
    wire \c0.data_in_3_Z0Z_2 ;
    wire \c0.data_in_5_Z0Z_1 ;
    wire \c0.data_in_5_Z0Z_0 ;
    wire \c0.N_132 ;
    wire \c0.un1_data_in_7__0_0_a2_1_a2_5_cascade_ ;
    wire \c0.N_121_cascade_ ;
    wire \c0.N_125 ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_4_3_cascade_ ;
    wire \c0.N_136 ;
    wire \c0.N_136_cascade_ ;
    wire \c0.un1_data_in_7__0_0_a2_1_a2_2 ;
    wire \c0.data_in_3_Z0Z_3 ;
    wire \c0.un1_data_in_7__1_0_a2_24_a2_3_cascade_ ;
    wire \c0.un1_data_in_7__1_0_a2_24_a2_4 ;
    wire \c0.data_in_5_Z0Z_4 ;
    wire \c0.data_in_5_Z0Z_2 ;
    wire \c0.data_in_2_Z0Z_0 ;
    wire \c0.d_4_33 ;
    wire \c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_ ;
    wire \c0.N_124 ;
    wire \c0.N_124_cascade_ ;
    wire \c0.N_108 ;
    wire \c0.un1_data_in_7__6_0_a2_5_a2_2_cascade_ ;
    wire \c0.un1_data_in_7__4_0_a2_0_a2_4 ;
    wire \c0.data_in_0_Z0Z_3 ;
    wire \c0.data_in_0_Z0Z_5 ;
    wire \c0.data_in_2_Z0Z_2 ;
    wire \c0.d_4_18 ;
    wire \c0.d_2_38 ;
    wire \c0.d_2_46 ;
    wire \c0.data_out_6_Z0Z_7 ;
    wire \c0.data_out_7_Z0Z_7 ;
    wire \c0.tx_data_RNO_1Z0Z_7 ;
    wire \c0.d_2_37 ;
    wire \c0.d_2_45 ;
    wire \c0.tx_data_RNO_0Z0Z_5 ;
    wire \c0.tx_data_RNO_3Z0Z_6_cascade_ ;
    wire \c0.tx_data_RNO_4Z0Z_6 ;
    wire \c0.d_2_42 ;
    wire \c0.nextCRC16_3_3_1 ;
    wire \c0.d_2_4 ;
    wire \c0.nextCRC16_3_3_1_cascade_ ;
    wire \c0.nextCRC16_3_0_a2_1_1 ;
    wire \c0.d_2_28 ;
    wire \c0.d_2_5 ;
    wire \c0.d_2_13 ;
    wire \c0.tx_data_RNO_3Z0Z_5_cascade_ ;
    wire \c0.tx_data_1_0_i_ns_1_5 ;
    wire \c0.tx_data_RNO_4Z0Z_5 ;
    wire \c0.tx_data_RNO_1Z0Z_0 ;
    wire \c0.tx_data_RNO_0Z0Z_0 ;
    wire \c0.tx_data_1_0_i_ns_1_0 ;
    wire \c0.tx.r_Tx_DataZ0Z_0 ;
    wire \c0.tx_data_RNO_0Z0Z_2 ;
    wire \c0.tx.r_Tx_DataZ0Z_2 ;
    wire \c0.d_2_25 ;
    wire \c0.tx_data_RNO_4Z0Z_1_cascade_ ;
    wire \c0.tx_data_RNO_0Z0Z_1 ;
    wire \c0.tx_data_1_0_i_ns_1_1_cascade_ ;
    wire \c0.tx.r_Tx_DataZ0Z_1 ;
    wire \c0.data_out_7_Z0Z_2 ;
    wire \c0.data_out_6_Z0Z_2 ;
    wire \c0.tx_data_RNO_1Z0Z_2 ;
    wire \c0.d_2_1 ;
    wire \c0.d_2_9 ;
    wire \c0.tx_data_RNO_3Z0Z_1 ;
    wire \c0.d_2_2 ;
    wire \c0.tx_data_RNO_3Z0Z_2_cascade_ ;
    wire \c0.tx_data_RNO_4Z0Z_2 ;
    wire \c0.tx_data_1_0_i_ns_1_2 ;
    wire \c0.d_2_39 ;
    wire \c0.d_2_47 ;
    wire \c0.tx_data_RNO_0Z0Z_7 ;
    wire \c0.d_2_36 ;
    wire \c0.d_2_44 ;
    wire \c0.tx_data_RNO_0Z0Z_4 ;
    wire \c0.data_out_6_Z0Z_1 ;
    wire \c0.data_out_7_Z0Z_1 ;
    wire \c0.tx_data_RNO_1Z0Z_1 ;
    wire \c0.m2_e_1_cascade_ ;
    wire \c0.data_out_7_Z0Z_3 ;
    wire \c0.data_out_6_Z0Z_3 ;
    wire \c0.N_132_mux_cascade_ ;
    wire \c0.tx_data_RNO_1Z0Z_3 ;
    wire \c0.byte_transmit_counterZ0Z_5 ;
    wire \c0.data_in_6_Z0Z_7 ;
    wire \c0.data_in_frame_6_Z0Z_7 ;
    wire \c0.data_in_7_Z0Z_7 ;
    wire \c0.data_in_frame_7_Z0Z_7 ;
    wire \c0.data_in_0_Z0Z_6 ;
    wire \c0.d_4_6 ;
    wire \c0.N_109 ;
    wire \c0.data_in_1_Z0Z_6 ;
    wire \c0.d_4_7 ;
    wire \c0.tx2_data_RNO_3Z0Z_7 ;
    wire \c0.data_in_4_Z0Z_4 ;
    wire \c0.data_in_6_Z0Z_1 ;
    wire \c0.N_34_cascade_ ;
    wire \c0.data_in_2_Z0Z_6 ;
    wire \c0.d_4_44 ;
    wire \c0.d_4_36 ;
    wire \c0.N_104 ;
    wire \c0.un1_data_in_6__3_0_a2_5_a2_2 ;
    wire \c0.un1_data_in_6__5_cascade_ ;
    wire \c0.un1_data_in_6__6 ;
    wire \c0.un1_data_in_6__1_0_a2_4_a2_2 ;
    wire \c0.m163_2_cascade_ ;
    wire \c0.N_126 ;
    wire \c0.m163_7_cascade_ ;
    wire \c0.m163_0 ;
    wire \c0.un1_data_in_6__5_0_a2_5_a2_2 ;
    wire \c0.N_120 ;
    wire \c0.data_in_1_Z0Z_4 ;
    wire \c0.N_121 ;
    wire \c0.m163_4 ;
    wire \c0.un1_data_in_7__1_0_a2_24_a2_7 ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_6 ;
    wire \c0.m163_8_cascade_ ;
    wire \c0.un1_data_in_7__1_3 ;
    wire \c0.m163_10 ;
    wire \c0.m163_1_cascade_ ;
    wire \c0.un1_data_in_7__0 ;
    wire \c0.N_164_0_cascade_ ;
    wire \c0.N_173_0_cascade_ ;
    wire \c0.data_in_3_Z0Z_7 ;
    wire \c0.d_4_RNIB3JJZ0Z_2 ;
    wire \c0.data_in_0_Z0Z_2 ;
    wire \c0.data_in_4_Z0Z_0 ;
    wire \c0.d_4_23 ;
    wire \c0.tx2_data_RNO_4Z0Z_7 ;
    wire \c0.d_4_2 ;
    wire \c0.tx2_data_RNO_4Z0Z_2 ;
    wire \c0.tx2_data_RNO_3Z0Z_2_cascade_ ;
    wire \c0.m131_ns_1 ;
    wire \c0.tx_data_RNO_1Z0Z_6 ;
    wire \c0.tx_data_RNO_0Z0Z_6 ;
    wire \c0.tx_data_1_0_i_ns_1_6 ;
    wire \c0.tx.r_Tx_DataZ0Z_6 ;
    wire \c0.tx.N_398_i ;
    wire \c0.rx.r_Bit_IndexZ0Z_1 ;
    wire \c0.rx.r_Bit_IndexZ0Z_2 ;
    wire \c0.rx.r_Bit_IndexZ0Z_0 ;
    wire \c0.rx.N_335 ;
    wire \c0.d_4_35 ;
    wire \c0.d_4_27 ;
    wire \c0.d_4_19 ;
    wire \c0.d_4_3 ;
    wire \c0.d_4_11 ;
    wire \c0.tx2_data_RNO_4Z0Z_3 ;
    wire \c0.tx2_data_RNO_3Z0Z_3_cascade_ ;
    wire \c0.tx2_data_RNO_0Z0Z_3 ;
    wire \c0.m105_ns_1_cascade_ ;
    wire \c0.tx2_data_RNO_1Z0Z_3 ;
    wire \c0.tx2.r_Tx_DataZ0Z_3 ;
    wire \c0.tx2_data_RNO_1Z0Z_7 ;
    wire \c0.m60_0_ns_1 ;
    wire \c0.tx2.r_Tx_DataZ0Z_7 ;
    wire \c0.d_2_6 ;
    wire \c0.d_2_22 ;
    wire \c0.d_2_14 ;
    wire \c0.d_2_30 ;
    wire \c0.d_2_16 ;
    wire \c0.d_2_17 ;
    wire \c0.d_2_12 ;
    wire \c0.d_2_21 ;
    wire \c0.d_2_11 ;
    wire \c0.d_2_26 ;
    wire \c0.d_2_18 ;
    wire \c0.d_2_10 ;
    wire \c0.byte_transmit_counterZ0Z_6 ;
    wire \c0.byte_transmit_counterZ0Z_7 ;
    wire \c0.byte_transmit_counterZ0Z_3 ;
    wire GNDG0;
    wire \c0.byte_transmit_counterZ0Z_4 ;
    wire \c0.byte_transmit_counterZ0Z_1 ;
    wire \c0.byte_transmit_counterZ0Z_0 ;
    wire \c0.N_132_mux ;
    wire \c0.byte_transmit_counterZ0Z_2 ;
    wire \c0.N_5_1_cascade_ ;
    wire \c0.byte_transmit_counter15 ;
    wire \c0.data_out_0__1_sqmuxa ;
    wire \c0.data_in_frame_6_Z0Z_4 ;
    wire \c0.data_in_frame_7_Z0Z_4 ;
    wire \c0.tx2_data_RNO_1Z0Z_4 ;
    wire \c0.tx2_data_RNO_0Z0Z_4 ;
    wire \c0.m120_ns_1_cascade_ ;
    wire \c0.tx2_data_RNO_3Z0Z_6 ;
    wire \c0.tx2_data_RNO_0Z0Z_6 ;
    wire \c0.m90_ns_1_cascade_ ;
    wire \c0.tx2_data_RNO_1Z0Z_6 ;
    wire \c0.data_in_7_Z0Z_4 ;
    wire \c0.rx_data_5 ;
    wire \c0.data_in_4_Z0Z_6 ;
    wire \c0.data_in_5_Z0Z_6 ;
    wire \c0.rx_data_6 ;
    wire \c0.d_4_26 ;
    wire \c0.data_in_6_Z0Z_4 ;
    wire \c0.d_4_41 ;
    wire \c0.un1_data_in_6__4_0_a2_5_a2_1 ;
    wire \c0.data_in_1_Z0Z_2 ;
    wire \c0.d_4_10 ;
    wire \c0.N_127 ;
    wire \c0.data_in_1_Z0Z_1 ;
    wire \c0.data_in_3_Z0Z_1 ;
    wire \c0.d_4_25 ;
    wire \c0.d_4_38 ;
    wire \c0.N_107 ;
    wire \c0.un1_data_in_6__2_0_a2_6_a2_2_cascade_ ;
    wire \c0.un1_data_in_6__2 ;
    wire \c0.d_4_46 ;
    wire \c0.d_4_42 ;
    wire \c0.N_133 ;
    wire \c0.un1_data_in_7__2_0_a2_0_a2_5_cascade_ ;
    wire \c0.un1_data_in_7__2 ;
    wire \c0.d_4_14 ;
    wire \c0.d_4_31 ;
    wire \c0.un1_data_in_7__2_0_a2_0_a2_4 ;
    wire \c0.un1_data_in_7__3_0_a2_0_a2_3 ;
    wire \c0.d_4_43 ;
    wire \c0.N_128 ;
    wire \c0.un1_data_in_7__3_0_a2_0_a2_4_cascade_ ;
    wire \c0.un1_data_in_7__5_0_a2_0_a2_1 ;
    wire \c0.m163_9 ;
    wire \c0.data_in_0_Z0Z_1 ;
    wire \c0.N_123 ;
    wire \c0.d_4_15 ;
    wire \c0.N_129 ;
    wire \c0.N_18 ;
    wire bfn_15_21_0_;
    wire \c0.un1_byte_transmit_counter2_1_cry_0 ;
    wire \c0.un1_byte_transmit_counter2_1_cry_1 ;
    wire \c0.un1_byte_transmit_counter2_1_cry_2 ;
    wire \c0.un1_byte_transmit_counter2_1_cry_3 ;
    wire \c0.un1_byte_transmit_counter2_1_cry_4 ;
    wire \c0.un1_byte_transmit_counter2_1_cry_5 ;
    wire \c0.un1_byte_transmit_counter2_1_cry_6 ;
    wire \c0.d_4_1 ;
    wire \c0.d_4_9 ;
    wire \c0.tx2_data_RNO_3Z0Z_1 ;
    wire \c0.tx2.r_Tx_DataZ0Z_1 ;
    wire \c0.data_in_frame_6_Z0Z_1 ;
    wire \c0.tx2_data_RNO_1Z0Z_1 ;
    wire \c0.tx2.r_Tx_DataZ0Z_4 ;
    wire \c0.N_173_0 ;
    wire \c0.tx2.r_Clock_Count_i_0 ;
    wire bfn_15_23_0_;
    wire \c0.tx2.r_Clock_Count_i_1 ;
    wire \c0.tx2.r_Clock_Count12_cry_0 ;
    wire \c0.tx2.r_Clock_Count_i_2 ;
    wire \c0.tx2.r_Clock_Count12_cry_1 ;
    wire \c0.tx2.r_Clock_Count_i_3 ;
    wire \c0.tx2.r_Clock_Count12_cry_2 ;
    wire \c0.tx2.r_Clock_Count12 ;
    wire CONSTANT_ONE_NET;
    wire \c0.d_2_29 ;
    wire \c0.data_out_0__1_sqmuxa_g ;
    wire \c0.tx2.r_Tx_DataZ0Z_6 ;
    wire \c0.tx2.r_Tx_DataZ0Z_2 ;
    wire \c0.tx2.o_Tx_Serial_RNOZ0Z_6_cascade_ ;
    wire \c0.tx2.o_Tx_Serial_RNOZ0Z_5 ;
    wire \c0.tx2.o_Tx_Serial_RNOZ0Z_3 ;
    wire \c0.tx2.m195_ns_1_cascade_ ;
    wire \c0.tx2.o_Tx_Serial_RNOZ0Z_2 ;
    wire \c0.tx2.N_196_0_cascade_ ;
    wire \c0.tx2.N_493_cascade_ ;
    wire \c0.tx2.N_205_mux ;
    wire PIN_3_c;
    wire \c0.data_in_7_Z0Z_0 ;
    wire \c0.data_in_7_Z0Z_1 ;
    wire \c0.data_in_frame_7_Z0Z_1 ;
    wire \c0.data_in_6_Z0Z_5 ;
    wire \c0.data_in_7_Z0Z_5 ;
    wire \c0.data_in_7_Z0Z_6 ;
    wire \c0.data_in_frame_7_Z0Z_6 ;
    wire \c0.data_in_6_Z0Z_6 ;
    wire \c0.data_in_frame_6_Z0Z_6 ;
    wire \c0.data_in_frame_0__0_sqmuxa_g ;
    wire \c0.data_in_7_Z0Z_2 ;
    wire \c0.data_in_6_Z0Z_2 ;
    wire \c0.rx_data_ready_g ;
    wire \c0.d_4_45 ;
    wire \c0.d_4_37 ;
    wire \c0.d_4_29 ;
    wire \c0.d_4_21 ;
    wire \c0.tx2_data_RNO_4Z0Z_5_cascade_ ;
    wire \c0.tx2_data_RNO_0Z0Z_5 ;
    wire \c0.m75_ns_1_cascade_ ;
    wire \c0.tx2.r_Tx_DataZ0Z_5 ;
    wire \c0.data_in_frame_6_Z0Z_5 ;
    wire \c0.data_in_frame_7_Z0Z_5 ;
    wire \c0.tx2_data_RNO_1Z0Z_5 ;
    wire \c0.d_4_47 ;
    wire \c0.d_4_39 ;
    wire \c0.tx2_data_RNO_0Z0Z_7 ;
    wire \c0.data_in_frame_6_Z0Z_0 ;
    wire \c0.data_in_frame_7_Z0Z_0 ;
    wire \c0.N_164_0 ;
    wire \c0.d_4_22 ;
    wire \c0.d_4_30 ;
    wire \c0.tx2_data_RNO_4Z0Z_6 ;
    wire \c0.d_4_4 ;
    wire \c0.d_4_12 ;
    wire \c0.tx2_data_RNO_3Z0Z_4 ;
    wire \c0.d_4_28 ;
    wire \c0.d_4_20 ;
    wire \c0.tx2_data_RNO_4Z0Z_4 ;
    wire \c0.d_4_13 ;
    wire \c0.d_4_5 ;
    wire \c0.tx2_data_RNO_3Z0Z_5 ;
    wire \c0.byte_transmit_counter2Z0Z_7 ;
    wire \c0.byte_transmit_counter2Z0Z_3 ;
    wire \c0.byte_transmit_counter2Z0Z_6 ;
    wire \c0.byte_transmit_counter2Z0Z_5 ;
    wire \c0.m45_0_0_cascade_ ;
    wire \c0.byte_transmit_counter2Z0Z_4 ;
    wire \c0.N_204_mux_cascade_ ;
    wire \c0.N_215_mux ;
    wire \c0.d_4_0 ;
    wire \c0.d_4_8 ;
    wire \c0.d_4_16 ;
    wire \c0.d_4_24 ;
    wire \c0.byte_transmit_counter2Z0Z_1 ;
    wire \c0.tx2_data_RNO_3Z0Z_0 ;
    wire \c0.tx2_data_RNO_4Z0Z_0_cascade_ ;
    wire \c0.byte_transmit_counter2Z0Z_2 ;
    wire \c0.tx2_data_RNO_1Z0Z_0 ;
    wire \c0.m146_ns_1_cascade_ ;
    wire \c0.tx2.r_Tx_DataZ0Z_0 ;
    wire \c0.byte_transmit_counter2Z0Z_0 ;
    wire \c0.d_4_32 ;
    wire \c0.N_204_mux ;
    wire \c0.d_4_40 ;
    wire \c0.tx2_data_RNO_0Z0Z_0 ;
    wire bfn_16_22_0_;
    wire \c0.tx2.un1_r_Clock_Count_cry_0 ;
    wire \c0.tx2.un1_r_Clock_Count_cry_1 ;
    wire \c0.tx2.un1_r_Clock_Count_cry_2 ;
    wire \c0.tx2.r_Clock_CountZ0Z_2 ;
    wire \c0.tx2.r_Clock_CountZ0Z_1 ;
    wire \c0.tx2.r_Clock_CountZ0Z_3 ;
    wire \c0.tx2.r_Clock_CountZ0Z_0 ;
    wire \c0.tx2.N_16_0 ;
    wire \c0.tx2.r_Clock_Count_0_sqmuxa ;
    wire \c0.tx2.N_83_0_cascade_ ;
    wire \c0.N_90_dup_cascade_ ;
    wire \c0.tx2.i97_mux_cascade_ ;
    wire \c0.tx2.r_SM_Main_illegal_0 ;
    wire \c0.tx2.N_214_0 ;
    wire \c0.tx2.r_Clock_Count12_THRU_CO ;
    wire \c0.tx2.N_17_0_cascade_ ;
    wire \c0.tx2.r_SM_Main_dup_4 ;
    wire \c0.tx2.r_Bit_IndexZ1Z_0 ;
    wire \c0.tx2.N_212_0_cascade_ ;
    wire \c0.tx2.r_SM_Main_dup_1 ;
    wire \c0.tx2.N_496_cascade_ ;
    wire \c0.tx2.r_SM_Main_dup_2 ;
    wire \c0.tx2.N_171_0 ;
    wire \c0.tx2.N_17_0 ;
    wire \c0.tx2.N_212_0 ;
    wire \c0.tx2.N_493 ;
    wire \c0.tx2.r_SM_Main_dup_3 ;
    wire \c0.tx2_transmitZ0 ;
    wire \c0.N_19_0 ;
    wire \c0.r_SM_Main_0 ;
    wire \c0.N_90_dup ;
    wire \c0.tx2.N_9_1_cascade_ ;
    wire \c0.tx2.r_Bit_IndexZ0Z_2 ;
    wire \c0.tx2.N_12_0 ;
    wire \c0.tx2.N_9_1 ;
    wire \c0.tx2.r_Bit_IndexZ0Z_1 ;
    wire \c0.tx2_active ;
    wire \c0.N_170_0 ;
    wire CLK_c_g;
    wire \c0.tx2_transmit_0_sqmuxa ;
    wire \c0.wait_for_transmissionZ0 ;
    wire \c0.i12_THRU_CO ;
    wire \c0.data_in_frame_0__0_sqmuxa ;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__20078),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__20080),
            .DIN(N__20079),
            .DOUT(N__20078),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__20080),
            .PADOUT(N__20079),
            .PADIN(N__20078),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD LED_obuf_iopad (
            .OE(N__20069),
            .DIN(N__20068),
            .DOUT(N__20067),
            .PACKAGEPIN(LED));
    defparam LED_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_preio (
            .PADOEN(N__20069),
            .PADOUT(N__20068),
            .PADIN(N__20067),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__9190),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PIN_1_obuf_iopad (
            .OE(N__20060),
            .DIN(N__20059),
            .DOUT(N__20058),
            .PACKAGEPIN(PIN_1));
    defparam PIN_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIN_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIN_1_obuf_preio (
            .PADOEN(N__20060),
            .PADOUT(N__20059),
            .PADIN(N__20058),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10288),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PIN_2_ibuf_iopad (
            .OE(N__20051),
            .DIN(N__20050),
            .DOUT(N__20049),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PIN_2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PIN_2_ibuf_preio (
            .PADOEN(N__20051),
            .PADOUT(N__20050),
            .PADIN(N__20049),
            .CLOCKENABLE(),
            .DIN0(PIN_2_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PIN_3_obuf_iopad (
            .OE(N__20042),
            .DIN(N__20041),
            .DOUT(N__20040),
            .PACKAGEPIN(PIN_3));
    defparam PIN_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIN_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIN_3_obuf_preio (
            .PADOEN(N__20042),
            .PADOUT(N__20041),
            .PADIN(N__20040),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__17404),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD USBPU_obuf_iopad (
            .OE(N__20033),
            .DIN(N__20032),
            .DOUT(N__20031),
            .PACKAGEPIN(USBPU));
    defparam USBPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam USBPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO USBPU_obuf_preio (
            .PADOEN(N__20033),
            .PADOUT(N__20032),
            .PADIN(N__20031),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__4707 (
            .O(N__20014),
            .I(N__20008));
    InMux I__4706 (
            .O(N__20013),
            .I(N__20005));
    InMux I__4705 (
            .O(N__20012),
            .I(N__20002));
    InMux I__4704 (
            .O(N__20011),
            .I(N__19999));
    LocalMux I__4703 (
            .O(N__20008),
            .I(N__19996));
    LocalMux I__4702 (
            .O(N__20005),
            .I(N__19993));
    LocalMux I__4701 (
            .O(N__20002),
            .I(N__19990));
    LocalMux I__4700 (
            .O(N__19999),
            .I(N__19983));
    Span4Mux_v I__4699 (
            .O(N__19996),
            .I(N__19983));
    Span4Mux_h I__4698 (
            .O(N__19993),
            .I(N__19983));
    Odrv4 I__4697 (
            .O(N__19990),
            .I(\c0.tx2_transmitZ0 ));
    Odrv4 I__4696 (
            .O(N__19983),
            .I(\c0.tx2_transmitZ0 ));
    CEMux I__4695 (
            .O(N__19978),
            .I(N__19974));
    CEMux I__4694 (
            .O(N__19977),
            .I(N__19970));
    LocalMux I__4693 (
            .O(N__19974),
            .I(N__19965));
    CEMux I__4692 (
            .O(N__19973),
            .I(N__19962));
    LocalMux I__4691 (
            .O(N__19970),
            .I(N__19959));
    CEMux I__4690 (
            .O(N__19969),
            .I(N__19956));
    CEMux I__4689 (
            .O(N__19968),
            .I(N__19953));
    Span4Mux_v I__4688 (
            .O(N__19965),
            .I(N__19947));
    LocalMux I__4687 (
            .O(N__19962),
            .I(N__19947));
    Span4Mux_h I__4686 (
            .O(N__19959),
            .I(N__19941));
    LocalMux I__4685 (
            .O(N__19956),
            .I(N__19941));
    LocalMux I__4684 (
            .O(N__19953),
            .I(N__19938));
    InMux I__4683 (
            .O(N__19952),
            .I(N__19935));
    Span4Mux_h I__4682 (
            .O(N__19947),
            .I(N__19932));
    InMux I__4681 (
            .O(N__19946),
            .I(N__19929));
    Span4Mux_v I__4680 (
            .O(N__19941),
            .I(N__19922));
    Span4Mux_h I__4679 (
            .O(N__19938),
            .I(N__19922));
    LocalMux I__4678 (
            .O(N__19935),
            .I(N__19922));
    Odrv4 I__4677 (
            .O(N__19932),
            .I(\c0.N_19_0 ));
    LocalMux I__4676 (
            .O(N__19929),
            .I(\c0.N_19_0 ));
    Odrv4 I__4675 (
            .O(N__19922),
            .I(\c0.N_19_0 ));
    CascadeMux I__4674 (
            .O(N__19915),
            .I(N__19909));
    InMux I__4673 (
            .O(N__19914),
            .I(N__19904));
    InMux I__4672 (
            .O(N__19913),
            .I(N__19904));
    CascadeMux I__4671 (
            .O(N__19912),
            .I(N__19900));
    InMux I__4670 (
            .O(N__19909),
            .I(N__19895));
    LocalMux I__4669 (
            .O(N__19904),
            .I(N__19892));
    InMux I__4668 (
            .O(N__19903),
            .I(N__19883));
    InMux I__4667 (
            .O(N__19900),
            .I(N__19883));
    InMux I__4666 (
            .O(N__19899),
            .I(N__19883));
    InMux I__4665 (
            .O(N__19898),
            .I(N__19883));
    LocalMux I__4664 (
            .O(N__19895),
            .I(\c0.r_SM_Main_0 ));
    Odrv4 I__4663 (
            .O(N__19892),
            .I(\c0.r_SM_Main_0 ));
    LocalMux I__4662 (
            .O(N__19883),
            .I(\c0.r_SM_Main_0 ));
    CascadeMux I__4661 (
            .O(N__19876),
            .I(N__19872));
    InMux I__4660 (
            .O(N__19875),
            .I(N__19867));
    InMux I__4659 (
            .O(N__19872),
            .I(N__19862));
    InMux I__4658 (
            .O(N__19871),
            .I(N__19862));
    InMux I__4657 (
            .O(N__19870),
            .I(N__19853));
    LocalMux I__4656 (
            .O(N__19867),
            .I(N__19848));
    LocalMux I__4655 (
            .O(N__19862),
            .I(N__19848));
    InMux I__4654 (
            .O(N__19861),
            .I(N__19841));
    InMux I__4653 (
            .O(N__19860),
            .I(N__19841));
    InMux I__4652 (
            .O(N__19859),
            .I(N__19841));
    InMux I__4651 (
            .O(N__19858),
            .I(N__19834));
    InMux I__4650 (
            .O(N__19857),
            .I(N__19834));
    InMux I__4649 (
            .O(N__19856),
            .I(N__19834));
    LocalMux I__4648 (
            .O(N__19853),
            .I(\c0.N_90_dup ));
    Odrv4 I__4647 (
            .O(N__19848),
            .I(\c0.N_90_dup ));
    LocalMux I__4646 (
            .O(N__19841),
            .I(\c0.N_90_dup ));
    LocalMux I__4645 (
            .O(N__19834),
            .I(\c0.N_90_dup ));
    CascadeMux I__4644 (
            .O(N__19825),
            .I(\c0.tx2.N_9_1_cascade_ ));
    InMux I__4643 (
            .O(N__19822),
            .I(N__19819));
    LocalMux I__4642 (
            .O(N__19819),
            .I(N__19812));
    InMux I__4641 (
            .O(N__19818),
            .I(N__19806));
    InMux I__4640 (
            .O(N__19817),
            .I(N__19806));
    InMux I__4639 (
            .O(N__19816),
            .I(N__19803));
    InMux I__4638 (
            .O(N__19815),
            .I(N__19800));
    Span4Mux_v I__4637 (
            .O(N__19812),
            .I(N__19797));
    InMux I__4636 (
            .O(N__19811),
            .I(N__19794));
    LocalMux I__4635 (
            .O(N__19806),
            .I(N__19791));
    LocalMux I__4634 (
            .O(N__19803),
            .I(\c0.tx2.r_Bit_IndexZ0Z_2 ));
    LocalMux I__4633 (
            .O(N__19800),
            .I(\c0.tx2.r_Bit_IndexZ0Z_2 ));
    Odrv4 I__4632 (
            .O(N__19797),
            .I(\c0.tx2.r_Bit_IndexZ0Z_2 ));
    LocalMux I__4631 (
            .O(N__19794),
            .I(\c0.tx2.r_Bit_IndexZ0Z_2 ));
    Odrv4 I__4630 (
            .O(N__19791),
            .I(\c0.tx2.r_Bit_IndexZ0Z_2 ));
    InMux I__4629 (
            .O(N__19780),
            .I(N__19774));
    InMux I__4628 (
            .O(N__19779),
            .I(N__19774));
    LocalMux I__4627 (
            .O(N__19774),
            .I(\c0.tx2.N_12_0 ));
    SRMux I__4626 (
            .O(N__19771),
            .I(N__19768));
    LocalMux I__4625 (
            .O(N__19768),
            .I(N__19765));
    Sp12to4 I__4624 (
            .O(N__19765),
            .I(N__19760));
    InMux I__4623 (
            .O(N__19764),
            .I(N__19757));
    InMux I__4622 (
            .O(N__19763),
            .I(N__19754));
    Odrv12 I__4621 (
            .O(N__19760),
            .I(\c0.tx2.N_9_1 ));
    LocalMux I__4620 (
            .O(N__19757),
            .I(\c0.tx2.N_9_1 ));
    LocalMux I__4619 (
            .O(N__19754),
            .I(\c0.tx2.N_9_1 ));
    InMux I__4618 (
            .O(N__19747),
            .I(N__19742));
    InMux I__4617 (
            .O(N__19746),
            .I(N__19736));
    InMux I__4616 (
            .O(N__19745),
            .I(N__19736));
    LocalMux I__4615 (
            .O(N__19742),
            .I(N__19733));
    InMux I__4614 (
            .O(N__19741),
            .I(N__19730));
    LocalMux I__4613 (
            .O(N__19736),
            .I(\c0.tx2.r_Bit_IndexZ0Z_1 ));
    Odrv4 I__4612 (
            .O(N__19733),
            .I(\c0.tx2.r_Bit_IndexZ0Z_1 ));
    LocalMux I__4611 (
            .O(N__19730),
            .I(\c0.tx2.r_Bit_IndexZ0Z_1 ));
    InMux I__4610 (
            .O(N__19723),
            .I(N__19717));
    InMux I__4609 (
            .O(N__19722),
            .I(N__19714));
    InMux I__4608 (
            .O(N__19721),
            .I(N__19711));
    CascadeMux I__4607 (
            .O(N__19720),
            .I(N__19708));
    LocalMux I__4606 (
            .O(N__19717),
            .I(N__19705));
    LocalMux I__4605 (
            .O(N__19714),
            .I(N__19700));
    LocalMux I__4604 (
            .O(N__19711),
            .I(N__19700));
    InMux I__4603 (
            .O(N__19708),
            .I(N__19697));
    Span12Mux_v I__4602 (
            .O(N__19705),
            .I(N__19694));
    Span4Mux_v I__4601 (
            .O(N__19700),
            .I(N__19691));
    LocalMux I__4600 (
            .O(N__19697),
            .I(\c0.tx2_active ));
    Odrv12 I__4599 (
            .O(N__19694),
            .I(\c0.tx2_active ));
    Odrv4 I__4598 (
            .O(N__19691),
            .I(\c0.tx2_active ));
    InMux I__4597 (
            .O(N__19684),
            .I(N__19681));
    LocalMux I__4596 (
            .O(N__19681),
            .I(\c0.N_170_0 ));
    ClkMux I__4595 (
            .O(N__19678),
            .I(N__19375));
    ClkMux I__4594 (
            .O(N__19677),
            .I(N__19375));
    ClkMux I__4593 (
            .O(N__19676),
            .I(N__19375));
    ClkMux I__4592 (
            .O(N__19675),
            .I(N__19375));
    ClkMux I__4591 (
            .O(N__19674),
            .I(N__19375));
    ClkMux I__4590 (
            .O(N__19673),
            .I(N__19375));
    ClkMux I__4589 (
            .O(N__19672),
            .I(N__19375));
    ClkMux I__4588 (
            .O(N__19671),
            .I(N__19375));
    ClkMux I__4587 (
            .O(N__19670),
            .I(N__19375));
    ClkMux I__4586 (
            .O(N__19669),
            .I(N__19375));
    ClkMux I__4585 (
            .O(N__19668),
            .I(N__19375));
    ClkMux I__4584 (
            .O(N__19667),
            .I(N__19375));
    ClkMux I__4583 (
            .O(N__19666),
            .I(N__19375));
    ClkMux I__4582 (
            .O(N__19665),
            .I(N__19375));
    ClkMux I__4581 (
            .O(N__19664),
            .I(N__19375));
    ClkMux I__4580 (
            .O(N__19663),
            .I(N__19375));
    ClkMux I__4579 (
            .O(N__19662),
            .I(N__19375));
    ClkMux I__4578 (
            .O(N__19661),
            .I(N__19375));
    ClkMux I__4577 (
            .O(N__19660),
            .I(N__19375));
    ClkMux I__4576 (
            .O(N__19659),
            .I(N__19375));
    ClkMux I__4575 (
            .O(N__19658),
            .I(N__19375));
    ClkMux I__4574 (
            .O(N__19657),
            .I(N__19375));
    ClkMux I__4573 (
            .O(N__19656),
            .I(N__19375));
    ClkMux I__4572 (
            .O(N__19655),
            .I(N__19375));
    ClkMux I__4571 (
            .O(N__19654),
            .I(N__19375));
    ClkMux I__4570 (
            .O(N__19653),
            .I(N__19375));
    ClkMux I__4569 (
            .O(N__19652),
            .I(N__19375));
    ClkMux I__4568 (
            .O(N__19651),
            .I(N__19375));
    ClkMux I__4567 (
            .O(N__19650),
            .I(N__19375));
    ClkMux I__4566 (
            .O(N__19649),
            .I(N__19375));
    ClkMux I__4565 (
            .O(N__19648),
            .I(N__19375));
    ClkMux I__4564 (
            .O(N__19647),
            .I(N__19375));
    ClkMux I__4563 (
            .O(N__19646),
            .I(N__19375));
    ClkMux I__4562 (
            .O(N__19645),
            .I(N__19375));
    ClkMux I__4561 (
            .O(N__19644),
            .I(N__19375));
    ClkMux I__4560 (
            .O(N__19643),
            .I(N__19375));
    ClkMux I__4559 (
            .O(N__19642),
            .I(N__19375));
    ClkMux I__4558 (
            .O(N__19641),
            .I(N__19375));
    ClkMux I__4557 (
            .O(N__19640),
            .I(N__19375));
    ClkMux I__4556 (
            .O(N__19639),
            .I(N__19375));
    ClkMux I__4555 (
            .O(N__19638),
            .I(N__19375));
    ClkMux I__4554 (
            .O(N__19637),
            .I(N__19375));
    ClkMux I__4553 (
            .O(N__19636),
            .I(N__19375));
    ClkMux I__4552 (
            .O(N__19635),
            .I(N__19375));
    ClkMux I__4551 (
            .O(N__19634),
            .I(N__19375));
    ClkMux I__4550 (
            .O(N__19633),
            .I(N__19375));
    ClkMux I__4549 (
            .O(N__19632),
            .I(N__19375));
    ClkMux I__4548 (
            .O(N__19631),
            .I(N__19375));
    ClkMux I__4547 (
            .O(N__19630),
            .I(N__19375));
    ClkMux I__4546 (
            .O(N__19629),
            .I(N__19375));
    ClkMux I__4545 (
            .O(N__19628),
            .I(N__19375));
    ClkMux I__4544 (
            .O(N__19627),
            .I(N__19375));
    ClkMux I__4543 (
            .O(N__19626),
            .I(N__19375));
    ClkMux I__4542 (
            .O(N__19625),
            .I(N__19375));
    ClkMux I__4541 (
            .O(N__19624),
            .I(N__19375));
    ClkMux I__4540 (
            .O(N__19623),
            .I(N__19375));
    ClkMux I__4539 (
            .O(N__19622),
            .I(N__19375));
    ClkMux I__4538 (
            .O(N__19621),
            .I(N__19375));
    ClkMux I__4537 (
            .O(N__19620),
            .I(N__19375));
    ClkMux I__4536 (
            .O(N__19619),
            .I(N__19375));
    ClkMux I__4535 (
            .O(N__19618),
            .I(N__19375));
    ClkMux I__4534 (
            .O(N__19617),
            .I(N__19375));
    ClkMux I__4533 (
            .O(N__19616),
            .I(N__19375));
    ClkMux I__4532 (
            .O(N__19615),
            .I(N__19375));
    ClkMux I__4531 (
            .O(N__19614),
            .I(N__19375));
    ClkMux I__4530 (
            .O(N__19613),
            .I(N__19375));
    ClkMux I__4529 (
            .O(N__19612),
            .I(N__19375));
    ClkMux I__4528 (
            .O(N__19611),
            .I(N__19375));
    ClkMux I__4527 (
            .O(N__19610),
            .I(N__19375));
    ClkMux I__4526 (
            .O(N__19609),
            .I(N__19375));
    ClkMux I__4525 (
            .O(N__19608),
            .I(N__19375));
    ClkMux I__4524 (
            .O(N__19607),
            .I(N__19375));
    ClkMux I__4523 (
            .O(N__19606),
            .I(N__19375));
    ClkMux I__4522 (
            .O(N__19605),
            .I(N__19375));
    ClkMux I__4521 (
            .O(N__19604),
            .I(N__19375));
    ClkMux I__4520 (
            .O(N__19603),
            .I(N__19375));
    ClkMux I__4519 (
            .O(N__19602),
            .I(N__19375));
    ClkMux I__4518 (
            .O(N__19601),
            .I(N__19375));
    ClkMux I__4517 (
            .O(N__19600),
            .I(N__19375));
    ClkMux I__4516 (
            .O(N__19599),
            .I(N__19375));
    ClkMux I__4515 (
            .O(N__19598),
            .I(N__19375));
    ClkMux I__4514 (
            .O(N__19597),
            .I(N__19375));
    ClkMux I__4513 (
            .O(N__19596),
            .I(N__19375));
    ClkMux I__4512 (
            .O(N__19595),
            .I(N__19375));
    ClkMux I__4511 (
            .O(N__19594),
            .I(N__19375));
    ClkMux I__4510 (
            .O(N__19593),
            .I(N__19375));
    ClkMux I__4509 (
            .O(N__19592),
            .I(N__19375));
    ClkMux I__4508 (
            .O(N__19591),
            .I(N__19375));
    ClkMux I__4507 (
            .O(N__19590),
            .I(N__19375));
    ClkMux I__4506 (
            .O(N__19589),
            .I(N__19375));
    ClkMux I__4505 (
            .O(N__19588),
            .I(N__19375));
    ClkMux I__4504 (
            .O(N__19587),
            .I(N__19375));
    ClkMux I__4503 (
            .O(N__19586),
            .I(N__19375));
    ClkMux I__4502 (
            .O(N__19585),
            .I(N__19375));
    ClkMux I__4501 (
            .O(N__19584),
            .I(N__19375));
    ClkMux I__4500 (
            .O(N__19583),
            .I(N__19375));
    ClkMux I__4499 (
            .O(N__19582),
            .I(N__19375));
    ClkMux I__4498 (
            .O(N__19581),
            .I(N__19375));
    ClkMux I__4497 (
            .O(N__19580),
            .I(N__19375));
    ClkMux I__4496 (
            .O(N__19579),
            .I(N__19375));
    ClkMux I__4495 (
            .O(N__19578),
            .I(N__19375));
    GlobalMux I__4494 (
            .O(N__19375),
            .I(N__19372));
    gio2CtrlBuf I__4493 (
            .O(N__19372),
            .I(CLK_c_g));
    SRMux I__4492 (
            .O(N__19369),
            .I(N__19366));
    LocalMux I__4491 (
            .O(N__19366),
            .I(N__19362));
    SRMux I__4490 (
            .O(N__19365),
            .I(N__19359));
    Span4Mux_v I__4489 (
            .O(N__19362),
            .I(N__19354));
    LocalMux I__4488 (
            .O(N__19359),
            .I(N__19354));
    Span4Mux_h I__4487 (
            .O(N__19354),
            .I(N__19350));
    InMux I__4486 (
            .O(N__19353),
            .I(N__19347));
    Odrv4 I__4485 (
            .O(N__19350),
            .I(\c0.tx2_transmit_0_sqmuxa ));
    LocalMux I__4484 (
            .O(N__19347),
            .I(\c0.tx2_transmit_0_sqmuxa ));
    InMux I__4483 (
            .O(N__19342),
            .I(N__19336));
    InMux I__4482 (
            .O(N__19341),
            .I(N__19333));
    CascadeMux I__4481 (
            .O(N__19340),
            .I(N__19330));
    InMux I__4480 (
            .O(N__19339),
            .I(N__19327));
    LocalMux I__4479 (
            .O(N__19336),
            .I(N__19323));
    LocalMux I__4478 (
            .O(N__19333),
            .I(N__19320));
    InMux I__4477 (
            .O(N__19330),
            .I(N__19317));
    LocalMux I__4476 (
            .O(N__19327),
            .I(N__19314));
    InMux I__4475 (
            .O(N__19326),
            .I(N__19311));
    Span4Mux_h I__4474 (
            .O(N__19323),
            .I(N__19308));
    Span4Mux_h I__4473 (
            .O(N__19320),
            .I(N__19305));
    LocalMux I__4472 (
            .O(N__19317),
            .I(N__19300));
    Span4Mux_h I__4471 (
            .O(N__19314),
            .I(N__19300));
    LocalMux I__4470 (
            .O(N__19311),
            .I(\c0.wait_for_transmissionZ0 ));
    Odrv4 I__4469 (
            .O(N__19308),
            .I(\c0.wait_for_transmissionZ0 ));
    Odrv4 I__4468 (
            .O(N__19305),
            .I(\c0.wait_for_transmissionZ0 ));
    Odrv4 I__4467 (
            .O(N__19300),
            .I(\c0.wait_for_transmissionZ0 ));
    InMux I__4466 (
            .O(N__19291),
            .I(N__19288));
    LocalMux I__4465 (
            .O(N__19288),
            .I(N__19284));
    InMux I__4464 (
            .O(N__19287),
            .I(N__19281));
    Span12Mux_h I__4463 (
            .O(N__19284),
            .I(N__19278));
    LocalMux I__4462 (
            .O(N__19281),
            .I(N__19275));
    Odrv12 I__4461 (
            .O(N__19278),
            .I(\c0.i12_THRU_CO ));
    Odrv12 I__4460 (
            .O(N__19275),
            .I(\c0.i12_THRU_CO ));
    IoInMux I__4459 (
            .O(N__19270),
            .I(N__19267));
    LocalMux I__4458 (
            .O(N__19267),
            .I(N__19264));
    Span12Mux_s4_h I__4457 (
            .O(N__19264),
            .I(N__19261));
    Odrv12 I__4456 (
            .O(N__19261),
            .I(\c0.data_in_frame_0__0_sqmuxa ));
    CascadeMux I__4455 (
            .O(N__19258),
            .I(N__19255));
    InMux I__4454 (
            .O(N__19255),
            .I(N__19252));
    LocalMux I__4453 (
            .O(N__19252),
            .I(\c0.tx2.N_214_0 ));
    InMux I__4452 (
            .O(N__19249),
            .I(N__19240));
    InMux I__4451 (
            .O(N__19248),
            .I(N__19240));
    InMux I__4450 (
            .O(N__19247),
            .I(N__19237));
    InMux I__4449 (
            .O(N__19246),
            .I(N__19232));
    InMux I__4448 (
            .O(N__19245),
            .I(N__19232));
    LocalMux I__4447 (
            .O(N__19240),
            .I(\c0.tx2.r_Clock_Count12_THRU_CO ));
    LocalMux I__4446 (
            .O(N__19237),
            .I(\c0.tx2.r_Clock_Count12_THRU_CO ));
    LocalMux I__4445 (
            .O(N__19232),
            .I(\c0.tx2.r_Clock_Count12_THRU_CO ));
    CascadeMux I__4444 (
            .O(N__19225),
            .I(\c0.tx2.N_17_0_cascade_ ));
    InMux I__4443 (
            .O(N__19222),
            .I(N__19215));
    InMux I__4442 (
            .O(N__19221),
            .I(N__19212));
    InMux I__4441 (
            .O(N__19220),
            .I(N__19205));
    InMux I__4440 (
            .O(N__19219),
            .I(N__19205));
    InMux I__4439 (
            .O(N__19218),
            .I(N__19205));
    LocalMux I__4438 (
            .O(N__19215),
            .I(\c0.tx2.r_SM_Main_dup_4 ));
    LocalMux I__4437 (
            .O(N__19212),
            .I(\c0.tx2.r_SM_Main_dup_4 ));
    LocalMux I__4436 (
            .O(N__19205),
            .I(\c0.tx2.r_SM_Main_dup_4 ));
    CascadeMux I__4435 (
            .O(N__19198),
            .I(N__19195));
    InMux I__4434 (
            .O(N__19195),
            .I(N__19186));
    InMux I__4433 (
            .O(N__19194),
            .I(N__19186));
    InMux I__4432 (
            .O(N__19193),
            .I(N__19183));
    InMux I__4431 (
            .O(N__19192),
            .I(N__19178));
    InMux I__4430 (
            .O(N__19191),
            .I(N__19178));
    LocalMux I__4429 (
            .O(N__19186),
            .I(\c0.tx2.r_Bit_IndexZ1Z_0 ));
    LocalMux I__4428 (
            .O(N__19183),
            .I(\c0.tx2.r_Bit_IndexZ1Z_0 ));
    LocalMux I__4427 (
            .O(N__19178),
            .I(\c0.tx2.r_Bit_IndexZ1Z_0 ));
    CascadeMux I__4426 (
            .O(N__19171),
            .I(\c0.tx2.N_212_0_cascade_ ));
    InMux I__4425 (
            .O(N__19168),
            .I(N__19161));
    InMux I__4424 (
            .O(N__19167),
            .I(N__19158));
    InMux I__4423 (
            .O(N__19166),
            .I(N__19151));
    InMux I__4422 (
            .O(N__19165),
            .I(N__19151));
    InMux I__4421 (
            .O(N__19164),
            .I(N__19151));
    LocalMux I__4420 (
            .O(N__19161),
            .I(\c0.tx2.r_SM_Main_dup_1 ));
    LocalMux I__4419 (
            .O(N__19158),
            .I(\c0.tx2.r_SM_Main_dup_1 ));
    LocalMux I__4418 (
            .O(N__19151),
            .I(\c0.tx2.r_SM_Main_dup_1 ));
    CascadeMux I__4417 (
            .O(N__19144),
            .I(\c0.tx2.N_496_cascade_ ));
    CascadeMux I__4416 (
            .O(N__19141),
            .I(N__19135));
    InMux I__4415 (
            .O(N__19140),
            .I(N__19127));
    InMux I__4414 (
            .O(N__19139),
            .I(N__19127));
    InMux I__4413 (
            .O(N__19138),
            .I(N__19122));
    InMux I__4412 (
            .O(N__19135),
            .I(N__19122));
    InMux I__4411 (
            .O(N__19134),
            .I(N__19115));
    InMux I__4410 (
            .O(N__19133),
            .I(N__19115));
    InMux I__4409 (
            .O(N__19132),
            .I(N__19115));
    LocalMux I__4408 (
            .O(N__19127),
            .I(\c0.tx2.r_SM_Main_dup_2 ));
    LocalMux I__4407 (
            .O(N__19122),
            .I(\c0.tx2.r_SM_Main_dup_2 ));
    LocalMux I__4406 (
            .O(N__19115),
            .I(\c0.tx2.r_SM_Main_dup_2 ));
    InMux I__4405 (
            .O(N__19108),
            .I(N__19100));
    InMux I__4404 (
            .O(N__19107),
            .I(N__19100));
    InMux I__4403 (
            .O(N__19106),
            .I(N__19097));
    InMux I__4402 (
            .O(N__19105),
            .I(N__19094));
    LocalMux I__4401 (
            .O(N__19100),
            .I(N__19091));
    LocalMux I__4400 (
            .O(N__19097),
            .I(N__19088));
    LocalMux I__4399 (
            .O(N__19094),
            .I(N__19085));
    Odrv12 I__4398 (
            .O(N__19091),
            .I(\c0.tx2.N_171_0 ));
    Odrv4 I__4397 (
            .O(N__19088),
            .I(\c0.tx2.N_171_0 ));
    Odrv4 I__4396 (
            .O(N__19085),
            .I(\c0.tx2.N_171_0 ));
    InMux I__4395 (
            .O(N__19078),
            .I(N__19074));
    InMux I__4394 (
            .O(N__19077),
            .I(N__19071));
    LocalMux I__4393 (
            .O(N__19074),
            .I(\c0.tx2.N_17_0 ));
    LocalMux I__4392 (
            .O(N__19071),
            .I(\c0.tx2.N_17_0 ));
    CascadeMux I__4391 (
            .O(N__19066),
            .I(N__19063));
    InMux I__4390 (
            .O(N__19063),
            .I(N__19060));
    LocalMux I__4389 (
            .O(N__19060),
            .I(\c0.tx2.N_212_0 ));
    InMux I__4388 (
            .O(N__19057),
            .I(N__19051));
    InMux I__4387 (
            .O(N__19056),
            .I(N__19051));
    LocalMux I__4386 (
            .O(N__19051),
            .I(\c0.tx2.N_493 ));
    InMux I__4385 (
            .O(N__19048),
            .I(N__19042));
    InMux I__4384 (
            .O(N__19047),
            .I(N__19039));
    InMux I__4383 (
            .O(N__19046),
            .I(N__19036));
    InMux I__4382 (
            .O(N__19045),
            .I(N__19033));
    LocalMux I__4381 (
            .O(N__19042),
            .I(\c0.tx2.r_SM_Main_dup_3 ));
    LocalMux I__4380 (
            .O(N__19039),
            .I(\c0.tx2.r_SM_Main_dup_3 ));
    LocalMux I__4379 (
            .O(N__19036),
            .I(\c0.tx2.r_SM_Main_dup_3 ));
    LocalMux I__4378 (
            .O(N__19033),
            .I(\c0.tx2.r_SM_Main_dup_3 ));
    CascadeMux I__4377 (
            .O(N__19024),
            .I(N__19021));
    InMux I__4376 (
            .O(N__19021),
            .I(N__19014));
    InMux I__4375 (
            .O(N__19020),
            .I(N__19014));
    InMux I__4374 (
            .O(N__19019),
            .I(N__19011));
    LocalMux I__4373 (
            .O(N__19014),
            .I(\c0.tx2.r_Clock_CountZ0Z_2 ));
    LocalMux I__4372 (
            .O(N__19011),
            .I(\c0.tx2.r_Clock_CountZ0Z_2 ));
    CascadeMux I__4371 (
            .O(N__19006),
            .I(N__19003));
    InMux I__4370 (
            .O(N__19003),
            .I(N__18996));
    InMux I__4369 (
            .O(N__19002),
            .I(N__18996));
    InMux I__4368 (
            .O(N__19001),
            .I(N__18993));
    LocalMux I__4367 (
            .O(N__18996),
            .I(\c0.tx2.r_Clock_CountZ0Z_1 ));
    LocalMux I__4366 (
            .O(N__18993),
            .I(\c0.tx2.r_Clock_CountZ0Z_1 ));
    CascadeMux I__4365 (
            .O(N__18988),
            .I(N__18984));
    InMux I__4364 (
            .O(N__18987),
            .I(N__18978));
    InMux I__4363 (
            .O(N__18984),
            .I(N__18978));
    InMux I__4362 (
            .O(N__18983),
            .I(N__18975));
    LocalMux I__4361 (
            .O(N__18978),
            .I(\c0.tx2.r_Clock_CountZ0Z_3 ));
    LocalMux I__4360 (
            .O(N__18975),
            .I(\c0.tx2.r_Clock_CountZ0Z_3 ));
    InMux I__4359 (
            .O(N__18970),
            .I(N__18963));
    InMux I__4358 (
            .O(N__18969),
            .I(N__18963));
    InMux I__4357 (
            .O(N__18968),
            .I(N__18960));
    LocalMux I__4356 (
            .O(N__18963),
            .I(\c0.tx2.r_Clock_CountZ0Z_0 ));
    LocalMux I__4355 (
            .O(N__18960),
            .I(\c0.tx2.r_Clock_CountZ0Z_0 ));
    InMux I__4354 (
            .O(N__18955),
            .I(N__18949));
    InMux I__4353 (
            .O(N__18954),
            .I(N__18949));
    LocalMux I__4352 (
            .O(N__18949),
            .I(N__18944));
    InMux I__4351 (
            .O(N__18948),
            .I(N__18939));
    InMux I__4350 (
            .O(N__18947),
            .I(N__18939));
    Odrv4 I__4349 (
            .O(N__18944),
            .I(\c0.tx2.N_16_0 ));
    LocalMux I__4348 (
            .O(N__18939),
            .I(\c0.tx2.N_16_0 ));
    InMux I__4347 (
            .O(N__18934),
            .I(N__18930));
    CascadeMux I__4346 (
            .O(N__18933),
            .I(N__18927));
    LocalMux I__4345 (
            .O(N__18930),
            .I(N__18924));
    InMux I__4344 (
            .O(N__18927),
            .I(N__18921));
    Odrv4 I__4343 (
            .O(N__18924),
            .I(\c0.tx2.r_Clock_Count_0_sqmuxa ));
    LocalMux I__4342 (
            .O(N__18921),
            .I(\c0.tx2.r_Clock_Count_0_sqmuxa ));
    CascadeMux I__4341 (
            .O(N__18916),
            .I(\c0.tx2.N_83_0_cascade_ ));
    CascadeMux I__4340 (
            .O(N__18913),
            .I(\c0.N_90_dup_cascade_ ));
    CascadeMux I__4339 (
            .O(N__18910),
            .I(\c0.tx2.i97_mux_cascade_ ));
    InMux I__4338 (
            .O(N__18907),
            .I(N__18904));
    LocalMux I__4337 (
            .O(N__18904),
            .I(\c0.tx2.r_SM_Main_illegal_0 ));
    InMux I__4336 (
            .O(N__18901),
            .I(N__18898));
    LocalMux I__4335 (
            .O(N__18898),
            .I(N__18895));
    Span4Mux_h I__4334 (
            .O(N__18895),
            .I(N__18891));
    InMux I__4333 (
            .O(N__18894),
            .I(N__18888));
    Odrv4 I__4332 (
            .O(N__18891),
            .I(\c0.d_4_0 ));
    LocalMux I__4331 (
            .O(N__18888),
            .I(\c0.d_4_0 ));
    InMux I__4330 (
            .O(N__18883),
            .I(N__18880));
    LocalMux I__4329 (
            .O(N__18880),
            .I(N__18877));
    Span4Mux_v I__4328 (
            .O(N__18877),
            .I(N__18873));
    InMux I__4327 (
            .O(N__18876),
            .I(N__18870));
    Sp12to4 I__4326 (
            .O(N__18873),
            .I(N__18864));
    LocalMux I__4325 (
            .O(N__18870),
            .I(N__18864));
    InMux I__4324 (
            .O(N__18869),
            .I(N__18861));
    Odrv12 I__4323 (
            .O(N__18864),
            .I(\c0.d_4_8 ));
    LocalMux I__4322 (
            .O(N__18861),
            .I(\c0.d_4_8 ));
    InMux I__4321 (
            .O(N__18856),
            .I(N__18853));
    LocalMux I__4320 (
            .O(N__18853),
            .I(N__18850));
    Span4Mux_h I__4319 (
            .O(N__18850),
            .I(N__18844));
    InMux I__4318 (
            .O(N__18849),
            .I(N__18839));
    InMux I__4317 (
            .O(N__18848),
            .I(N__18839));
    InMux I__4316 (
            .O(N__18847),
            .I(N__18836));
    Odrv4 I__4315 (
            .O(N__18844),
            .I(\c0.d_4_16 ));
    LocalMux I__4314 (
            .O(N__18839),
            .I(\c0.d_4_16 ));
    LocalMux I__4313 (
            .O(N__18836),
            .I(\c0.d_4_16 ));
    CascadeMux I__4312 (
            .O(N__18829),
            .I(N__18826));
    InMux I__4311 (
            .O(N__18826),
            .I(N__18823));
    LocalMux I__4310 (
            .O(N__18823),
            .I(N__18820));
    Span4Mux_v I__4309 (
            .O(N__18820),
            .I(N__18815));
    InMux I__4308 (
            .O(N__18819),
            .I(N__18812));
    InMux I__4307 (
            .O(N__18818),
            .I(N__18809));
    Span4Mux_h I__4306 (
            .O(N__18815),
            .I(N__18804));
    LocalMux I__4305 (
            .O(N__18812),
            .I(N__18804));
    LocalMux I__4304 (
            .O(N__18809),
            .I(\c0.d_4_24 ));
    Odrv4 I__4303 (
            .O(N__18804),
            .I(\c0.d_4_24 ));
    InMux I__4302 (
            .O(N__18799),
            .I(N__18792));
    InMux I__4301 (
            .O(N__18798),
            .I(N__18788));
    InMux I__4300 (
            .O(N__18797),
            .I(N__18785));
    InMux I__4299 (
            .O(N__18796),
            .I(N__18779));
    InMux I__4298 (
            .O(N__18795),
            .I(N__18779));
    LocalMux I__4297 (
            .O(N__18792),
            .I(N__18776));
    InMux I__4296 (
            .O(N__18791),
            .I(N__18773));
    LocalMux I__4295 (
            .O(N__18788),
            .I(N__18768));
    LocalMux I__4294 (
            .O(N__18785),
            .I(N__18768));
    InMux I__4293 (
            .O(N__18784),
            .I(N__18765));
    LocalMux I__4292 (
            .O(N__18779),
            .I(N__18759));
    Span4Mux_h I__4291 (
            .O(N__18776),
            .I(N__18754));
    LocalMux I__4290 (
            .O(N__18773),
            .I(N__18754));
    Span4Mux_v I__4289 (
            .O(N__18768),
            .I(N__18749));
    LocalMux I__4288 (
            .O(N__18765),
            .I(N__18749));
    InMux I__4287 (
            .O(N__18764),
            .I(N__18746));
    InMux I__4286 (
            .O(N__18763),
            .I(N__18741));
    InMux I__4285 (
            .O(N__18762),
            .I(N__18741));
    Odrv12 I__4284 (
            .O(N__18759),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    Odrv4 I__4283 (
            .O(N__18754),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    Odrv4 I__4282 (
            .O(N__18749),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    LocalMux I__4281 (
            .O(N__18746),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    LocalMux I__4280 (
            .O(N__18741),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    InMux I__4279 (
            .O(N__18730),
            .I(N__18727));
    LocalMux I__4278 (
            .O(N__18727),
            .I(\c0.tx2_data_RNO_3Z0Z_0 ));
    CascadeMux I__4277 (
            .O(N__18724),
            .I(\c0.tx2_data_RNO_4Z0Z_0_cascade_ ));
    InMux I__4276 (
            .O(N__18721),
            .I(N__18705));
    InMux I__4275 (
            .O(N__18720),
            .I(N__18700));
    InMux I__4274 (
            .O(N__18719),
            .I(N__18700));
    InMux I__4273 (
            .O(N__18718),
            .I(N__18697));
    InMux I__4272 (
            .O(N__18717),
            .I(N__18690));
    InMux I__4271 (
            .O(N__18716),
            .I(N__18690));
    InMux I__4270 (
            .O(N__18715),
            .I(N__18690));
    InMux I__4269 (
            .O(N__18714),
            .I(N__18687));
    InMux I__4268 (
            .O(N__18713),
            .I(N__18684));
    InMux I__4267 (
            .O(N__18712),
            .I(N__18681));
    InMux I__4266 (
            .O(N__18711),
            .I(N__18674));
    InMux I__4265 (
            .O(N__18710),
            .I(N__18674));
    InMux I__4264 (
            .O(N__18709),
            .I(N__18674));
    InMux I__4263 (
            .O(N__18708),
            .I(N__18671));
    LocalMux I__4262 (
            .O(N__18705),
            .I(N__18666));
    LocalMux I__4261 (
            .O(N__18700),
            .I(N__18666));
    LocalMux I__4260 (
            .O(N__18697),
            .I(N__18663));
    LocalMux I__4259 (
            .O(N__18690),
            .I(N__18658));
    LocalMux I__4258 (
            .O(N__18687),
            .I(N__18658));
    LocalMux I__4257 (
            .O(N__18684),
            .I(N__18649));
    LocalMux I__4256 (
            .O(N__18681),
            .I(N__18649));
    LocalMux I__4255 (
            .O(N__18674),
            .I(N__18646));
    LocalMux I__4254 (
            .O(N__18671),
            .I(N__18641));
    Span4Mux_v I__4253 (
            .O(N__18666),
            .I(N__18641));
    Span4Mux_v I__4252 (
            .O(N__18663),
            .I(N__18636));
    Span4Mux_h I__4251 (
            .O(N__18658),
            .I(N__18636));
    InMux I__4250 (
            .O(N__18657),
            .I(N__18633));
    InMux I__4249 (
            .O(N__18656),
            .I(N__18626));
    InMux I__4248 (
            .O(N__18655),
            .I(N__18626));
    InMux I__4247 (
            .O(N__18654),
            .I(N__18626));
    Odrv4 I__4246 (
            .O(N__18649),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    Odrv12 I__4245 (
            .O(N__18646),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    Odrv4 I__4244 (
            .O(N__18641),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    Odrv4 I__4243 (
            .O(N__18636),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    LocalMux I__4242 (
            .O(N__18633),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    LocalMux I__4241 (
            .O(N__18626),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    InMux I__4240 (
            .O(N__18613),
            .I(N__18610));
    LocalMux I__4239 (
            .O(N__18610),
            .I(N__18607));
    Odrv12 I__4238 (
            .O(N__18607),
            .I(\c0.tx2_data_RNO_1Z0Z_0 ));
    CascadeMux I__4237 (
            .O(N__18604),
            .I(\c0.m146_ns_1_cascade_ ));
    InMux I__4236 (
            .O(N__18601),
            .I(N__18598));
    LocalMux I__4235 (
            .O(N__18598),
            .I(\c0.tx2.r_Tx_DataZ0Z_0 ));
    CascadeMux I__4234 (
            .O(N__18595),
            .I(N__18583));
    CascadeMux I__4233 (
            .O(N__18594),
            .I(N__18579));
    CascadeMux I__4232 (
            .O(N__18593),
            .I(N__18573));
    InMux I__4231 (
            .O(N__18592),
            .I(N__18562));
    InMux I__4230 (
            .O(N__18591),
            .I(N__18555));
    InMux I__4229 (
            .O(N__18590),
            .I(N__18555));
    InMux I__4228 (
            .O(N__18589),
            .I(N__18555));
    InMux I__4227 (
            .O(N__18588),
            .I(N__18550));
    InMux I__4226 (
            .O(N__18587),
            .I(N__18550));
    InMux I__4225 (
            .O(N__18586),
            .I(N__18543));
    InMux I__4224 (
            .O(N__18583),
            .I(N__18543));
    InMux I__4223 (
            .O(N__18582),
            .I(N__18543));
    InMux I__4222 (
            .O(N__18579),
            .I(N__18536));
    InMux I__4221 (
            .O(N__18578),
            .I(N__18536));
    InMux I__4220 (
            .O(N__18577),
            .I(N__18536));
    InMux I__4219 (
            .O(N__18576),
            .I(N__18533));
    InMux I__4218 (
            .O(N__18573),
            .I(N__18528));
    InMux I__4217 (
            .O(N__18572),
            .I(N__18521));
    InMux I__4216 (
            .O(N__18571),
            .I(N__18521));
    CascadeMux I__4215 (
            .O(N__18570),
            .I(N__18515));
    InMux I__4214 (
            .O(N__18569),
            .I(N__18510));
    InMux I__4213 (
            .O(N__18568),
            .I(N__18501));
    InMux I__4212 (
            .O(N__18567),
            .I(N__18501));
    InMux I__4211 (
            .O(N__18566),
            .I(N__18501));
    InMux I__4210 (
            .O(N__18565),
            .I(N__18501));
    LocalMux I__4209 (
            .O(N__18562),
            .I(N__18496));
    LocalMux I__4208 (
            .O(N__18555),
            .I(N__18496));
    LocalMux I__4207 (
            .O(N__18550),
            .I(N__18493));
    LocalMux I__4206 (
            .O(N__18543),
            .I(N__18490));
    LocalMux I__4205 (
            .O(N__18536),
            .I(N__18485));
    LocalMux I__4204 (
            .O(N__18533),
            .I(N__18485));
    InMux I__4203 (
            .O(N__18532),
            .I(N__18479));
    InMux I__4202 (
            .O(N__18531),
            .I(N__18476));
    LocalMux I__4201 (
            .O(N__18528),
            .I(N__18473));
    InMux I__4200 (
            .O(N__18527),
            .I(N__18468));
    InMux I__4199 (
            .O(N__18526),
            .I(N__18468));
    LocalMux I__4198 (
            .O(N__18521),
            .I(N__18465));
    InMux I__4197 (
            .O(N__18520),
            .I(N__18458));
    InMux I__4196 (
            .O(N__18519),
            .I(N__18458));
    InMux I__4195 (
            .O(N__18518),
            .I(N__18458));
    InMux I__4194 (
            .O(N__18515),
            .I(N__18453));
    InMux I__4193 (
            .O(N__18514),
            .I(N__18453));
    InMux I__4192 (
            .O(N__18513),
            .I(N__18450));
    LocalMux I__4191 (
            .O(N__18510),
            .I(N__18443));
    LocalMux I__4190 (
            .O(N__18501),
            .I(N__18443));
    Span4Mux_h I__4189 (
            .O(N__18496),
            .I(N__18443));
    Span4Mux_h I__4188 (
            .O(N__18493),
            .I(N__18436));
    Span4Mux_v I__4187 (
            .O(N__18490),
            .I(N__18436));
    Span4Mux_h I__4186 (
            .O(N__18485),
            .I(N__18436));
    InMux I__4185 (
            .O(N__18484),
            .I(N__18429));
    InMux I__4184 (
            .O(N__18483),
            .I(N__18429));
    InMux I__4183 (
            .O(N__18482),
            .I(N__18429));
    LocalMux I__4182 (
            .O(N__18479),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4181 (
            .O(N__18476),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    Odrv12 I__4180 (
            .O(N__18473),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4179 (
            .O(N__18468),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    Odrv12 I__4178 (
            .O(N__18465),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4177 (
            .O(N__18458),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4176 (
            .O(N__18453),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4175 (
            .O(N__18450),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    Odrv4 I__4174 (
            .O(N__18443),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    Odrv4 I__4173 (
            .O(N__18436),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4172 (
            .O(N__18429),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    InMux I__4171 (
            .O(N__18406),
            .I(N__18403));
    LocalMux I__4170 (
            .O(N__18403),
            .I(N__18396));
    InMux I__4169 (
            .O(N__18402),
            .I(N__18393));
    InMux I__4168 (
            .O(N__18401),
            .I(N__18390));
    InMux I__4167 (
            .O(N__18400),
            .I(N__18385));
    InMux I__4166 (
            .O(N__18399),
            .I(N__18385));
    Odrv4 I__4165 (
            .O(N__18396),
            .I(\c0.d_4_32 ));
    LocalMux I__4164 (
            .O(N__18393),
            .I(\c0.d_4_32 ));
    LocalMux I__4163 (
            .O(N__18390),
            .I(\c0.d_4_32 ));
    LocalMux I__4162 (
            .O(N__18385),
            .I(\c0.d_4_32 ));
    CascadeMux I__4161 (
            .O(N__18376),
            .I(N__18366));
    CascadeMux I__4160 (
            .O(N__18375),
            .I(N__18362));
    CascadeMux I__4159 (
            .O(N__18374),
            .I(N__18358));
    CascadeMux I__4158 (
            .O(N__18373),
            .I(N__18349));
    CascadeMux I__4157 (
            .O(N__18372),
            .I(N__18344));
    CascadeMux I__4156 (
            .O(N__18371),
            .I(N__18341));
    InMux I__4155 (
            .O(N__18370),
            .I(N__18334));
    InMux I__4154 (
            .O(N__18369),
            .I(N__18334));
    InMux I__4153 (
            .O(N__18366),
            .I(N__18334));
    InMux I__4152 (
            .O(N__18365),
            .I(N__18324));
    InMux I__4151 (
            .O(N__18362),
            .I(N__18324));
    InMux I__4150 (
            .O(N__18361),
            .I(N__18319));
    InMux I__4149 (
            .O(N__18358),
            .I(N__18319));
    InMux I__4148 (
            .O(N__18357),
            .I(N__18312));
    InMux I__4147 (
            .O(N__18356),
            .I(N__18312));
    InMux I__4146 (
            .O(N__18355),
            .I(N__18312));
    InMux I__4145 (
            .O(N__18354),
            .I(N__18309));
    CascadeMux I__4144 (
            .O(N__18353),
            .I(N__18306));
    CascadeMux I__4143 (
            .O(N__18352),
            .I(N__18298));
    InMux I__4142 (
            .O(N__18349),
            .I(N__18293));
    InMux I__4141 (
            .O(N__18348),
            .I(N__18293));
    InMux I__4140 (
            .O(N__18347),
            .I(N__18286));
    InMux I__4139 (
            .O(N__18344),
            .I(N__18286));
    InMux I__4138 (
            .O(N__18341),
            .I(N__18286));
    LocalMux I__4137 (
            .O(N__18334),
            .I(N__18283));
    CascadeMux I__4136 (
            .O(N__18333),
            .I(N__18279));
    CascadeMux I__4135 (
            .O(N__18332),
            .I(N__18275));
    CascadeMux I__4134 (
            .O(N__18331),
            .I(N__18271));
    CascadeMux I__4133 (
            .O(N__18330),
            .I(N__18268));
    CascadeMux I__4132 (
            .O(N__18329),
            .I(N__18264));
    LocalMux I__4131 (
            .O(N__18324),
            .I(N__18261));
    LocalMux I__4130 (
            .O(N__18319),
            .I(N__18258));
    LocalMux I__4129 (
            .O(N__18312),
            .I(N__18253));
    LocalMux I__4128 (
            .O(N__18309),
            .I(N__18253));
    InMux I__4127 (
            .O(N__18306),
            .I(N__18248));
    InMux I__4126 (
            .O(N__18305),
            .I(N__18248));
    InMux I__4125 (
            .O(N__18304),
            .I(N__18237));
    InMux I__4124 (
            .O(N__18303),
            .I(N__18237));
    InMux I__4123 (
            .O(N__18302),
            .I(N__18237));
    InMux I__4122 (
            .O(N__18301),
            .I(N__18237));
    InMux I__4121 (
            .O(N__18298),
            .I(N__18237));
    LocalMux I__4120 (
            .O(N__18293),
            .I(N__18232));
    LocalMux I__4119 (
            .O(N__18286),
            .I(N__18232));
    Span4Mux_h I__4118 (
            .O(N__18283),
            .I(N__18229));
    InMux I__4117 (
            .O(N__18282),
            .I(N__18224));
    InMux I__4116 (
            .O(N__18279),
            .I(N__18224));
    InMux I__4115 (
            .O(N__18278),
            .I(N__18215));
    InMux I__4114 (
            .O(N__18275),
            .I(N__18215));
    InMux I__4113 (
            .O(N__18274),
            .I(N__18215));
    InMux I__4112 (
            .O(N__18271),
            .I(N__18215));
    InMux I__4111 (
            .O(N__18268),
            .I(N__18208));
    InMux I__4110 (
            .O(N__18267),
            .I(N__18208));
    InMux I__4109 (
            .O(N__18264),
            .I(N__18208));
    Span4Mux_v I__4108 (
            .O(N__18261),
            .I(N__18199));
    Span4Mux_h I__4107 (
            .O(N__18258),
            .I(N__18199));
    Span4Mux_v I__4106 (
            .O(N__18253),
            .I(N__18199));
    LocalMux I__4105 (
            .O(N__18248),
            .I(N__18199));
    LocalMux I__4104 (
            .O(N__18237),
            .I(N__18194));
    Span4Mux_h I__4103 (
            .O(N__18232),
            .I(N__18194));
    Odrv4 I__4102 (
            .O(N__18229),
            .I(\c0.N_204_mux ));
    LocalMux I__4101 (
            .O(N__18224),
            .I(\c0.N_204_mux ));
    LocalMux I__4100 (
            .O(N__18215),
            .I(\c0.N_204_mux ));
    LocalMux I__4099 (
            .O(N__18208),
            .I(\c0.N_204_mux ));
    Odrv4 I__4098 (
            .O(N__18199),
            .I(\c0.N_204_mux ));
    Odrv4 I__4097 (
            .O(N__18194),
            .I(\c0.N_204_mux ));
    InMux I__4096 (
            .O(N__18181),
            .I(N__18178));
    LocalMux I__4095 (
            .O(N__18178),
            .I(N__18175));
    Span4Mux_h I__4094 (
            .O(N__18175),
            .I(N__18170));
    InMux I__4093 (
            .O(N__18174),
            .I(N__18167));
    InMux I__4092 (
            .O(N__18173),
            .I(N__18164));
    Odrv4 I__4091 (
            .O(N__18170),
            .I(\c0.d_4_40 ));
    LocalMux I__4090 (
            .O(N__18167),
            .I(\c0.d_4_40 ));
    LocalMux I__4089 (
            .O(N__18164),
            .I(\c0.d_4_40 ));
    InMux I__4088 (
            .O(N__18157),
            .I(N__18154));
    LocalMux I__4087 (
            .O(N__18154),
            .I(\c0.tx2_data_RNO_0Z0Z_0 ));
    InMux I__4086 (
            .O(N__18151),
            .I(\c0.tx2.un1_r_Clock_Count_cry_0 ));
    InMux I__4085 (
            .O(N__18148),
            .I(\c0.tx2.un1_r_Clock_Count_cry_1 ));
    InMux I__4084 (
            .O(N__18145),
            .I(\c0.tx2.un1_r_Clock_Count_cry_2 ));
    InMux I__4083 (
            .O(N__18142),
            .I(N__18138));
    InMux I__4082 (
            .O(N__18141),
            .I(N__18135));
    LocalMux I__4081 (
            .O(N__18138),
            .I(N__18132));
    LocalMux I__4080 (
            .O(N__18135),
            .I(N__18129));
    Odrv4 I__4079 (
            .O(N__18132),
            .I(\c0.N_164_0 ));
    Odrv4 I__4078 (
            .O(N__18129),
            .I(\c0.N_164_0 ));
    InMux I__4077 (
            .O(N__18124),
            .I(N__18121));
    LocalMux I__4076 (
            .O(N__18121),
            .I(N__18118));
    Span4Mux_h I__4075 (
            .O(N__18118),
            .I(N__18114));
    InMux I__4074 (
            .O(N__18117),
            .I(N__18111));
    Odrv4 I__4073 (
            .O(N__18114),
            .I(\c0.d_4_22 ));
    LocalMux I__4072 (
            .O(N__18111),
            .I(\c0.d_4_22 ));
    CascadeMux I__4071 (
            .O(N__18106),
            .I(N__18103));
    InMux I__4070 (
            .O(N__18103),
            .I(N__18100));
    LocalMux I__4069 (
            .O(N__18100),
            .I(N__18097));
    Span4Mux_v I__4068 (
            .O(N__18097),
            .I(N__18091));
    InMux I__4067 (
            .O(N__18096),
            .I(N__18088));
    InMux I__4066 (
            .O(N__18095),
            .I(N__18085));
    InMux I__4065 (
            .O(N__18094),
            .I(N__18082));
    Odrv4 I__4064 (
            .O(N__18091),
            .I(\c0.d_4_30 ));
    LocalMux I__4063 (
            .O(N__18088),
            .I(\c0.d_4_30 ));
    LocalMux I__4062 (
            .O(N__18085),
            .I(\c0.d_4_30 ));
    LocalMux I__4061 (
            .O(N__18082),
            .I(\c0.d_4_30 ));
    CascadeMux I__4060 (
            .O(N__18073),
            .I(N__18070));
    InMux I__4059 (
            .O(N__18070),
            .I(N__18067));
    LocalMux I__4058 (
            .O(N__18067),
            .I(N__18064));
    Odrv4 I__4057 (
            .O(N__18064),
            .I(\c0.tx2_data_RNO_4Z0Z_6 ));
    InMux I__4056 (
            .O(N__18061),
            .I(N__18058));
    LocalMux I__4055 (
            .O(N__18058),
            .I(N__18055));
    Span12Mux_h I__4054 (
            .O(N__18055),
            .I(N__18051));
    InMux I__4053 (
            .O(N__18054),
            .I(N__18048));
    Odrv12 I__4052 (
            .O(N__18051),
            .I(\c0.d_4_4 ));
    LocalMux I__4051 (
            .O(N__18048),
            .I(\c0.d_4_4 ));
    InMux I__4050 (
            .O(N__18043),
            .I(N__18040));
    LocalMux I__4049 (
            .O(N__18040),
            .I(N__18037));
    Span4Mux_h I__4048 (
            .O(N__18037),
            .I(N__18031));
    InMux I__4047 (
            .O(N__18036),
            .I(N__18026));
    InMux I__4046 (
            .O(N__18035),
            .I(N__18026));
    InMux I__4045 (
            .O(N__18034),
            .I(N__18023));
    Odrv4 I__4044 (
            .O(N__18031),
            .I(\c0.d_4_12 ));
    LocalMux I__4043 (
            .O(N__18026),
            .I(\c0.d_4_12 ));
    LocalMux I__4042 (
            .O(N__18023),
            .I(\c0.d_4_12 ));
    CascadeMux I__4041 (
            .O(N__18016),
            .I(N__18013));
    InMux I__4040 (
            .O(N__18013),
            .I(N__18010));
    LocalMux I__4039 (
            .O(N__18010),
            .I(N__18007));
    Odrv4 I__4038 (
            .O(N__18007),
            .I(\c0.tx2_data_RNO_3Z0Z_4 ));
    CascadeMux I__4037 (
            .O(N__18004),
            .I(N__18000));
    InMux I__4036 (
            .O(N__18003),
            .I(N__17997));
    InMux I__4035 (
            .O(N__18000),
            .I(N__17994));
    LocalMux I__4034 (
            .O(N__17997),
            .I(N__17988));
    LocalMux I__4033 (
            .O(N__17994),
            .I(N__17988));
    InMux I__4032 (
            .O(N__17993),
            .I(N__17985));
    Span4Mux_v I__4031 (
            .O(N__17988),
            .I(N__17981));
    LocalMux I__4030 (
            .O(N__17985),
            .I(N__17978));
    InMux I__4029 (
            .O(N__17984),
            .I(N__17975));
    Odrv4 I__4028 (
            .O(N__17981),
            .I(\c0.d_4_28 ));
    Odrv12 I__4027 (
            .O(N__17978),
            .I(\c0.d_4_28 ));
    LocalMux I__4026 (
            .O(N__17975),
            .I(\c0.d_4_28 ));
    InMux I__4025 (
            .O(N__17968),
            .I(N__17965));
    LocalMux I__4024 (
            .O(N__17965),
            .I(N__17961));
    InMux I__4023 (
            .O(N__17964),
            .I(N__17957));
    Span4Mux_h I__4022 (
            .O(N__17961),
            .I(N__17954));
    InMux I__4021 (
            .O(N__17960),
            .I(N__17951));
    LocalMux I__4020 (
            .O(N__17957),
            .I(N__17948));
    Odrv4 I__4019 (
            .O(N__17954),
            .I(\c0.d_4_20 ));
    LocalMux I__4018 (
            .O(N__17951),
            .I(\c0.d_4_20 ));
    Odrv4 I__4017 (
            .O(N__17948),
            .I(\c0.d_4_20 ));
    InMux I__4016 (
            .O(N__17941),
            .I(N__17938));
    LocalMux I__4015 (
            .O(N__17938),
            .I(N__17935));
    Span4Mux_v I__4014 (
            .O(N__17935),
            .I(N__17932));
    Odrv4 I__4013 (
            .O(N__17932),
            .I(\c0.tx2_data_RNO_4Z0Z_4 ));
    InMux I__4012 (
            .O(N__17929),
            .I(N__17926));
    LocalMux I__4011 (
            .O(N__17926),
            .I(N__17923));
    Span4Mux_h I__4010 (
            .O(N__17923),
            .I(N__17919));
    InMux I__4009 (
            .O(N__17922),
            .I(N__17916));
    Odrv4 I__4008 (
            .O(N__17919),
            .I(\c0.d_4_13 ));
    LocalMux I__4007 (
            .O(N__17916),
            .I(\c0.d_4_13 ));
    CascadeMux I__4006 (
            .O(N__17911),
            .I(N__17908));
    InMux I__4005 (
            .O(N__17908),
            .I(N__17905));
    LocalMux I__4004 (
            .O(N__17905),
            .I(N__17901));
    InMux I__4003 (
            .O(N__17904),
            .I(N__17897));
    Span4Mux_h I__4002 (
            .O(N__17901),
            .I(N__17894));
    InMux I__4001 (
            .O(N__17900),
            .I(N__17891));
    LocalMux I__4000 (
            .O(N__17897),
            .I(N__17888));
    Odrv4 I__3999 (
            .O(N__17894),
            .I(\c0.d_4_5 ));
    LocalMux I__3998 (
            .O(N__17891),
            .I(\c0.d_4_5 ));
    Odrv12 I__3997 (
            .O(N__17888),
            .I(\c0.d_4_5 ));
    InMux I__3996 (
            .O(N__17881),
            .I(N__17878));
    LocalMux I__3995 (
            .O(N__17878),
            .I(\c0.tx2_data_RNO_3Z0Z_5 ));
    InMux I__3994 (
            .O(N__17875),
            .I(N__17871));
    InMux I__3993 (
            .O(N__17874),
            .I(N__17868));
    LocalMux I__3992 (
            .O(N__17871),
            .I(\c0.byte_transmit_counter2Z0Z_7 ));
    LocalMux I__3991 (
            .O(N__17868),
            .I(\c0.byte_transmit_counter2Z0Z_7 ));
    InMux I__3990 (
            .O(N__17863),
            .I(N__17859));
    InMux I__3989 (
            .O(N__17862),
            .I(N__17856));
    LocalMux I__3988 (
            .O(N__17859),
            .I(\c0.byte_transmit_counter2Z0Z_3 ));
    LocalMux I__3987 (
            .O(N__17856),
            .I(\c0.byte_transmit_counter2Z0Z_3 ));
    InMux I__3986 (
            .O(N__17851),
            .I(N__17847));
    InMux I__3985 (
            .O(N__17850),
            .I(N__17844));
    LocalMux I__3984 (
            .O(N__17847),
            .I(\c0.byte_transmit_counter2Z0Z_6 ));
    LocalMux I__3983 (
            .O(N__17844),
            .I(\c0.byte_transmit_counter2Z0Z_6 ));
    InMux I__3982 (
            .O(N__17839),
            .I(N__17835));
    InMux I__3981 (
            .O(N__17838),
            .I(N__17832));
    LocalMux I__3980 (
            .O(N__17835),
            .I(\c0.byte_transmit_counter2Z0Z_5 ));
    LocalMux I__3979 (
            .O(N__17832),
            .I(\c0.byte_transmit_counter2Z0Z_5 ));
    CascadeMux I__3978 (
            .O(N__17827),
            .I(\c0.m45_0_0_cascade_ ));
    InMux I__3977 (
            .O(N__17824),
            .I(N__17820));
    InMux I__3976 (
            .O(N__17823),
            .I(N__17817));
    LocalMux I__3975 (
            .O(N__17820),
            .I(\c0.byte_transmit_counter2Z0Z_4 ));
    LocalMux I__3974 (
            .O(N__17817),
            .I(\c0.byte_transmit_counter2Z0Z_4 ));
    CascadeMux I__3973 (
            .O(N__17812),
            .I(\c0.N_204_mux_cascade_ ));
    InMux I__3972 (
            .O(N__17809),
            .I(N__17806));
    LocalMux I__3971 (
            .O(N__17806),
            .I(N__17802));
    InMux I__3970 (
            .O(N__17805),
            .I(N__17799));
    Span4Mux_h I__3969 (
            .O(N__17802),
            .I(N__17796));
    LocalMux I__3968 (
            .O(N__17799),
            .I(\c0.N_215_mux ));
    Odrv4 I__3967 (
            .O(N__17796),
            .I(\c0.N_215_mux ));
    CascadeMux I__3966 (
            .O(N__17791),
            .I(N__17787));
    InMux I__3965 (
            .O(N__17790),
            .I(N__17784));
    InMux I__3964 (
            .O(N__17787),
            .I(N__17781));
    LocalMux I__3963 (
            .O(N__17784),
            .I(N__17776));
    LocalMux I__3962 (
            .O(N__17781),
            .I(N__17776));
    Span4Mux_v I__3961 (
            .O(N__17776),
            .I(N__17772));
    InMux I__3960 (
            .O(N__17775),
            .I(N__17769));
    Span4Mux_h I__3959 (
            .O(N__17772),
            .I(N__17766));
    LocalMux I__3958 (
            .O(N__17769),
            .I(\c0.data_in_7_Z0Z_2 ));
    Odrv4 I__3957 (
            .O(N__17766),
            .I(\c0.data_in_7_Z0Z_2 ));
    InMux I__3956 (
            .O(N__17761),
            .I(N__17758));
    LocalMux I__3955 (
            .O(N__17758),
            .I(N__17754));
    InMux I__3954 (
            .O(N__17757),
            .I(N__17751));
    Span4Mux_h I__3953 (
            .O(N__17754),
            .I(N__17746));
    LocalMux I__3952 (
            .O(N__17751),
            .I(N__17746));
    Span4Mux_h I__3951 (
            .O(N__17746),
            .I(N__17742));
    InMux I__3950 (
            .O(N__17745),
            .I(N__17739));
    Odrv4 I__3949 (
            .O(N__17742),
            .I(\c0.data_in_6_Z0Z_2 ));
    LocalMux I__3948 (
            .O(N__17739),
            .I(\c0.data_in_6_Z0Z_2 ));
    CascadeMux I__3947 (
            .O(N__17734),
            .I(N__17731));
    InMux I__3946 (
            .O(N__17731),
            .I(N__17728));
    LocalMux I__3945 (
            .O(N__17728),
            .I(N__17712));
    CEMux I__3944 (
            .O(N__17727),
            .I(N__17683));
    CEMux I__3943 (
            .O(N__17726),
            .I(N__17683));
    CEMux I__3942 (
            .O(N__17725),
            .I(N__17683));
    CEMux I__3941 (
            .O(N__17724),
            .I(N__17683));
    CEMux I__3940 (
            .O(N__17723),
            .I(N__17683));
    CEMux I__3939 (
            .O(N__17722),
            .I(N__17683));
    CEMux I__3938 (
            .O(N__17721),
            .I(N__17683));
    CEMux I__3937 (
            .O(N__17720),
            .I(N__17683));
    CEMux I__3936 (
            .O(N__17719),
            .I(N__17683));
    CEMux I__3935 (
            .O(N__17718),
            .I(N__17683));
    CEMux I__3934 (
            .O(N__17717),
            .I(N__17683));
    CEMux I__3933 (
            .O(N__17716),
            .I(N__17683));
    CEMux I__3932 (
            .O(N__17715),
            .I(N__17683));
    Glb2LocalMux I__3931 (
            .O(N__17712),
            .I(N__17683));
    GlobalMux I__3930 (
            .O(N__17683),
            .I(N__17680));
    gio2CtrlBuf I__3929 (
            .O(N__17680),
            .I(\c0.rx_data_ready_g ));
    InMux I__3928 (
            .O(N__17677),
            .I(N__17673));
    InMux I__3927 (
            .O(N__17676),
            .I(N__17670));
    LocalMux I__3926 (
            .O(N__17673),
            .I(N__17667));
    LocalMux I__3925 (
            .O(N__17670),
            .I(N__17664));
    Span4Mux_v I__3924 (
            .O(N__17667),
            .I(N__17659));
    Span4Mux_v I__3923 (
            .O(N__17664),
            .I(N__17659));
    Odrv4 I__3922 (
            .O(N__17659),
            .I(\c0.d_4_45 ));
    CascadeMux I__3921 (
            .O(N__17656),
            .I(N__17653));
    InMux I__3920 (
            .O(N__17653),
            .I(N__17650));
    LocalMux I__3919 (
            .O(N__17650),
            .I(N__17644));
    CascadeMux I__3918 (
            .O(N__17649),
            .I(N__17641));
    InMux I__3917 (
            .O(N__17648),
            .I(N__17636));
    InMux I__3916 (
            .O(N__17647),
            .I(N__17636));
    Span4Mux_h I__3915 (
            .O(N__17644),
            .I(N__17633));
    InMux I__3914 (
            .O(N__17641),
            .I(N__17630));
    LocalMux I__3913 (
            .O(N__17636),
            .I(N__17627));
    Odrv4 I__3912 (
            .O(N__17633),
            .I(\c0.d_4_37 ));
    LocalMux I__3911 (
            .O(N__17630),
            .I(\c0.d_4_37 ));
    Odrv4 I__3910 (
            .O(N__17627),
            .I(\c0.d_4_37 ));
    InMux I__3909 (
            .O(N__17620),
            .I(N__17613));
    InMux I__3908 (
            .O(N__17619),
            .I(N__17613));
    InMux I__3907 (
            .O(N__17618),
            .I(N__17610));
    LocalMux I__3906 (
            .O(N__17613),
            .I(N__17607));
    LocalMux I__3905 (
            .O(N__17610),
            .I(N__17603));
    Span4Mux_v I__3904 (
            .O(N__17607),
            .I(N__17600));
    InMux I__3903 (
            .O(N__17606),
            .I(N__17597));
    Odrv12 I__3902 (
            .O(N__17603),
            .I(\c0.d_4_29 ));
    Odrv4 I__3901 (
            .O(N__17600),
            .I(\c0.d_4_29 ));
    LocalMux I__3900 (
            .O(N__17597),
            .I(\c0.d_4_29 ));
    InMux I__3899 (
            .O(N__17590),
            .I(N__17587));
    LocalMux I__3898 (
            .O(N__17587),
            .I(N__17584));
    Span4Mux_v I__3897 (
            .O(N__17584),
            .I(N__17579));
    InMux I__3896 (
            .O(N__17583),
            .I(N__17576));
    InMux I__3895 (
            .O(N__17582),
            .I(N__17573));
    Odrv4 I__3894 (
            .O(N__17579),
            .I(\c0.d_4_21 ));
    LocalMux I__3893 (
            .O(N__17576),
            .I(\c0.d_4_21 ));
    LocalMux I__3892 (
            .O(N__17573),
            .I(\c0.d_4_21 ));
    CascadeMux I__3891 (
            .O(N__17566),
            .I(\c0.tx2_data_RNO_4Z0Z_5_cascade_ ));
    InMux I__3890 (
            .O(N__17563),
            .I(N__17560));
    LocalMux I__3889 (
            .O(N__17560),
            .I(\c0.tx2_data_RNO_0Z0Z_5 ));
    CascadeMux I__3888 (
            .O(N__17557),
            .I(\c0.m75_ns_1_cascade_ ));
    InMux I__3887 (
            .O(N__17554),
            .I(N__17551));
    LocalMux I__3886 (
            .O(N__17551),
            .I(N__17548));
    Span4Mux_h I__3885 (
            .O(N__17548),
            .I(N__17545));
    Odrv4 I__3884 (
            .O(N__17545),
            .I(\c0.tx2.r_Tx_DataZ0Z_5 ));
    InMux I__3883 (
            .O(N__17542),
            .I(N__17539));
    LocalMux I__3882 (
            .O(N__17539),
            .I(N__17536));
    Odrv4 I__3881 (
            .O(N__17536),
            .I(\c0.data_in_frame_6_Z0Z_5 ));
    CascadeMux I__3880 (
            .O(N__17533),
            .I(N__17530));
    InMux I__3879 (
            .O(N__17530),
            .I(N__17527));
    LocalMux I__3878 (
            .O(N__17527),
            .I(N__17524));
    Odrv4 I__3877 (
            .O(N__17524),
            .I(\c0.data_in_frame_7_Z0Z_5 ));
    InMux I__3876 (
            .O(N__17521),
            .I(N__17518));
    LocalMux I__3875 (
            .O(N__17518),
            .I(\c0.tx2_data_RNO_1Z0Z_5 ));
    InMux I__3874 (
            .O(N__17515),
            .I(N__17511));
    InMux I__3873 (
            .O(N__17514),
            .I(N__17508));
    LocalMux I__3872 (
            .O(N__17511),
            .I(N__17505));
    LocalMux I__3871 (
            .O(N__17508),
            .I(N__17501));
    Span4Mux_v I__3870 (
            .O(N__17505),
            .I(N__17498));
    InMux I__3869 (
            .O(N__17504),
            .I(N__17495));
    Span12Mux_v I__3868 (
            .O(N__17501),
            .I(N__17492));
    Odrv4 I__3867 (
            .O(N__17498),
            .I(\c0.d_4_47 ));
    LocalMux I__3866 (
            .O(N__17495),
            .I(\c0.d_4_47 ));
    Odrv12 I__3865 (
            .O(N__17492),
            .I(\c0.d_4_47 ));
    CascadeMux I__3864 (
            .O(N__17485),
            .I(N__17481));
    CascadeMux I__3863 (
            .O(N__17484),
            .I(N__17478));
    InMux I__3862 (
            .O(N__17481),
            .I(N__17475));
    InMux I__3861 (
            .O(N__17478),
            .I(N__17472));
    LocalMux I__3860 (
            .O(N__17475),
            .I(N__17469));
    LocalMux I__3859 (
            .O(N__17472),
            .I(N__17466));
    Span4Mux_h I__3858 (
            .O(N__17469),
            .I(N__17460));
    Span4Mux_h I__3857 (
            .O(N__17466),
            .I(N__17460));
    InMux I__3856 (
            .O(N__17465),
            .I(N__17457));
    Odrv4 I__3855 (
            .O(N__17460),
            .I(\c0.d_4_39 ));
    LocalMux I__3854 (
            .O(N__17457),
            .I(\c0.d_4_39 ));
    InMux I__3853 (
            .O(N__17452),
            .I(N__17449));
    LocalMux I__3852 (
            .O(N__17449),
            .I(N__17446));
    Span4Mux_v I__3851 (
            .O(N__17446),
            .I(N__17443));
    Odrv4 I__3850 (
            .O(N__17443),
            .I(\c0.tx2_data_RNO_0Z0Z_7 ));
    InMux I__3849 (
            .O(N__17440),
            .I(N__17437));
    LocalMux I__3848 (
            .O(N__17437),
            .I(N__17434));
    Span4Mux_v I__3847 (
            .O(N__17434),
            .I(N__17431));
    Span4Mux_h I__3846 (
            .O(N__17431),
            .I(N__17428));
    Odrv4 I__3845 (
            .O(N__17428),
            .I(\c0.data_in_frame_6_Z0Z_0 ));
    CascadeMux I__3844 (
            .O(N__17425),
            .I(N__17422));
    InMux I__3843 (
            .O(N__17422),
            .I(N__17419));
    LocalMux I__3842 (
            .O(N__17419),
            .I(N__17416));
    Odrv12 I__3841 (
            .O(N__17416),
            .I(\c0.data_in_frame_7_Z0Z_0 ));
    CascadeMux I__3840 (
            .O(N__17413),
            .I(\c0.tx2.N_493_cascade_ ));
    InMux I__3839 (
            .O(N__17410),
            .I(N__17407));
    LocalMux I__3838 (
            .O(N__17407),
            .I(\c0.tx2.N_205_mux ));
    IoInMux I__3837 (
            .O(N__17404),
            .I(N__17401));
    LocalMux I__3836 (
            .O(N__17401),
            .I(N__17398));
    IoSpan4Mux I__3835 (
            .O(N__17398),
            .I(N__17395));
    Span4Mux_s1_h I__3834 (
            .O(N__17395),
            .I(N__17392));
    Sp12to4 I__3833 (
            .O(N__17392),
            .I(N__17388));
    CascadeMux I__3832 (
            .O(N__17391),
            .I(N__17385));
    Span12Mux_h I__3831 (
            .O(N__17388),
            .I(N__17382));
    InMux I__3830 (
            .O(N__17385),
            .I(N__17379));
    Odrv12 I__3829 (
            .O(N__17382),
            .I(PIN_3_c));
    LocalMux I__3828 (
            .O(N__17379),
            .I(PIN_3_c));
    InMux I__3827 (
            .O(N__17374),
            .I(N__17371));
    LocalMux I__3826 (
            .O(N__17371),
            .I(N__17366));
    CascadeMux I__3825 (
            .O(N__17370),
            .I(N__17363));
    InMux I__3824 (
            .O(N__17369),
            .I(N__17360));
    Span4Mux_v I__3823 (
            .O(N__17366),
            .I(N__17357));
    InMux I__3822 (
            .O(N__17363),
            .I(N__17354));
    LocalMux I__3821 (
            .O(N__17360),
            .I(N__17351));
    Sp12to4 I__3820 (
            .O(N__17357),
            .I(N__17346));
    LocalMux I__3819 (
            .O(N__17354),
            .I(N__17346));
    Odrv12 I__3818 (
            .O(N__17351),
            .I(\c0.data_in_7_Z0Z_0 ));
    Odrv12 I__3817 (
            .O(N__17346),
            .I(\c0.data_in_7_Z0Z_0 ));
    InMux I__3816 (
            .O(N__17341),
            .I(N__17338));
    LocalMux I__3815 (
            .O(N__17338),
            .I(N__17334));
    InMux I__3814 (
            .O(N__17337),
            .I(N__17330));
    Span4Mux_v I__3813 (
            .O(N__17334),
            .I(N__17327));
    InMux I__3812 (
            .O(N__17333),
            .I(N__17324));
    LocalMux I__3811 (
            .O(N__17330),
            .I(N__17321));
    Sp12to4 I__3810 (
            .O(N__17327),
            .I(N__17316));
    LocalMux I__3809 (
            .O(N__17324),
            .I(N__17316));
    Odrv4 I__3808 (
            .O(N__17321),
            .I(\c0.data_in_7_Z0Z_1 ));
    Odrv12 I__3807 (
            .O(N__17316),
            .I(\c0.data_in_7_Z0Z_1 ));
    InMux I__3806 (
            .O(N__17311),
            .I(N__17308));
    LocalMux I__3805 (
            .O(N__17308),
            .I(N__17305));
    Span4Mux_v I__3804 (
            .O(N__17305),
            .I(N__17302));
    Odrv4 I__3803 (
            .O(N__17302),
            .I(\c0.data_in_frame_7_Z0Z_1 ));
    InMux I__3802 (
            .O(N__17299),
            .I(N__17296));
    LocalMux I__3801 (
            .O(N__17296),
            .I(N__17293));
    Span4Mux_v I__3800 (
            .O(N__17293),
            .I(N__17288));
    InMux I__3799 (
            .O(N__17292),
            .I(N__17285));
    InMux I__3798 (
            .O(N__17291),
            .I(N__17282));
    Odrv4 I__3797 (
            .O(N__17288),
            .I(\c0.data_in_6_Z0Z_5 ));
    LocalMux I__3796 (
            .O(N__17285),
            .I(\c0.data_in_6_Z0Z_5 ));
    LocalMux I__3795 (
            .O(N__17282),
            .I(\c0.data_in_6_Z0Z_5 ));
    CascadeMux I__3794 (
            .O(N__17275),
            .I(N__17272));
    InMux I__3793 (
            .O(N__17272),
            .I(N__17267));
    InMux I__3792 (
            .O(N__17271),
            .I(N__17264));
    InMux I__3791 (
            .O(N__17270),
            .I(N__17261));
    LocalMux I__3790 (
            .O(N__17267),
            .I(N__17258));
    LocalMux I__3789 (
            .O(N__17264),
            .I(\c0.data_in_7_Z0Z_5 ));
    LocalMux I__3788 (
            .O(N__17261),
            .I(\c0.data_in_7_Z0Z_5 ));
    Odrv4 I__3787 (
            .O(N__17258),
            .I(\c0.data_in_7_Z0Z_5 ));
    InMux I__3786 (
            .O(N__17251),
            .I(N__17248));
    LocalMux I__3785 (
            .O(N__17248),
            .I(N__17243));
    InMux I__3784 (
            .O(N__17247),
            .I(N__17240));
    InMux I__3783 (
            .O(N__17246),
            .I(N__17237));
    Span4Mux_h I__3782 (
            .O(N__17243),
            .I(N__17234));
    LocalMux I__3781 (
            .O(N__17240),
            .I(\c0.data_in_7_Z0Z_6 ));
    LocalMux I__3780 (
            .O(N__17237),
            .I(\c0.data_in_7_Z0Z_6 ));
    Odrv4 I__3779 (
            .O(N__17234),
            .I(\c0.data_in_7_Z0Z_6 ));
    InMux I__3778 (
            .O(N__17227),
            .I(N__17224));
    LocalMux I__3777 (
            .O(N__17224),
            .I(\c0.data_in_frame_7_Z0Z_6 ));
    CascadeMux I__3776 (
            .O(N__17221),
            .I(N__17218));
    InMux I__3775 (
            .O(N__17218),
            .I(N__17213));
    InMux I__3774 (
            .O(N__17217),
            .I(N__17210));
    InMux I__3773 (
            .O(N__17216),
            .I(N__17207));
    LocalMux I__3772 (
            .O(N__17213),
            .I(N__17204));
    LocalMux I__3771 (
            .O(N__17210),
            .I(\c0.data_in_6_Z0Z_6 ));
    LocalMux I__3770 (
            .O(N__17207),
            .I(\c0.data_in_6_Z0Z_6 ));
    Odrv12 I__3769 (
            .O(N__17204),
            .I(\c0.data_in_6_Z0Z_6 ));
    InMux I__3768 (
            .O(N__17197),
            .I(N__17194));
    LocalMux I__3767 (
            .O(N__17194),
            .I(N__17191));
    Odrv4 I__3766 (
            .O(N__17191),
            .I(\c0.data_in_frame_6_Z0Z_6 ));
    CEMux I__3765 (
            .O(N__17188),
            .I(N__17131));
    CEMux I__3764 (
            .O(N__17187),
            .I(N__17131));
    CEMux I__3763 (
            .O(N__17186),
            .I(N__17131));
    CEMux I__3762 (
            .O(N__17185),
            .I(N__17131));
    CEMux I__3761 (
            .O(N__17184),
            .I(N__17131));
    CEMux I__3760 (
            .O(N__17183),
            .I(N__17131));
    CEMux I__3759 (
            .O(N__17182),
            .I(N__17131));
    CEMux I__3758 (
            .O(N__17181),
            .I(N__17131));
    CEMux I__3757 (
            .O(N__17180),
            .I(N__17131));
    CEMux I__3756 (
            .O(N__17179),
            .I(N__17131));
    CEMux I__3755 (
            .O(N__17178),
            .I(N__17131));
    CEMux I__3754 (
            .O(N__17177),
            .I(N__17131));
    CEMux I__3753 (
            .O(N__17176),
            .I(N__17131));
    CEMux I__3752 (
            .O(N__17175),
            .I(N__17131));
    CEMux I__3751 (
            .O(N__17174),
            .I(N__17131));
    CEMux I__3750 (
            .O(N__17173),
            .I(N__17131));
    CEMux I__3749 (
            .O(N__17172),
            .I(N__17131));
    CEMux I__3748 (
            .O(N__17171),
            .I(N__17131));
    CEMux I__3747 (
            .O(N__17170),
            .I(N__17131));
    GlobalMux I__3746 (
            .O(N__17131),
            .I(N__17128));
    gio2CtrlBuf I__3745 (
            .O(N__17128),
            .I(\c0.data_in_frame_0__0_sqmuxa_g ));
    InMux I__3744 (
            .O(N__17125),
            .I(N__17122));
    LocalMux I__3743 (
            .O(N__17122),
            .I(\c0.tx2.r_Clock_Count_i_3 ));
    InMux I__3742 (
            .O(N__17119),
            .I(\c0.tx2.r_Clock_Count12 ));
    CascadeMux I__3741 (
            .O(N__17116),
            .I(N__17109));
    CascadeMux I__3740 (
            .O(N__17115),
            .I(N__17106));
    CascadeMux I__3739 (
            .O(N__17114),
            .I(N__17100));
    CascadeMux I__3738 (
            .O(N__17113),
            .I(N__17097));
    CascadeMux I__3737 (
            .O(N__17112),
            .I(N__17094));
    InMux I__3736 (
            .O(N__17109),
            .I(N__17076));
    InMux I__3735 (
            .O(N__17106),
            .I(N__17076));
    InMux I__3734 (
            .O(N__17105),
            .I(N__17076));
    InMux I__3733 (
            .O(N__17104),
            .I(N__17076));
    InMux I__3732 (
            .O(N__17103),
            .I(N__17071));
    InMux I__3731 (
            .O(N__17100),
            .I(N__17068));
    InMux I__3730 (
            .O(N__17097),
            .I(N__17061));
    InMux I__3729 (
            .O(N__17094),
            .I(N__17061));
    InMux I__3728 (
            .O(N__17093),
            .I(N__17061));
    CascadeMux I__3727 (
            .O(N__17092),
            .I(N__17057));
    InMux I__3726 (
            .O(N__17091),
            .I(N__17053));
    InMux I__3725 (
            .O(N__17090),
            .I(N__17040));
    InMux I__3724 (
            .O(N__17089),
            .I(N__17040));
    InMux I__3723 (
            .O(N__17088),
            .I(N__17040));
    InMux I__3722 (
            .O(N__17087),
            .I(N__17040));
    InMux I__3721 (
            .O(N__17086),
            .I(N__17040));
    InMux I__3720 (
            .O(N__17085),
            .I(N__17040));
    LocalMux I__3719 (
            .O(N__17076),
            .I(N__17037));
    InMux I__3718 (
            .O(N__17075),
            .I(N__17032));
    InMux I__3717 (
            .O(N__17074),
            .I(N__17032));
    LocalMux I__3716 (
            .O(N__17071),
            .I(N__17029));
    LocalMux I__3715 (
            .O(N__17068),
            .I(N__17024));
    LocalMux I__3714 (
            .O(N__17061),
            .I(N__17024));
    InMux I__3713 (
            .O(N__17060),
            .I(N__17021));
    InMux I__3712 (
            .O(N__17057),
            .I(N__17015));
    InMux I__3711 (
            .O(N__17056),
            .I(N__17012));
    LocalMux I__3710 (
            .O(N__17053),
            .I(N__17001));
    LocalMux I__3709 (
            .O(N__17040),
            .I(N__17001));
    Span4Mux_v I__3708 (
            .O(N__17037),
            .I(N__16996));
    LocalMux I__3707 (
            .O(N__17032),
            .I(N__16996));
    Span4Mux_h I__3706 (
            .O(N__17029),
            .I(N__16991));
    Span4Mux_v I__3705 (
            .O(N__17024),
            .I(N__16991));
    LocalMux I__3704 (
            .O(N__17021),
            .I(N__16988));
    InMux I__3703 (
            .O(N__17020),
            .I(N__16981));
    InMux I__3702 (
            .O(N__17019),
            .I(N__16981));
    InMux I__3701 (
            .O(N__17018),
            .I(N__16981));
    LocalMux I__3700 (
            .O(N__17015),
            .I(N__16976));
    LocalMux I__3699 (
            .O(N__17012),
            .I(N__16976));
    InMux I__3698 (
            .O(N__17011),
            .I(N__16967));
    InMux I__3697 (
            .O(N__17010),
            .I(N__16967));
    InMux I__3696 (
            .O(N__17009),
            .I(N__16967));
    InMux I__3695 (
            .O(N__17008),
            .I(N__16967));
    InMux I__3694 (
            .O(N__17007),
            .I(N__16962));
    InMux I__3693 (
            .O(N__17006),
            .I(N__16962));
    Span4Mux_v I__3692 (
            .O(N__17001),
            .I(N__16952));
    Span4Mux_h I__3691 (
            .O(N__16996),
            .I(N__16949));
    Span4Mux_h I__3690 (
            .O(N__16991),
            .I(N__16942));
    Span4Mux_h I__3689 (
            .O(N__16988),
            .I(N__16942));
    LocalMux I__3688 (
            .O(N__16981),
            .I(N__16942));
    Span12Mux_v I__3687 (
            .O(N__16976),
            .I(N__16935));
    LocalMux I__3686 (
            .O(N__16967),
            .I(N__16935));
    LocalMux I__3685 (
            .O(N__16962),
            .I(N__16935));
    InMux I__3684 (
            .O(N__16961),
            .I(N__16920));
    InMux I__3683 (
            .O(N__16960),
            .I(N__16920));
    InMux I__3682 (
            .O(N__16959),
            .I(N__16920));
    InMux I__3681 (
            .O(N__16958),
            .I(N__16920));
    InMux I__3680 (
            .O(N__16957),
            .I(N__16920));
    InMux I__3679 (
            .O(N__16956),
            .I(N__16920));
    InMux I__3678 (
            .O(N__16955),
            .I(N__16920));
    Odrv4 I__3677 (
            .O(N__16952),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3676 (
            .O(N__16949),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3675 (
            .O(N__16942),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3674 (
            .O(N__16935),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3673 (
            .O(N__16920),
            .I(CONSTANT_ONE_NET));
    InMux I__3672 (
            .O(N__16909),
            .I(N__16906));
    LocalMux I__3671 (
            .O(N__16906),
            .I(N__16902));
    InMux I__3670 (
            .O(N__16905),
            .I(N__16899));
    Span4Mux_v I__3669 (
            .O(N__16902),
            .I(N__16896));
    LocalMux I__3668 (
            .O(N__16899),
            .I(N__16893));
    Span4Mux_h I__3667 (
            .O(N__16896),
            .I(N__16890));
    Span4Mux_h I__3666 (
            .O(N__16893),
            .I(N__16887));
    Odrv4 I__3665 (
            .O(N__16890),
            .I(\c0.d_2_29 ));
    Odrv4 I__3664 (
            .O(N__16887),
            .I(\c0.d_2_29 ));
    SRMux I__3663 (
            .O(N__16882),
            .I(N__16869));
    SRMux I__3662 (
            .O(N__16881),
            .I(N__16866));
    SRMux I__3661 (
            .O(N__16880),
            .I(N__16863));
    SRMux I__3660 (
            .O(N__16879),
            .I(N__16860));
    SRMux I__3659 (
            .O(N__16878),
            .I(N__16857));
    SRMux I__3658 (
            .O(N__16877),
            .I(N__16854));
    SRMux I__3657 (
            .O(N__16876),
            .I(N__16851));
    SRMux I__3656 (
            .O(N__16875),
            .I(N__16848));
    SRMux I__3655 (
            .O(N__16874),
            .I(N__16845));
    SRMux I__3654 (
            .O(N__16873),
            .I(N__16842));
    SRMux I__3653 (
            .O(N__16872),
            .I(N__16839));
    LocalMux I__3652 (
            .O(N__16869),
            .I(N__16821));
    LocalMux I__3651 (
            .O(N__16866),
            .I(N__16818));
    LocalMux I__3650 (
            .O(N__16863),
            .I(N__16815));
    LocalMux I__3649 (
            .O(N__16860),
            .I(N__16812));
    LocalMux I__3648 (
            .O(N__16857),
            .I(N__16809));
    LocalMux I__3647 (
            .O(N__16854),
            .I(N__16806));
    LocalMux I__3646 (
            .O(N__16851),
            .I(N__16803));
    LocalMux I__3645 (
            .O(N__16848),
            .I(N__16800));
    LocalMux I__3644 (
            .O(N__16845),
            .I(N__16797));
    LocalMux I__3643 (
            .O(N__16842),
            .I(N__16794));
    LocalMux I__3642 (
            .O(N__16839),
            .I(N__16791));
    CEMux I__3641 (
            .O(N__16838),
            .I(N__16738));
    CEMux I__3640 (
            .O(N__16837),
            .I(N__16738));
    CEMux I__3639 (
            .O(N__16836),
            .I(N__16738));
    CEMux I__3638 (
            .O(N__16835),
            .I(N__16738));
    CEMux I__3637 (
            .O(N__16834),
            .I(N__16738));
    CEMux I__3636 (
            .O(N__16833),
            .I(N__16738));
    CEMux I__3635 (
            .O(N__16832),
            .I(N__16738));
    CEMux I__3634 (
            .O(N__16831),
            .I(N__16738));
    CEMux I__3633 (
            .O(N__16830),
            .I(N__16738));
    CEMux I__3632 (
            .O(N__16829),
            .I(N__16738));
    CEMux I__3631 (
            .O(N__16828),
            .I(N__16738));
    CEMux I__3630 (
            .O(N__16827),
            .I(N__16738));
    CEMux I__3629 (
            .O(N__16826),
            .I(N__16738));
    CEMux I__3628 (
            .O(N__16825),
            .I(N__16738));
    CEMux I__3627 (
            .O(N__16824),
            .I(N__16738));
    Glb2LocalMux I__3626 (
            .O(N__16821),
            .I(N__16738));
    Glb2LocalMux I__3625 (
            .O(N__16818),
            .I(N__16738));
    Glb2LocalMux I__3624 (
            .O(N__16815),
            .I(N__16738));
    Glb2LocalMux I__3623 (
            .O(N__16812),
            .I(N__16738));
    Glb2LocalMux I__3622 (
            .O(N__16809),
            .I(N__16738));
    Glb2LocalMux I__3621 (
            .O(N__16806),
            .I(N__16738));
    Glb2LocalMux I__3620 (
            .O(N__16803),
            .I(N__16738));
    Glb2LocalMux I__3619 (
            .O(N__16800),
            .I(N__16738));
    Glb2LocalMux I__3618 (
            .O(N__16797),
            .I(N__16738));
    Glb2LocalMux I__3617 (
            .O(N__16794),
            .I(N__16738));
    Glb2LocalMux I__3616 (
            .O(N__16791),
            .I(N__16738));
    GlobalMux I__3615 (
            .O(N__16738),
            .I(N__16735));
    gio2CtrlBuf I__3614 (
            .O(N__16735),
            .I(\c0.data_out_0__1_sqmuxa_g ));
    InMux I__3613 (
            .O(N__16732),
            .I(N__16729));
    LocalMux I__3612 (
            .O(N__16729),
            .I(N__16726));
    Span4Mux_v I__3611 (
            .O(N__16726),
            .I(N__16723));
    Odrv4 I__3610 (
            .O(N__16723),
            .I(\c0.tx2.r_Tx_DataZ0Z_6 ));
    InMux I__3609 (
            .O(N__16720),
            .I(N__16717));
    LocalMux I__3608 (
            .O(N__16717),
            .I(N__16714));
    Span4Mux_h I__3607 (
            .O(N__16714),
            .I(N__16711));
    Odrv4 I__3606 (
            .O(N__16711),
            .I(\c0.tx2.r_Tx_DataZ0Z_2 ));
    CascadeMux I__3605 (
            .O(N__16708),
            .I(\c0.tx2.o_Tx_Serial_RNOZ0Z_6_cascade_ ));
    InMux I__3604 (
            .O(N__16705),
            .I(N__16702));
    LocalMux I__3603 (
            .O(N__16702),
            .I(N__16699));
    Odrv4 I__3602 (
            .O(N__16699),
            .I(\c0.tx2.o_Tx_Serial_RNOZ0Z_5 ));
    InMux I__3601 (
            .O(N__16696),
            .I(N__16693));
    LocalMux I__3600 (
            .O(N__16693),
            .I(\c0.tx2.o_Tx_Serial_RNOZ0Z_3 ));
    CascadeMux I__3599 (
            .O(N__16690),
            .I(\c0.tx2.m195_ns_1_cascade_ ));
    InMux I__3598 (
            .O(N__16687),
            .I(N__16684));
    LocalMux I__3597 (
            .O(N__16684),
            .I(N__16681));
    Odrv4 I__3596 (
            .O(N__16681),
            .I(\c0.tx2.o_Tx_Serial_RNOZ0Z_2 ));
    CascadeMux I__3595 (
            .O(N__16678),
            .I(\c0.tx2.N_196_0_cascade_ ));
    CascadeMux I__3594 (
            .O(N__16675),
            .I(N__16671));
    InMux I__3593 (
            .O(N__16674),
            .I(N__16667));
    InMux I__3592 (
            .O(N__16671),
            .I(N__16664));
    InMux I__3591 (
            .O(N__16670),
            .I(N__16661));
    LocalMux I__3590 (
            .O(N__16667),
            .I(N__16656));
    LocalMux I__3589 (
            .O(N__16664),
            .I(N__16656));
    LocalMux I__3588 (
            .O(N__16661),
            .I(\c0.d_4_1 ));
    Odrv4 I__3587 (
            .O(N__16656),
            .I(\c0.d_4_1 ));
    InMux I__3586 (
            .O(N__16651),
            .I(N__16648));
    LocalMux I__3585 (
            .O(N__16648),
            .I(N__16643));
    InMux I__3584 (
            .O(N__16647),
            .I(N__16638));
    InMux I__3583 (
            .O(N__16646),
            .I(N__16638));
    Odrv4 I__3582 (
            .O(N__16643),
            .I(\c0.d_4_9 ));
    LocalMux I__3581 (
            .O(N__16638),
            .I(\c0.d_4_9 ));
    InMux I__3580 (
            .O(N__16633),
            .I(N__16630));
    LocalMux I__3579 (
            .O(N__16630),
            .I(N__16627));
    Odrv12 I__3578 (
            .O(N__16627),
            .I(\c0.tx2_data_RNO_3Z0Z_1 ));
    InMux I__3577 (
            .O(N__16624),
            .I(N__16621));
    LocalMux I__3576 (
            .O(N__16621),
            .I(N__16618));
    Odrv4 I__3575 (
            .O(N__16618),
            .I(\c0.tx2.r_Tx_DataZ0Z_1 ));
    CascadeMux I__3574 (
            .O(N__16615),
            .I(N__16612));
    InMux I__3573 (
            .O(N__16612),
            .I(N__16609));
    LocalMux I__3572 (
            .O(N__16609),
            .I(N__16606));
    Span4Mux_h I__3571 (
            .O(N__16606),
            .I(N__16603));
    Span4Mux_h I__3570 (
            .O(N__16603),
            .I(N__16600));
    Odrv4 I__3569 (
            .O(N__16600),
            .I(\c0.data_in_frame_6_Z0Z_1 ));
    InMux I__3568 (
            .O(N__16597),
            .I(N__16594));
    LocalMux I__3567 (
            .O(N__16594),
            .I(N__16591));
    Odrv12 I__3566 (
            .O(N__16591),
            .I(\c0.tx2_data_RNO_1Z0Z_1 ));
    InMux I__3565 (
            .O(N__16588),
            .I(N__16585));
    LocalMux I__3564 (
            .O(N__16585),
            .I(N__16582));
    Odrv12 I__3563 (
            .O(N__16582),
            .I(\c0.tx2.r_Tx_DataZ0Z_4 ));
    InMux I__3562 (
            .O(N__16579),
            .I(N__16576));
    LocalMux I__3561 (
            .O(N__16576),
            .I(N__16573));
    Odrv4 I__3560 (
            .O(N__16573),
            .I(\c0.N_173_0 ));
    InMux I__3559 (
            .O(N__16570),
            .I(N__16566));
    InMux I__3558 (
            .O(N__16569),
            .I(N__16563));
    LocalMux I__3557 (
            .O(N__16566),
            .I(\c0.tx2.r_Clock_Count_i_0 ));
    LocalMux I__3556 (
            .O(N__16563),
            .I(\c0.tx2.r_Clock_Count_i_0 ));
    InMux I__3555 (
            .O(N__16558),
            .I(N__16555));
    LocalMux I__3554 (
            .O(N__16555),
            .I(\c0.tx2.r_Clock_Count_i_1 ));
    InMux I__3553 (
            .O(N__16552),
            .I(N__16549));
    LocalMux I__3552 (
            .O(N__16549),
            .I(\c0.tx2.r_Clock_Count_i_2 ));
    InMux I__3551 (
            .O(N__16546),
            .I(N__16539));
    InMux I__3550 (
            .O(N__16545),
            .I(N__16539));
    InMux I__3549 (
            .O(N__16544),
            .I(N__16536));
    LocalMux I__3548 (
            .O(N__16539),
            .I(N__16533));
    LocalMux I__3547 (
            .O(N__16536),
            .I(N__16529));
    Span4Mux_h I__3546 (
            .O(N__16533),
            .I(N__16526));
    InMux I__3545 (
            .O(N__16532),
            .I(N__16523));
    Odrv4 I__3544 (
            .O(N__16529),
            .I(\c0.N_123 ));
    Odrv4 I__3543 (
            .O(N__16526),
            .I(\c0.N_123 ));
    LocalMux I__3542 (
            .O(N__16523),
            .I(\c0.N_123 ));
    InMux I__3541 (
            .O(N__16516),
            .I(N__16512));
    InMux I__3540 (
            .O(N__16515),
            .I(N__16509));
    LocalMux I__3539 (
            .O(N__16512),
            .I(N__16506));
    LocalMux I__3538 (
            .O(N__16509),
            .I(N__16502));
    Span4Mux_v I__3537 (
            .O(N__16506),
            .I(N__16498));
    InMux I__3536 (
            .O(N__16505),
            .I(N__16495));
    Span4Mux_h I__3535 (
            .O(N__16502),
            .I(N__16492));
    InMux I__3534 (
            .O(N__16501),
            .I(N__16489));
    Odrv4 I__3533 (
            .O(N__16498),
            .I(\c0.d_4_15 ));
    LocalMux I__3532 (
            .O(N__16495),
            .I(\c0.d_4_15 ));
    Odrv4 I__3531 (
            .O(N__16492),
            .I(\c0.d_4_15 ));
    LocalMux I__3530 (
            .O(N__16489),
            .I(\c0.d_4_15 ));
    InMux I__3529 (
            .O(N__16480),
            .I(N__16477));
    LocalMux I__3528 (
            .O(N__16477),
            .I(\c0.N_129 ));
    CascadeMux I__3527 (
            .O(N__16474),
            .I(N__16470));
    InMux I__3526 (
            .O(N__16473),
            .I(N__16467));
    InMux I__3525 (
            .O(N__16470),
            .I(N__16464));
    LocalMux I__3524 (
            .O(N__16467),
            .I(\c0.N_18 ));
    LocalMux I__3523 (
            .O(N__16464),
            .I(\c0.N_18 ));
    InMux I__3522 (
            .O(N__16459),
            .I(\c0.un1_byte_transmit_counter2_1_cry_0 ));
    InMux I__3521 (
            .O(N__16456),
            .I(\c0.un1_byte_transmit_counter2_1_cry_1 ));
    InMux I__3520 (
            .O(N__16453),
            .I(\c0.un1_byte_transmit_counter2_1_cry_2 ));
    InMux I__3519 (
            .O(N__16450),
            .I(\c0.un1_byte_transmit_counter2_1_cry_3 ));
    InMux I__3518 (
            .O(N__16447),
            .I(\c0.un1_byte_transmit_counter2_1_cry_4 ));
    InMux I__3517 (
            .O(N__16444),
            .I(\c0.un1_byte_transmit_counter2_1_cry_5 ));
    InMux I__3516 (
            .O(N__16441),
            .I(\c0.un1_byte_transmit_counter2_1_cry_6 ));
    CascadeMux I__3515 (
            .O(N__16438),
            .I(N__16431));
    InMux I__3514 (
            .O(N__16437),
            .I(N__16428));
    InMux I__3513 (
            .O(N__16436),
            .I(N__16423));
    InMux I__3512 (
            .O(N__16435),
            .I(N__16423));
    InMux I__3511 (
            .O(N__16434),
            .I(N__16420));
    InMux I__3510 (
            .O(N__16431),
            .I(N__16417));
    LocalMux I__3509 (
            .O(N__16428),
            .I(N__16414));
    LocalMux I__3508 (
            .O(N__16423),
            .I(\c0.d_4_38 ));
    LocalMux I__3507 (
            .O(N__16420),
            .I(\c0.d_4_38 ));
    LocalMux I__3506 (
            .O(N__16417),
            .I(\c0.d_4_38 ));
    Odrv4 I__3505 (
            .O(N__16414),
            .I(\c0.d_4_38 ));
    InMux I__3504 (
            .O(N__16405),
            .I(N__16400));
    InMux I__3503 (
            .O(N__16404),
            .I(N__16397));
    InMux I__3502 (
            .O(N__16403),
            .I(N__16394));
    LocalMux I__3501 (
            .O(N__16400),
            .I(N__16391));
    LocalMux I__3500 (
            .O(N__16397),
            .I(\c0.N_107 ));
    LocalMux I__3499 (
            .O(N__16394),
            .I(\c0.N_107 ));
    Odrv4 I__3498 (
            .O(N__16391),
            .I(\c0.N_107 ));
    CascadeMux I__3497 (
            .O(N__16384),
            .I(\c0.un1_data_in_6__2_0_a2_6_a2_2_cascade_ ));
    InMux I__3496 (
            .O(N__16381),
            .I(N__16378));
    LocalMux I__3495 (
            .O(N__16378),
            .I(N__16375));
    Odrv4 I__3494 (
            .O(N__16375),
            .I(\c0.un1_data_in_6__2 ));
    CascadeMux I__3493 (
            .O(N__16372),
            .I(N__16368));
    CascadeMux I__3492 (
            .O(N__16371),
            .I(N__16364));
    InMux I__3491 (
            .O(N__16368),
            .I(N__16361));
    InMux I__3490 (
            .O(N__16367),
            .I(N__16358));
    InMux I__3489 (
            .O(N__16364),
            .I(N__16355));
    LocalMux I__3488 (
            .O(N__16361),
            .I(N__16350));
    LocalMux I__3487 (
            .O(N__16358),
            .I(N__16350));
    LocalMux I__3486 (
            .O(N__16355),
            .I(N__16347));
    Span4Mux_v I__3485 (
            .O(N__16350),
            .I(N__16344));
    Span4Mux_v I__3484 (
            .O(N__16347),
            .I(N__16341));
    Odrv4 I__3483 (
            .O(N__16344),
            .I(\c0.d_4_46 ));
    Odrv4 I__3482 (
            .O(N__16341),
            .I(\c0.d_4_46 ));
    InMux I__3481 (
            .O(N__16336),
            .I(N__16332));
    InMux I__3480 (
            .O(N__16335),
            .I(N__16329));
    LocalMux I__3479 (
            .O(N__16332),
            .I(N__16324));
    LocalMux I__3478 (
            .O(N__16329),
            .I(N__16321));
    InMux I__3477 (
            .O(N__16328),
            .I(N__16318));
    InMux I__3476 (
            .O(N__16327),
            .I(N__16315));
    Odrv4 I__3475 (
            .O(N__16324),
            .I(\c0.d_4_42 ));
    Odrv4 I__3474 (
            .O(N__16321),
            .I(\c0.d_4_42 ));
    LocalMux I__3473 (
            .O(N__16318),
            .I(\c0.d_4_42 ));
    LocalMux I__3472 (
            .O(N__16315),
            .I(\c0.d_4_42 ));
    InMux I__3471 (
            .O(N__16306),
            .I(N__16303));
    LocalMux I__3470 (
            .O(N__16303),
            .I(N__16298));
    InMux I__3469 (
            .O(N__16302),
            .I(N__16295));
    InMux I__3468 (
            .O(N__16301),
            .I(N__16292));
    Odrv4 I__3467 (
            .O(N__16298),
            .I(\c0.N_133 ));
    LocalMux I__3466 (
            .O(N__16295),
            .I(\c0.N_133 ));
    LocalMux I__3465 (
            .O(N__16292),
            .I(\c0.N_133 ));
    CascadeMux I__3464 (
            .O(N__16285),
            .I(\c0.un1_data_in_7__2_0_a2_0_a2_5_cascade_ ));
    InMux I__3463 (
            .O(N__16282),
            .I(N__16279));
    LocalMux I__3462 (
            .O(N__16279),
            .I(N__16276));
    Odrv4 I__3461 (
            .O(N__16276),
            .I(\c0.un1_data_in_7__2 ));
    InMux I__3460 (
            .O(N__16273),
            .I(N__16269));
    InMux I__3459 (
            .O(N__16272),
            .I(N__16265));
    LocalMux I__3458 (
            .O(N__16269),
            .I(N__16262));
    InMux I__3457 (
            .O(N__16268),
            .I(N__16259));
    LocalMux I__3456 (
            .O(N__16265),
            .I(N__16256));
    Span4Mux_v I__3455 (
            .O(N__16262),
            .I(N__16253));
    LocalMux I__3454 (
            .O(N__16259),
            .I(\c0.d_4_14 ));
    Odrv4 I__3453 (
            .O(N__16256),
            .I(\c0.d_4_14 ));
    Odrv4 I__3452 (
            .O(N__16253),
            .I(\c0.d_4_14 ));
    InMux I__3451 (
            .O(N__16246),
            .I(N__16239));
    InMux I__3450 (
            .O(N__16245),
            .I(N__16236));
    InMux I__3449 (
            .O(N__16244),
            .I(N__16229));
    InMux I__3448 (
            .O(N__16243),
            .I(N__16229));
    InMux I__3447 (
            .O(N__16242),
            .I(N__16229));
    LocalMux I__3446 (
            .O(N__16239),
            .I(\c0.d_4_31 ));
    LocalMux I__3445 (
            .O(N__16236),
            .I(\c0.d_4_31 ));
    LocalMux I__3444 (
            .O(N__16229),
            .I(\c0.d_4_31 ));
    InMux I__3443 (
            .O(N__16222),
            .I(N__16219));
    LocalMux I__3442 (
            .O(N__16219),
            .I(N__16216));
    Odrv4 I__3441 (
            .O(N__16216),
            .I(\c0.un1_data_in_7__2_0_a2_0_a2_4 ));
    InMux I__3440 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__3439 (
            .O(N__16210),
            .I(N__16207));
    Span4Mux_v I__3438 (
            .O(N__16207),
            .I(N__16204));
    Span4Mux_h I__3437 (
            .O(N__16204),
            .I(N__16201));
    Odrv4 I__3436 (
            .O(N__16201),
            .I(\c0.un1_data_in_7__3_0_a2_0_a2_3 ));
    InMux I__3435 (
            .O(N__16198),
            .I(N__16194));
    InMux I__3434 (
            .O(N__16197),
            .I(N__16191));
    LocalMux I__3433 (
            .O(N__16194),
            .I(N__16188));
    LocalMux I__3432 (
            .O(N__16191),
            .I(N__16185));
    Span4Mux_v I__3431 (
            .O(N__16188),
            .I(N__16180));
    Span4Mux_h I__3430 (
            .O(N__16185),
            .I(N__16177));
    InMux I__3429 (
            .O(N__16184),
            .I(N__16174));
    InMux I__3428 (
            .O(N__16183),
            .I(N__16171));
    Odrv4 I__3427 (
            .O(N__16180),
            .I(\c0.d_4_43 ));
    Odrv4 I__3426 (
            .O(N__16177),
            .I(\c0.d_4_43 ));
    LocalMux I__3425 (
            .O(N__16174),
            .I(\c0.d_4_43 ));
    LocalMux I__3424 (
            .O(N__16171),
            .I(\c0.d_4_43 ));
    InMux I__3423 (
            .O(N__16162),
            .I(N__16158));
    InMux I__3422 (
            .O(N__16161),
            .I(N__16154));
    LocalMux I__3421 (
            .O(N__16158),
            .I(N__16151));
    InMux I__3420 (
            .O(N__16157),
            .I(N__16148));
    LocalMux I__3419 (
            .O(N__16154),
            .I(\c0.N_128 ));
    Odrv4 I__3418 (
            .O(N__16151),
            .I(\c0.N_128 ));
    LocalMux I__3417 (
            .O(N__16148),
            .I(\c0.N_128 ));
    CascadeMux I__3416 (
            .O(N__16141),
            .I(\c0.un1_data_in_7__3_0_a2_0_a2_4_cascade_ ));
    InMux I__3415 (
            .O(N__16138),
            .I(N__16135));
    LocalMux I__3414 (
            .O(N__16135),
            .I(\c0.un1_data_in_7__5_0_a2_0_a2_1 ));
    InMux I__3413 (
            .O(N__16132),
            .I(N__16129));
    LocalMux I__3412 (
            .O(N__16129),
            .I(N__16126));
    Odrv4 I__3411 (
            .O(N__16126),
            .I(\c0.m163_9 ));
    InMux I__3410 (
            .O(N__16123),
            .I(N__16120));
    LocalMux I__3409 (
            .O(N__16120),
            .I(N__16117));
    Span4Mux_h I__3408 (
            .O(N__16117),
            .I(N__16114));
    Span4Mux_h I__3407 (
            .O(N__16114),
            .I(N__16110));
    InMux I__3406 (
            .O(N__16113),
            .I(N__16107));
    Odrv4 I__3405 (
            .O(N__16110),
            .I(\c0.data_in_0_Z0Z_1 ));
    LocalMux I__3404 (
            .O(N__16107),
            .I(\c0.data_in_0_Z0Z_1 ));
    InMux I__3403 (
            .O(N__16102),
            .I(N__16099));
    LocalMux I__3402 (
            .O(N__16099),
            .I(N__16095));
    InMux I__3401 (
            .O(N__16098),
            .I(N__16092));
    Odrv12 I__3400 (
            .O(N__16095),
            .I(\c0.data_in_4_Z0Z_6 ));
    LocalMux I__3399 (
            .O(N__16092),
            .I(\c0.data_in_4_Z0Z_6 ));
    InMux I__3398 (
            .O(N__16087),
            .I(N__16084));
    LocalMux I__3397 (
            .O(N__16084),
            .I(N__16081));
    Span4Mux_v I__3396 (
            .O(N__16081),
            .I(N__16077));
    InMux I__3395 (
            .O(N__16080),
            .I(N__16074));
    Odrv4 I__3394 (
            .O(N__16077),
            .I(\c0.data_in_5_Z0Z_6 ));
    LocalMux I__3393 (
            .O(N__16074),
            .I(\c0.data_in_5_Z0Z_6 ));
    InMux I__3392 (
            .O(N__16069),
            .I(N__16065));
    InMux I__3391 (
            .O(N__16068),
            .I(N__16062));
    LocalMux I__3390 (
            .O(N__16065),
            .I(N__16059));
    LocalMux I__3389 (
            .O(N__16062),
            .I(N__16056));
    Odrv12 I__3388 (
            .O(N__16059),
            .I(\c0.rx_data_6 ));
    Odrv4 I__3387 (
            .O(N__16056),
            .I(\c0.rx_data_6 ));
    InMux I__3386 (
            .O(N__16051),
            .I(N__16047));
    InMux I__3385 (
            .O(N__16050),
            .I(N__16043));
    LocalMux I__3384 (
            .O(N__16047),
            .I(N__16040));
    InMux I__3383 (
            .O(N__16046),
            .I(N__16036));
    LocalMux I__3382 (
            .O(N__16043),
            .I(N__16033));
    Span4Mux_v I__3381 (
            .O(N__16040),
            .I(N__16030));
    InMux I__3380 (
            .O(N__16039),
            .I(N__16027));
    LocalMux I__3379 (
            .O(N__16036),
            .I(N__16024));
    Odrv12 I__3378 (
            .O(N__16033),
            .I(\c0.d_4_26 ));
    Odrv4 I__3377 (
            .O(N__16030),
            .I(\c0.d_4_26 ));
    LocalMux I__3376 (
            .O(N__16027),
            .I(\c0.d_4_26 ));
    Odrv4 I__3375 (
            .O(N__16024),
            .I(\c0.d_4_26 ));
    InMux I__3374 (
            .O(N__16015),
            .I(N__16012));
    LocalMux I__3373 (
            .O(N__16012),
            .I(N__16007));
    InMux I__3372 (
            .O(N__16011),
            .I(N__16004));
    CascadeMux I__3371 (
            .O(N__16010),
            .I(N__16001));
    Span4Mux_h I__3370 (
            .O(N__16007),
            .I(N__15998));
    LocalMux I__3369 (
            .O(N__16004),
            .I(N__15995));
    InMux I__3368 (
            .O(N__16001),
            .I(N__15992));
    Odrv4 I__3367 (
            .O(N__15998),
            .I(\c0.data_in_6_Z0Z_4 ));
    Odrv4 I__3366 (
            .O(N__15995),
            .I(\c0.data_in_6_Z0Z_4 ));
    LocalMux I__3365 (
            .O(N__15992),
            .I(\c0.data_in_6_Z0Z_4 ));
    InMux I__3364 (
            .O(N__15985),
            .I(N__15982));
    LocalMux I__3363 (
            .O(N__15982),
            .I(N__15977));
    InMux I__3362 (
            .O(N__15981),
            .I(N__15974));
    CascadeMux I__3361 (
            .O(N__15980),
            .I(N__15971));
    Span4Mux_v I__3360 (
            .O(N__15977),
            .I(N__15966));
    LocalMux I__3359 (
            .O(N__15974),
            .I(N__15966));
    InMux I__3358 (
            .O(N__15971),
            .I(N__15963));
    Span4Mux_h I__3357 (
            .O(N__15966),
            .I(N__15959));
    LocalMux I__3356 (
            .O(N__15963),
            .I(N__15956));
    InMux I__3355 (
            .O(N__15962),
            .I(N__15953));
    Odrv4 I__3354 (
            .O(N__15959),
            .I(\c0.d_4_41 ));
    Odrv4 I__3353 (
            .O(N__15956),
            .I(\c0.d_4_41 ));
    LocalMux I__3352 (
            .O(N__15953),
            .I(\c0.d_4_41 ));
    CascadeMux I__3351 (
            .O(N__15946),
            .I(N__15943));
    InMux I__3350 (
            .O(N__15943),
            .I(N__15940));
    LocalMux I__3349 (
            .O(N__15940),
            .I(\c0.un1_data_in_6__4_0_a2_5_a2_1 ));
    InMux I__3348 (
            .O(N__15937),
            .I(N__15934));
    LocalMux I__3347 (
            .O(N__15934),
            .I(N__15930));
    CascadeMux I__3346 (
            .O(N__15933),
            .I(N__15926));
    Span4Mux_v I__3345 (
            .O(N__15930),
            .I(N__15923));
    InMux I__3344 (
            .O(N__15929),
            .I(N__15918));
    InMux I__3343 (
            .O(N__15926),
            .I(N__15918));
    Span4Mux_h I__3342 (
            .O(N__15923),
            .I(N__15913));
    LocalMux I__3341 (
            .O(N__15918),
            .I(N__15913));
    Odrv4 I__3340 (
            .O(N__15913),
            .I(\c0.data_in_1_Z0Z_2 ));
    InMux I__3339 (
            .O(N__15910),
            .I(N__15907));
    LocalMux I__3338 (
            .O(N__15907),
            .I(N__15902));
    InMux I__3337 (
            .O(N__15906),
            .I(N__15897));
    InMux I__3336 (
            .O(N__15905),
            .I(N__15897));
    Odrv4 I__3335 (
            .O(N__15902),
            .I(\c0.d_4_10 ));
    LocalMux I__3334 (
            .O(N__15897),
            .I(\c0.d_4_10 ));
    InMux I__3333 (
            .O(N__15892),
            .I(N__15888));
    InMux I__3332 (
            .O(N__15891),
            .I(N__15885));
    LocalMux I__3331 (
            .O(N__15888),
            .I(N__15882));
    LocalMux I__3330 (
            .O(N__15885),
            .I(\c0.N_127 ));
    Odrv12 I__3329 (
            .O(N__15882),
            .I(\c0.N_127 ));
    InMux I__3328 (
            .O(N__15877),
            .I(N__15874));
    LocalMux I__3327 (
            .O(N__15874),
            .I(N__15871));
    Span12Mux_h I__3326 (
            .O(N__15871),
            .I(N__15866));
    InMux I__3325 (
            .O(N__15870),
            .I(N__15863));
    InMux I__3324 (
            .O(N__15869),
            .I(N__15860));
    Odrv12 I__3323 (
            .O(N__15866),
            .I(\c0.data_in_1_Z0Z_1 ));
    LocalMux I__3322 (
            .O(N__15863),
            .I(\c0.data_in_1_Z0Z_1 ));
    LocalMux I__3321 (
            .O(N__15860),
            .I(\c0.data_in_1_Z0Z_1 ));
    InMux I__3320 (
            .O(N__15853),
            .I(N__15850));
    LocalMux I__3319 (
            .O(N__15850),
            .I(N__15846));
    InMux I__3318 (
            .O(N__15849),
            .I(N__15843));
    Span4Mux_h I__3317 (
            .O(N__15846),
            .I(N__15839));
    LocalMux I__3316 (
            .O(N__15843),
            .I(N__15836));
    InMux I__3315 (
            .O(N__15842),
            .I(N__15833));
    Odrv4 I__3314 (
            .O(N__15839),
            .I(\c0.data_in_3_Z0Z_1 ));
    Odrv4 I__3313 (
            .O(N__15836),
            .I(\c0.data_in_3_Z0Z_1 ));
    LocalMux I__3312 (
            .O(N__15833),
            .I(\c0.data_in_3_Z0Z_1 ));
    InMux I__3311 (
            .O(N__15826),
            .I(N__15823));
    LocalMux I__3310 (
            .O(N__15823),
            .I(N__15820));
    Span4Mux_h I__3309 (
            .O(N__15820),
            .I(N__15815));
    InMux I__3308 (
            .O(N__15819),
            .I(N__15812));
    InMux I__3307 (
            .O(N__15818),
            .I(N__15809));
    Odrv4 I__3306 (
            .O(N__15815),
            .I(\c0.d_4_25 ));
    LocalMux I__3305 (
            .O(N__15812),
            .I(\c0.d_4_25 ));
    LocalMux I__3304 (
            .O(N__15809),
            .I(\c0.d_4_25 ));
    InMux I__3303 (
            .O(N__15802),
            .I(N__15799));
    LocalMux I__3302 (
            .O(N__15799),
            .I(\c0.data_in_frame_6_Z0Z_4 ));
    InMux I__3301 (
            .O(N__15796),
            .I(N__15793));
    LocalMux I__3300 (
            .O(N__15793),
            .I(\c0.data_in_frame_7_Z0Z_4 ));
    InMux I__3299 (
            .O(N__15790),
            .I(N__15787));
    LocalMux I__3298 (
            .O(N__15787),
            .I(\c0.tx2_data_RNO_1Z0Z_4 ));
    InMux I__3297 (
            .O(N__15784),
            .I(N__15781));
    LocalMux I__3296 (
            .O(N__15781),
            .I(\c0.tx2_data_RNO_0Z0Z_4 ));
    CascadeMux I__3295 (
            .O(N__15778),
            .I(\c0.m120_ns_1_cascade_ ));
    InMux I__3294 (
            .O(N__15775),
            .I(N__15772));
    LocalMux I__3293 (
            .O(N__15772),
            .I(\c0.tx2_data_RNO_3Z0Z_6 ));
    InMux I__3292 (
            .O(N__15769),
            .I(N__15766));
    LocalMux I__3291 (
            .O(N__15766),
            .I(\c0.tx2_data_RNO_0Z0Z_6 ));
    CascadeMux I__3290 (
            .O(N__15763),
            .I(\c0.m90_ns_1_cascade_ ));
    InMux I__3289 (
            .O(N__15760),
            .I(N__15757));
    LocalMux I__3288 (
            .O(N__15757),
            .I(\c0.tx2_data_RNO_1Z0Z_6 ));
    InMux I__3287 (
            .O(N__15754),
            .I(N__15751));
    LocalMux I__3286 (
            .O(N__15751),
            .I(N__15747));
    InMux I__3285 (
            .O(N__15750),
            .I(N__15743));
    Span4Mux_h I__3284 (
            .O(N__15747),
            .I(N__15740));
    InMux I__3283 (
            .O(N__15746),
            .I(N__15737));
    LocalMux I__3282 (
            .O(N__15743),
            .I(N__15734));
    Odrv4 I__3281 (
            .O(N__15740),
            .I(\c0.data_in_7_Z0Z_4 ));
    LocalMux I__3280 (
            .O(N__15737),
            .I(\c0.data_in_7_Z0Z_4 ));
    Odrv12 I__3279 (
            .O(N__15734),
            .I(\c0.data_in_7_Z0Z_4 ));
    InMux I__3278 (
            .O(N__15727),
            .I(N__15724));
    LocalMux I__3277 (
            .O(N__15724),
            .I(N__15721));
    Span4Mux_h I__3276 (
            .O(N__15721),
            .I(N__15718));
    Span4Mux_h I__3275 (
            .O(N__15718),
            .I(N__15714));
    InMux I__3274 (
            .O(N__15717),
            .I(N__15711));
    Odrv4 I__3273 (
            .O(N__15714),
            .I(\c0.rx_data_5 ));
    LocalMux I__3272 (
            .O(N__15711),
            .I(\c0.rx_data_5 ));
    InMux I__3271 (
            .O(N__15706),
            .I(N__15699));
    InMux I__3270 (
            .O(N__15705),
            .I(N__15699));
    InMux I__3269 (
            .O(N__15704),
            .I(N__15696));
    LocalMux I__3268 (
            .O(N__15699),
            .I(N__15693));
    LocalMux I__3267 (
            .O(N__15696),
            .I(N__15690));
    Span4Mux_h I__3266 (
            .O(N__15693),
            .I(N__15687));
    Odrv4 I__3265 (
            .O(N__15690),
            .I(\c0.d_2_10 ));
    Odrv4 I__3264 (
            .O(N__15687),
            .I(\c0.d_2_10 ));
    InMux I__3263 (
            .O(N__15682),
            .I(N__15679));
    LocalMux I__3262 (
            .O(N__15679),
            .I(\c0.byte_transmit_counterZ0Z_6 ));
    InMux I__3261 (
            .O(N__15676),
            .I(N__15673));
    LocalMux I__3260 (
            .O(N__15673),
            .I(\c0.byte_transmit_counterZ0Z_7 ));
    InMux I__3259 (
            .O(N__15670),
            .I(N__15667));
    LocalMux I__3258 (
            .O(N__15667),
            .I(\c0.byte_transmit_counterZ0Z_3 ));
    InMux I__3257 (
            .O(N__15664),
            .I(N__15661));
    LocalMux I__3256 (
            .O(N__15661),
            .I(\c0.byte_transmit_counterZ0Z_4 ));
    InMux I__3255 (
            .O(N__15658),
            .I(N__15653));
    InMux I__3254 (
            .O(N__15657),
            .I(N__15647));
    InMux I__3253 (
            .O(N__15656),
            .I(N__15644));
    LocalMux I__3252 (
            .O(N__15653),
            .I(N__15641));
    InMux I__3251 (
            .O(N__15652),
            .I(N__15637));
    InMux I__3250 (
            .O(N__15651),
            .I(N__15634));
    InMux I__3249 (
            .O(N__15650),
            .I(N__15628));
    LocalMux I__3248 (
            .O(N__15647),
            .I(N__15625));
    LocalMux I__3247 (
            .O(N__15644),
            .I(N__15622));
    Span4Mux_h I__3246 (
            .O(N__15641),
            .I(N__15619));
    InMux I__3245 (
            .O(N__15640),
            .I(N__15616));
    LocalMux I__3244 (
            .O(N__15637),
            .I(N__15611));
    LocalMux I__3243 (
            .O(N__15634),
            .I(N__15611));
    InMux I__3242 (
            .O(N__15633),
            .I(N__15607));
    InMux I__3241 (
            .O(N__15632),
            .I(N__15604));
    InMux I__3240 (
            .O(N__15631),
            .I(N__15601));
    LocalMux I__3239 (
            .O(N__15628),
            .I(N__15596));
    Span4Mux_h I__3238 (
            .O(N__15625),
            .I(N__15596));
    Span4Mux_h I__3237 (
            .O(N__15622),
            .I(N__15593));
    Span4Mux_h I__3236 (
            .O(N__15619),
            .I(N__15586));
    LocalMux I__3235 (
            .O(N__15616),
            .I(N__15586));
    Span4Mux_h I__3234 (
            .O(N__15611),
            .I(N__15586));
    InMux I__3233 (
            .O(N__15610),
            .I(N__15583));
    LocalMux I__3232 (
            .O(N__15607),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    LocalMux I__3231 (
            .O(N__15604),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    LocalMux I__3230 (
            .O(N__15601),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    Odrv4 I__3229 (
            .O(N__15596),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    Odrv4 I__3228 (
            .O(N__15593),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    Odrv4 I__3227 (
            .O(N__15586),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    LocalMux I__3226 (
            .O(N__15583),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    CascadeMux I__3225 (
            .O(N__15568),
            .I(N__15562));
    CascadeMux I__3224 (
            .O(N__15567),
            .I(N__15559));
    InMux I__3223 (
            .O(N__15566),
            .I(N__15550));
    InMux I__3222 (
            .O(N__15565),
            .I(N__15550));
    InMux I__3221 (
            .O(N__15562),
            .I(N__15541));
    InMux I__3220 (
            .O(N__15559),
            .I(N__15541));
    InMux I__3219 (
            .O(N__15558),
            .I(N__15541));
    InMux I__3218 (
            .O(N__15557),
            .I(N__15541));
    InMux I__3217 (
            .O(N__15556),
            .I(N__15523));
    InMux I__3216 (
            .O(N__15555),
            .I(N__15523));
    LocalMux I__3215 (
            .O(N__15550),
            .I(N__15518));
    LocalMux I__3214 (
            .O(N__15541),
            .I(N__15518));
    CascadeMux I__3213 (
            .O(N__15540),
            .I(N__15512));
    CascadeMux I__3212 (
            .O(N__15539),
            .I(N__15507));
    CascadeMux I__3211 (
            .O(N__15538),
            .I(N__15504));
    InMux I__3210 (
            .O(N__15537),
            .I(N__15489));
    InMux I__3209 (
            .O(N__15536),
            .I(N__15489));
    InMux I__3208 (
            .O(N__15535),
            .I(N__15489));
    InMux I__3207 (
            .O(N__15534),
            .I(N__15489));
    InMux I__3206 (
            .O(N__15533),
            .I(N__15489));
    InMux I__3205 (
            .O(N__15532),
            .I(N__15482));
    InMux I__3204 (
            .O(N__15531),
            .I(N__15482));
    InMux I__3203 (
            .O(N__15530),
            .I(N__15482));
    InMux I__3202 (
            .O(N__15529),
            .I(N__15479));
    CascadeMux I__3201 (
            .O(N__15528),
            .I(N__15475));
    LocalMux I__3200 (
            .O(N__15523),
            .I(N__15466));
    Span4Mux_h I__3199 (
            .O(N__15518),
            .I(N__15466));
    InMux I__3198 (
            .O(N__15517),
            .I(N__15463));
    InMux I__3197 (
            .O(N__15516),
            .I(N__15460));
    InMux I__3196 (
            .O(N__15515),
            .I(N__15451));
    InMux I__3195 (
            .O(N__15512),
            .I(N__15451));
    InMux I__3194 (
            .O(N__15511),
            .I(N__15451));
    InMux I__3193 (
            .O(N__15510),
            .I(N__15451));
    InMux I__3192 (
            .O(N__15507),
            .I(N__15438));
    InMux I__3191 (
            .O(N__15504),
            .I(N__15438));
    InMux I__3190 (
            .O(N__15503),
            .I(N__15438));
    InMux I__3189 (
            .O(N__15502),
            .I(N__15438));
    InMux I__3188 (
            .O(N__15501),
            .I(N__15438));
    InMux I__3187 (
            .O(N__15500),
            .I(N__15438));
    LocalMux I__3186 (
            .O(N__15489),
            .I(N__15435));
    LocalMux I__3185 (
            .O(N__15482),
            .I(N__15430));
    LocalMux I__3184 (
            .O(N__15479),
            .I(N__15430));
    InMux I__3183 (
            .O(N__15478),
            .I(N__15426));
    InMux I__3182 (
            .O(N__15475),
            .I(N__15421));
    InMux I__3181 (
            .O(N__15474),
            .I(N__15421));
    InMux I__3180 (
            .O(N__15473),
            .I(N__15416));
    InMux I__3179 (
            .O(N__15472),
            .I(N__15416));
    InMux I__3178 (
            .O(N__15471),
            .I(N__15413));
    Span4Mux_v I__3177 (
            .O(N__15466),
            .I(N__15410));
    LocalMux I__3176 (
            .O(N__15463),
            .I(N__15397));
    LocalMux I__3175 (
            .O(N__15460),
            .I(N__15397));
    LocalMux I__3174 (
            .O(N__15451),
            .I(N__15397));
    LocalMux I__3173 (
            .O(N__15438),
            .I(N__15397));
    Span4Mux_v I__3172 (
            .O(N__15435),
            .I(N__15397));
    Span4Mux_h I__3171 (
            .O(N__15430),
            .I(N__15397));
    InMux I__3170 (
            .O(N__15429),
            .I(N__15394));
    LocalMux I__3169 (
            .O(N__15426),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    LocalMux I__3168 (
            .O(N__15421),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    LocalMux I__3167 (
            .O(N__15416),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    LocalMux I__3166 (
            .O(N__15413),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    Odrv4 I__3165 (
            .O(N__15410),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    Odrv4 I__3164 (
            .O(N__15397),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    LocalMux I__3163 (
            .O(N__15394),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    InMux I__3162 (
            .O(N__15379),
            .I(N__15376));
    LocalMux I__3161 (
            .O(N__15376),
            .I(N__15361));
    InMux I__3160 (
            .O(N__15375),
            .I(N__15356));
    InMux I__3159 (
            .O(N__15374),
            .I(N__15356));
    InMux I__3158 (
            .O(N__15373),
            .I(N__15347));
    InMux I__3157 (
            .O(N__15372),
            .I(N__15347));
    InMux I__3156 (
            .O(N__15371),
            .I(N__15347));
    InMux I__3155 (
            .O(N__15370),
            .I(N__15347));
    InMux I__3154 (
            .O(N__15369),
            .I(N__15321));
    InMux I__3153 (
            .O(N__15368),
            .I(N__15321));
    InMux I__3152 (
            .O(N__15367),
            .I(N__15321));
    InMux I__3151 (
            .O(N__15366),
            .I(N__15321));
    InMux I__3150 (
            .O(N__15365),
            .I(N__15321));
    InMux I__3149 (
            .O(N__15364),
            .I(N__15318));
    Span4Mux_v I__3148 (
            .O(N__15361),
            .I(N__15311));
    LocalMux I__3147 (
            .O(N__15356),
            .I(N__15311));
    LocalMux I__3146 (
            .O(N__15347),
            .I(N__15311));
    InMux I__3145 (
            .O(N__15346),
            .I(N__15304));
    InMux I__3144 (
            .O(N__15345),
            .I(N__15304));
    InMux I__3143 (
            .O(N__15344),
            .I(N__15304));
    InMux I__3142 (
            .O(N__15343),
            .I(N__15295));
    InMux I__3141 (
            .O(N__15342),
            .I(N__15295));
    InMux I__3140 (
            .O(N__15341),
            .I(N__15295));
    InMux I__3139 (
            .O(N__15340),
            .I(N__15295));
    InMux I__3138 (
            .O(N__15339),
            .I(N__15290));
    InMux I__3137 (
            .O(N__15338),
            .I(N__15290));
    InMux I__3136 (
            .O(N__15337),
            .I(N__15279));
    InMux I__3135 (
            .O(N__15336),
            .I(N__15274));
    InMux I__3134 (
            .O(N__15335),
            .I(N__15274));
    InMux I__3133 (
            .O(N__15334),
            .I(N__15271));
    InMux I__3132 (
            .O(N__15333),
            .I(N__15268));
    InMux I__3131 (
            .O(N__15332),
            .I(N__15265));
    LocalMux I__3130 (
            .O(N__15321),
            .I(N__15262));
    LocalMux I__3129 (
            .O(N__15318),
            .I(N__15251));
    Span4Mux_h I__3128 (
            .O(N__15311),
            .I(N__15251));
    LocalMux I__3127 (
            .O(N__15304),
            .I(N__15251));
    LocalMux I__3126 (
            .O(N__15295),
            .I(N__15251));
    LocalMux I__3125 (
            .O(N__15290),
            .I(N__15251));
    InMux I__3124 (
            .O(N__15289),
            .I(N__15238));
    InMux I__3123 (
            .O(N__15288),
            .I(N__15238));
    InMux I__3122 (
            .O(N__15287),
            .I(N__15238));
    InMux I__3121 (
            .O(N__15286),
            .I(N__15238));
    InMux I__3120 (
            .O(N__15285),
            .I(N__15238));
    InMux I__3119 (
            .O(N__15284),
            .I(N__15238));
    InMux I__3118 (
            .O(N__15283),
            .I(N__15233));
    InMux I__3117 (
            .O(N__15282),
            .I(N__15233));
    LocalMux I__3116 (
            .O(N__15279),
            .I(\c0.N_132_mux ));
    LocalMux I__3115 (
            .O(N__15274),
            .I(\c0.N_132_mux ));
    LocalMux I__3114 (
            .O(N__15271),
            .I(\c0.N_132_mux ));
    LocalMux I__3113 (
            .O(N__15268),
            .I(\c0.N_132_mux ));
    LocalMux I__3112 (
            .O(N__15265),
            .I(\c0.N_132_mux ));
    Odrv12 I__3111 (
            .O(N__15262),
            .I(\c0.N_132_mux ));
    Odrv4 I__3110 (
            .O(N__15251),
            .I(\c0.N_132_mux ));
    LocalMux I__3109 (
            .O(N__15238),
            .I(\c0.N_132_mux ));
    LocalMux I__3108 (
            .O(N__15233),
            .I(\c0.N_132_mux ));
    CascadeMux I__3107 (
            .O(N__15214),
            .I(N__15206));
    CascadeMux I__3106 (
            .O(N__15213),
            .I(N__15203));
    CascadeMux I__3105 (
            .O(N__15212),
            .I(N__15200));
    CascadeMux I__3104 (
            .O(N__15211),
            .I(N__15194));
    CascadeMux I__3103 (
            .O(N__15210),
            .I(N__15191));
    CascadeMux I__3102 (
            .O(N__15209),
            .I(N__15188));
    InMux I__3101 (
            .O(N__15206),
            .I(N__15183));
    InMux I__3100 (
            .O(N__15203),
            .I(N__15174));
    InMux I__3099 (
            .O(N__15200),
            .I(N__15174));
    InMux I__3098 (
            .O(N__15199),
            .I(N__15174));
    InMux I__3097 (
            .O(N__15198),
            .I(N__15174));
    InMux I__3096 (
            .O(N__15197),
            .I(N__15171));
    InMux I__3095 (
            .O(N__15194),
            .I(N__15168));
    InMux I__3094 (
            .O(N__15191),
            .I(N__15156));
    InMux I__3093 (
            .O(N__15188),
            .I(N__15156));
    InMux I__3092 (
            .O(N__15187),
            .I(N__15156));
    InMux I__3091 (
            .O(N__15186),
            .I(N__15153));
    LocalMux I__3090 (
            .O(N__15183),
            .I(N__15146));
    LocalMux I__3089 (
            .O(N__15174),
            .I(N__15146));
    LocalMux I__3088 (
            .O(N__15171),
            .I(N__15146));
    LocalMux I__3087 (
            .O(N__15168),
            .I(N__15143));
    InMux I__3086 (
            .O(N__15167),
            .I(N__15140));
    InMux I__3085 (
            .O(N__15166),
            .I(N__15137));
    InMux I__3084 (
            .O(N__15165),
            .I(N__15134));
    InMux I__3083 (
            .O(N__15164),
            .I(N__15130));
    InMux I__3082 (
            .O(N__15163),
            .I(N__15127));
    LocalMux I__3081 (
            .O(N__15156),
            .I(N__15120));
    LocalMux I__3080 (
            .O(N__15153),
            .I(N__15120));
    Span4Mux_h I__3079 (
            .O(N__15146),
            .I(N__15120));
    Span4Mux_h I__3078 (
            .O(N__15143),
            .I(N__15111));
    LocalMux I__3077 (
            .O(N__15140),
            .I(N__15111));
    LocalMux I__3076 (
            .O(N__15137),
            .I(N__15111));
    LocalMux I__3075 (
            .O(N__15134),
            .I(N__15111));
    InMux I__3074 (
            .O(N__15133),
            .I(N__15107));
    LocalMux I__3073 (
            .O(N__15130),
            .I(N__15102));
    LocalMux I__3072 (
            .O(N__15127),
            .I(N__15102));
    Span4Mux_v I__3071 (
            .O(N__15120),
            .I(N__15099));
    Span4Mux_v I__3070 (
            .O(N__15111),
            .I(N__15096));
    InMux I__3069 (
            .O(N__15110),
            .I(N__15093));
    LocalMux I__3068 (
            .O(N__15107),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    Odrv12 I__3067 (
            .O(N__15102),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    Odrv4 I__3066 (
            .O(N__15099),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    Odrv4 I__3065 (
            .O(N__15096),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    LocalMux I__3064 (
            .O(N__15093),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    CascadeMux I__3063 (
            .O(N__15082),
            .I(\c0.N_5_1_cascade_ ));
    CEMux I__3062 (
            .O(N__15079),
            .I(N__15076));
    LocalMux I__3061 (
            .O(N__15076),
            .I(N__15072));
    CEMux I__3060 (
            .O(N__15075),
            .I(N__15069));
    Span4Mux_h I__3059 (
            .O(N__15072),
            .I(N__15064));
    LocalMux I__3058 (
            .O(N__15069),
            .I(N__15064));
    Span4Mux_v I__3057 (
            .O(N__15064),
            .I(N__15060));
    InMux I__3056 (
            .O(N__15063),
            .I(N__15057));
    Sp12to4 I__3055 (
            .O(N__15060),
            .I(N__15052));
    LocalMux I__3054 (
            .O(N__15057),
            .I(N__15052));
    Span12Mux_s11_v I__3053 (
            .O(N__15052),
            .I(N__15049));
    Odrv12 I__3052 (
            .O(N__15049),
            .I(\c0.byte_transmit_counter15 ));
    IoInMux I__3051 (
            .O(N__15046),
            .I(N__15043));
    LocalMux I__3050 (
            .O(N__15043),
            .I(N__15040));
    Span4Mux_s0_v I__3049 (
            .O(N__15040),
            .I(N__15037));
    Span4Mux_v I__3048 (
            .O(N__15037),
            .I(N__15034));
    Odrv4 I__3047 (
            .O(N__15034),
            .I(\c0.data_out_0__1_sqmuxa ));
    InMux I__3046 (
            .O(N__15031),
            .I(N__15027));
    InMux I__3045 (
            .O(N__15030),
            .I(N__15023));
    LocalMux I__3044 (
            .O(N__15027),
            .I(N__15020));
    CascadeMux I__3043 (
            .O(N__15026),
            .I(N__15017));
    LocalMux I__3042 (
            .O(N__15023),
            .I(N__15014));
    Span4Mux_h I__3041 (
            .O(N__15020),
            .I(N__15011));
    InMux I__3040 (
            .O(N__15017),
            .I(N__15008));
    Odrv12 I__3039 (
            .O(N__15014),
            .I(\c0.d_2_14 ));
    Odrv4 I__3038 (
            .O(N__15011),
            .I(\c0.d_2_14 ));
    LocalMux I__3037 (
            .O(N__15008),
            .I(\c0.d_2_14 ));
    CascadeMux I__3036 (
            .O(N__15001),
            .I(N__14998));
    InMux I__3035 (
            .O(N__14998),
            .I(N__14994));
    InMux I__3034 (
            .O(N__14997),
            .I(N__14990));
    LocalMux I__3033 (
            .O(N__14994),
            .I(N__14987));
    InMux I__3032 (
            .O(N__14993),
            .I(N__14984));
    LocalMux I__3031 (
            .O(N__14990),
            .I(N__14980));
    Span4Mux_h I__3030 (
            .O(N__14987),
            .I(N__14977));
    LocalMux I__3029 (
            .O(N__14984),
            .I(N__14974));
    InMux I__3028 (
            .O(N__14983),
            .I(N__14971));
    Span4Mux_h I__3027 (
            .O(N__14980),
            .I(N__14968));
    Odrv4 I__3026 (
            .O(N__14977),
            .I(\c0.d_2_30 ));
    Odrv4 I__3025 (
            .O(N__14974),
            .I(\c0.d_2_30 ));
    LocalMux I__3024 (
            .O(N__14971),
            .I(\c0.d_2_30 ));
    Odrv4 I__3023 (
            .O(N__14968),
            .I(\c0.d_2_30 ));
    InMux I__3022 (
            .O(N__14959),
            .I(N__14954));
    InMux I__3021 (
            .O(N__14958),
            .I(N__14949));
    InMux I__3020 (
            .O(N__14957),
            .I(N__14949));
    LocalMux I__3019 (
            .O(N__14954),
            .I(N__14946));
    LocalMux I__3018 (
            .O(N__14949),
            .I(N__14941));
    Span4Mux_v I__3017 (
            .O(N__14946),
            .I(N__14941));
    Odrv4 I__3016 (
            .O(N__14941),
            .I(\c0.d_2_16 ));
    CascadeMux I__3015 (
            .O(N__14938),
            .I(N__14935));
    InMux I__3014 (
            .O(N__14935),
            .I(N__14930));
    InMux I__3013 (
            .O(N__14934),
            .I(N__14927));
    InMux I__3012 (
            .O(N__14933),
            .I(N__14923));
    LocalMux I__3011 (
            .O(N__14930),
            .I(N__14920));
    LocalMux I__3010 (
            .O(N__14927),
            .I(N__14917));
    InMux I__3009 (
            .O(N__14926),
            .I(N__14914));
    LocalMux I__3008 (
            .O(N__14923),
            .I(N__14907));
    Span4Mux_v I__3007 (
            .O(N__14920),
            .I(N__14907));
    Span4Mux_v I__3006 (
            .O(N__14917),
            .I(N__14907));
    LocalMux I__3005 (
            .O(N__14914),
            .I(\c0.d_2_17 ));
    Odrv4 I__3004 (
            .O(N__14907),
            .I(\c0.d_2_17 ));
    CascadeMux I__3003 (
            .O(N__14902),
            .I(N__14899));
    InMux I__3002 (
            .O(N__14899),
            .I(N__14896));
    LocalMux I__3001 (
            .O(N__14896),
            .I(N__14891));
    InMux I__3000 (
            .O(N__14895),
            .I(N__14886));
    InMux I__2999 (
            .O(N__14894),
            .I(N__14886));
    Span4Mux_h I__2998 (
            .O(N__14891),
            .I(N__14883));
    LocalMux I__2997 (
            .O(N__14886),
            .I(N__14880));
    Odrv4 I__2996 (
            .O(N__14883),
            .I(\c0.d_2_12 ));
    Odrv4 I__2995 (
            .O(N__14880),
            .I(\c0.d_2_12 ));
    InMux I__2994 (
            .O(N__14875),
            .I(N__14870));
    InMux I__2993 (
            .O(N__14874),
            .I(N__14867));
    CascadeMux I__2992 (
            .O(N__14873),
            .I(N__14863));
    LocalMux I__2991 (
            .O(N__14870),
            .I(N__14860));
    LocalMux I__2990 (
            .O(N__14867),
            .I(N__14857));
    CascadeMux I__2989 (
            .O(N__14866),
            .I(N__14854));
    InMux I__2988 (
            .O(N__14863),
            .I(N__14851));
    Span12Mux_h I__2987 (
            .O(N__14860),
            .I(N__14848));
    Span4Mux_v I__2986 (
            .O(N__14857),
            .I(N__14845));
    InMux I__2985 (
            .O(N__14854),
            .I(N__14842));
    LocalMux I__2984 (
            .O(N__14851),
            .I(N__14839));
    Odrv12 I__2983 (
            .O(N__14848),
            .I(\c0.d_2_21 ));
    Odrv4 I__2982 (
            .O(N__14845),
            .I(\c0.d_2_21 ));
    LocalMux I__2981 (
            .O(N__14842),
            .I(\c0.d_2_21 ));
    Odrv12 I__2980 (
            .O(N__14839),
            .I(\c0.d_2_21 ));
    CascadeMux I__2979 (
            .O(N__14830),
            .I(N__14826));
    InMux I__2978 (
            .O(N__14829),
            .I(N__14823));
    InMux I__2977 (
            .O(N__14826),
            .I(N__14820));
    LocalMux I__2976 (
            .O(N__14823),
            .I(N__14815));
    LocalMux I__2975 (
            .O(N__14820),
            .I(N__14812));
    InMux I__2974 (
            .O(N__14819),
            .I(N__14807));
    InMux I__2973 (
            .O(N__14818),
            .I(N__14807));
    Span4Mux_h I__2972 (
            .O(N__14815),
            .I(N__14804));
    Span4Mux_v I__2971 (
            .O(N__14812),
            .I(N__14799));
    LocalMux I__2970 (
            .O(N__14807),
            .I(N__14799));
    Odrv4 I__2969 (
            .O(N__14804),
            .I(\c0.d_2_11 ));
    Odrv4 I__2968 (
            .O(N__14799),
            .I(\c0.d_2_11 ));
    InMux I__2967 (
            .O(N__14794),
            .I(N__14790));
    InMux I__2966 (
            .O(N__14793),
            .I(N__14786));
    LocalMux I__2965 (
            .O(N__14790),
            .I(N__14783));
    InMux I__2964 (
            .O(N__14789),
            .I(N__14780));
    LocalMux I__2963 (
            .O(N__14786),
            .I(N__14777));
    Span4Mux_h I__2962 (
            .O(N__14783),
            .I(N__14772));
    LocalMux I__2961 (
            .O(N__14780),
            .I(N__14769));
    Span4Mux_h I__2960 (
            .O(N__14777),
            .I(N__14766));
    InMux I__2959 (
            .O(N__14776),
            .I(N__14763));
    InMux I__2958 (
            .O(N__14775),
            .I(N__14760));
    Odrv4 I__2957 (
            .O(N__14772),
            .I(\c0.d_2_26 ));
    Odrv4 I__2956 (
            .O(N__14769),
            .I(\c0.d_2_26 ));
    Odrv4 I__2955 (
            .O(N__14766),
            .I(\c0.d_2_26 ));
    LocalMux I__2954 (
            .O(N__14763),
            .I(\c0.d_2_26 ));
    LocalMux I__2953 (
            .O(N__14760),
            .I(\c0.d_2_26 ));
    InMux I__2952 (
            .O(N__14749),
            .I(N__14744));
    InMux I__2951 (
            .O(N__14748),
            .I(N__14738));
    InMux I__2950 (
            .O(N__14747),
            .I(N__14738));
    LocalMux I__2949 (
            .O(N__14744),
            .I(N__14735));
    CascadeMux I__2948 (
            .O(N__14743),
            .I(N__14732));
    LocalMux I__2947 (
            .O(N__14738),
            .I(N__14729));
    Span4Mux_h I__2946 (
            .O(N__14735),
            .I(N__14726));
    InMux I__2945 (
            .O(N__14732),
            .I(N__14723));
    Span4Mux_h I__2944 (
            .O(N__14729),
            .I(N__14720));
    Odrv4 I__2943 (
            .O(N__14726),
            .I(\c0.d_2_18 ));
    LocalMux I__2942 (
            .O(N__14723),
            .I(\c0.d_2_18 ));
    Odrv4 I__2941 (
            .O(N__14720),
            .I(\c0.d_2_18 ));
    InMux I__2940 (
            .O(N__14713),
            .I(N__14710));
    LocalMux I__2939 (
            .O(N__14710),
            .I(N__14706));
    InMux I__2938 (
            .O(N__14709),
            .I(N__14701));
    Span4Mux_v I__2937 (
            .O(N__14706),
            .I(N__14697));
    InMux I__2936 (
            .O(N__14705),
            .I(N__14694));
    InMux I__2935 (
            .O(N__14704),
            .I(N__14691));
    LocalMux I__2934 (
            .O(N__14701),
            .I(N__14688));
    InMux I__2933 (
            .O(N__14700),
            .I(N__14685));
    Odrv4 I__2932 (
            .O(N__14697),
            .I(\c0.d_4_35 ));
    LocalMux I__2931 (
            .O(N__14694),
            .I(\c0.d_4_35 ));
    LocalMux I__2930 (
            .O(N__14691),
            .I(\c0.d_4_35 ));
    Odrv12 I__2929 (
            .O(N__14688),
            .I(\c0.d_4_35 ));
    LocalMux I__2928 (
            .O(N__14685),
            .I(\c0.d_4_35 ));
    InMux I__2927 (
            .O(N__14674),
            .I(N__14671));
    LocalMux I__2926 (
            .O(N__14671),
            .I(N__14668));
    Span4Mux_v I__2925 (
            .O(N__14668),
            .I(N__14662));
    InMux I__2924 (
            .O(N__14667),
            .I(N__14657));
    InMux I__2923 (
            .O(N__14666),
            .I(N__14657));
    InMux I__2922 (
            .O(N__14665),
            .I(N__14654));
    Odrv4 I__2921 (
            .O(N__14662),
            .I(\c0.d_4_27 ));
    LocalMux I__2920 (
            .O(N__14657),
            .I(\c0.d_4_27 ));
    LocalMux I__2919 (
            .O(N__14654),
            .I(\c0.d_4_27 ));
    CascadeMux I__2918 (
            .O(N__14647),
            .I(N__14644));
    InMux I__2917 (
            .O(N__14644),
            .I(N__14641));
    LocalMux I__2916 (
            .O(N__14641),
            .I(N__14637));
    InMux I__2915 (
            .O(N__14640),
            .I(N__14634));
    Span4Mux_v I__2914 (
            .O(N__14637),
            .I(N__14629));
    LocalMux I__2913 (
            .O(N__14634),
            .I(N__14629));
    Span4Mux_v I__2912 (
            .O(N__14629),
            .I(N__14625));
    InMux I__2911 (
            .O(N__14628),
            .I(N__14622));
    Odrv4 I__2910 (
            .O(N__14625),
            .I(\c0.d_4_19 ));
    LocalMux I__2909 (
            .O(N__14622),
            .I(\c0.d_4_19 ));
    InMux I__2908 (
            .O(N__14617),
            .I(N__14614));
    LocalMux I__2907 (
            .O(N__14614),
            .I(N__14608));
    InMux I__2906 (
            .O(N__14613),
            .I(N__14603));
    InMux I__2905 (
            .O(N__14612),
            .I(N__14603));
    InMux I__2904 (
            .O(N__14611),
            .I(N__14600));
    Odrv4 I__2903 (
            .O(N__14608),
            .I(\c0.d_4_3 ));
    LocalMux I__2902 (
            .O(N__14603),
            .I(\c0.d_4_3 ));
    LocalMux I__2901 (
            .O(N__14600),
            .I(\c0.d_4_3 ));
    CascadeMux I__2900 (
            .O(N__14593),
            .I(N__14590));
    InMux I__2899 (
            .O(N__14590),
            .I(N__14587));
    LocalMux I__2898 (
            .O(N__14587),
            .I(N__14583));
    InMux I__2897 (
            .O(N__14586),
            .I(N__14580));
    Span4Mux_v I__2896 (
            .O(N__14583),
            .I(N__14574));
    LocalMux I__2895 (
            .O(N__14580),
            .I(N__14574));
    InMux I__2894 (
            .O(N__14579),
            .I(N__14571));
    Odrv4 I__2893 (
            .O(N__14574),
            .I(\c0.d_4_11 ));
    LocalMux I__2892 (
            .O(N__14571),
            .I(\c0.d_4_11 ));
    InMux I__2891 (
            .O(N__14566),
            .I(N__14563));
    LocalMux I__2890 (
            .O(N__14563),
            .I(\c0.tx2_data_RNO_4Z0Z_3 ));
    CascadeMux I__2889 (
            .O(N__14560),
            .I(\c0.tx2_data_RNO_3Z0Z_3_cascade_ ));
    InMux I__2888 (
            .O(N__14557),
            .I(N__14554));
    LocalMux I__2887 (
            .O(N__14554),
            .I(\c0.tx2_data_RNO_0Z0Z_3 ));
    CascadeMux I__2886 (
            .O(N__14551),
            .I(\c0.m105_ns_1_cascade_ ));
    InMux I__2885 (
            .O(N__14548),
            .I(N__14545));
    LocalMux I__2884 (
            .O(N__14545),
            .I(N__14542));
    Span4Mux_h I__2883 (
            .O(N__14542),
            .I(N__14539));
    Odrv4 I__2882 (
            .O(N__14539),
            .I(\c0.tx2_data_RNO_1Z0Z_3 ));
    InMux I__2881 (
            .O(N__14536),
            .I(N__14533));
    LocalMux I__2880 (
            .O(N__14533),
            .I(\c0.tx2.r_Tx_DataZ0Z_3 ));
    CascadeMux I__2879 (
            .O(N__14530),
            .I(N__14527));
    InMux I__2878 (
            .O(N__14527),
            .I(N__14524));
    LocalMux I__2877 (
            .O(N__14524),
            .I(N__14521));
    Span4Mux_v I__2876 (
            .O(N__14521),
            .I(N__14518));
    Odrv4 I__2875 (
            .O(N__14518),
            .I(\c0.tx2_data_RNO_1Z0Z_7 ));
    InMux I__2874 (
            .O(N__14515),
            .I(N__14512));
    LocalMux I__2873 (
            .O(N__14512),
            .I(\c0.m60_0_ns_1 ));
    InMux I__2872 (
            .O(N__14509),
            .I(N__14506));
    LocalMux I__2871 (
            .O(N__14506),
            .I(\c0.tx2.r_Tx_DataZ0Z_7 ));
    InMux I__2870 (
            .O(N__14503),
            .I(N__14499));
    InMux I__2869 (
            .O(N__14502),
            .I(N__14494));
    LocalMux I__2868 (
            .O(N__14499),
            .I(N__14491));
    InMux I__2867 (
            .O(N__14498),
            .I(N__14488));
    InMux I__2866 (
            .O(N__14497),
            .I(N__14485));
    LocalMux I__2865 (
            .O(N__14494),
            .I(N__14482));
    Span12Mux_v I__2864 (
            .O(N__14491),
            .I(N__14475));
    LocalMux I__2863 (
            .O(N__14488),
            .I(N__14475));
    LocalMux I__2862 (
            .O(N__14485),
            .I(N__14475));
    Odrv4 I__2861 (
            .O(N__14482),
            .I(\c0.d_2_6 ));
    Odrv12 I__2860 (
            .O(N__14475),
            .I(\c0.d_2_6 ));
    InMux I__2859 (
            .O(N__14470),
            .I(N__14467));
    LocalMux I__2858 (
            .O(N__14467),
            .I(N__14461));
    InMux I__2857 (
            .O(N__14466),
            .I(N__14456));
    InMux I__2856 (
            .O(N__14465),
            .I(N__14456));
    CascadeMux I__2855 (
            .O(N__14464),
            .I(N__14453));
    Span4Mux_h I__2854 (
            .O(N__14461),
            .I(N__14448));
    LocalMux I__2853 (
            .O(N__14456),
            .I(N__14448));
    InMux I__2852 (
            .O(N__14453),
            .I(N__14445));
    Span4Mux_h I__2851 (
            .O(N__14448),
            .I(N__14442));
    LocalMux I__2850 (
            .O(N__14445),
            .I(\c0.d_2_22 ));
    Odrv4 I__2849 (
            .O(N__14442),
            .I(\c0.d_2_22 ));
    InMux I__2848 (
            .O(N__14437),
            .I(N__14434));
    LocalMux I__2847 (
            .O(N__14434),
            .I(N__14431));
    Span4Mux_h I__2846 (
            .O(N__14431),
            .I(N__14427));
    InMux I__2845 (
            .O(N__14430),
            .I(N__14424));
    Odrv4 I__2844 (
            .O(N__14427),
            .I(\c0.data_in_0_Z0Z_2 ));
    LocalMux I__2843 (
            .O(N__14424),
            .I(\c0.data_in_0_Z0Z_2 ));
    InMux I__2842 (
            .O(N__14419),
            .I(N__14416));
    LocalMux I__2841 (
            .O(N__14416),
            .I(N__14413));
    Span4Mux_h I__2840 (
            .O(N__14413),
            .I(N__14410));
    Span4Mux_v I__2839 (
            .O(N__14410),
            .I(N__14406));
    InMux I__2838 (
            .O(N__14409),
            .I(N__14403));
    Odrv4 I__2837 (
            .O(N__14406),
            .I(\c0.data_in_4_Z0Z_0 ));
    LocalMux I__2836 (
            .O(N__14403),
            .I(\c0.data_in_4_Z0Z_0 ));
    InMux I__2835 (
            .O(N__14398),
            .I(N__14395));
    LocalMux I__2834 (
            .O(N__14395),
            .I(N__14391));
    CascadeMux I__2833 (
            .O(N__14394),
            .I(N__14387));
    Span4Mux_h I__2832 (
            .O(N__14391),
            .I(N__14384));
    InMux I__2831 (
            .O(N__14390),
            .I(N__14379));
    InMux I__2830 (
            .O(N__14387),
            .I(N__14379));
    Odrv4 I__2829 (
            .O(N__14384),
            .I(\c0.d_4_23 ));
    LocalMux I__2828 (
            .O(N__14379),
            .I(\c0.d_4_23 ));
    CascadeMux I__2827 (
            .O(N__14374),
            .I(N__14371));
    InMux I__2826 (
            .O(N__14371),
            .I(N__14368));
    LocalMux I__2825 (
            .O(N__14368),
            .I(\c0.tx2_data_RNO_4Z0Z_7 ));
    InMux I__2824 (
            .O(N__14365),
            .I(N__14362));
    LocalMux I__2823 (
            .O(N__14362),
            .I(N__14357));
    InMux I__2822 (
            .O(N__14361),
            .I(N__14352));
    InMux I__2821 (
            .O(N__14360),
            .I(N__14352));
    Odrv4 I__2820 (
            .O(N__14357),
            .I(\c0.d_4_2 ));
    LocalMux I__2819 (
            .O(N__14352),
            .I(\c0.d_4_2 ));
    InMux I__2818 (
            .O(N__14347),
            .I(N__14344));
    LocalMux I__2817 (
            .O(N__14344),
            .I(N__14341));
    Odrv4 I__2816 (
            .O(N__14341),
            .I(\c0.tx2_data_RNO_4Z0Z_2 ));
    CascadeMux I__2815 (
            .O(N__14338),
            .I(\c0.tx2_data_RNO_3Z0Z_2_cascade_ ));
    InMux I__2814 (
            .O(N__14335),
            .I(N__14332));
    LocalMux I__2813 (
            .O(N__14332),
            .I(N__14329));
    Span4Mux_h I__2812 (
            .O(N__14329),
            .I(N__14326));
    Odrv4 I__2811 (
            .O(N__14326),
            .I(\c0.m131_ns_1 ));
    InMux I__2810 (
            .O(N__14323),
            .I(N__14320));
    LocalMux I__2809 (
            .O(N__14320),
            .I(N__14317));
    Span4Mux_v I__2808 (
            .O(N__14317),
            .I(N__14314));
    Odrv4 I__2807 (
            .O(N__14314),
            .I(\c0.tx_data_RNO_1Z0Z_6 ));
    InMux I__2806 (
            .O(N__14311),
            .I(N__14308));
    LocalMux I__2805 (
            .O(N__14308),
            .I(\c0.tx_data_RNO_0Z0Z_6 ));
    InMux I__2804 (
            .O(N__14305),
            .I(N__14302));
    LocalMux I__2803 (
            .O(N__14302),
            .I(\c0.tx_data_1_0_i_ns_1_6 ));
    InMux I__2802 (
            .O(N__14299),
            .I(N__14296));
    LocalMux I__2801 (
            .O(N__14296),
            .I(N__14293));
    Span4Mux_v I__2800 (
            .O(N__14293),
            .I(N__14290));
    Odrv4 I__2799 (
            .O(N__14290),
            .I(\c0.tx.r_Tx_DataZ0Z_6 ));
    CEMux I__2798 (
            .O(N__14287),
            .I(N__14284));
    LocalMux I__2797 (
            .O(N__14284),
            .I(N__14280));
    CEMux I__2796 (
            .O(N__14283),
            .I(N__14276));
    Span4Mux_v I__2795 (
            .O(N__14280),
            .I(N__14273));
    CEMux I__2794 (
            .O(N__14279),
            .I(N__14270));
    LocalMux I__2793 (
            .O(N__14276),
            .I(N__14267));
    Span4Mux_h I__2792 (
            .O(N__14273),
            .I(N__14262));
    LocalMux I__2791 (
            .O(N__14270),
            .I(N__14262));
    Span4Mux_h I__2790 (
            .O(N__14267),
            .I(N__14259));
    Span4Mux_h I__2789 (
            .O(N__14262),
            .I(N__14256));
    Odrv4 I__2788 (
            .O(N__14259),
            .I(\c0.tx.N_398_i ));
    Odrv4 I__2787 (
            .O(N__14256),
            .I(\c0.tx.N_398_i ));
    CascadeMux I__2786 (
            .O(N__14251),
            .I(N__14248));
    InMux I__2785 (
            .O(N__14248),
            .I(N__14241));
    InMux I__2784 (
            .O(N__14247),
            .I(N__14238));
    CascadeMux I__2783 (
            .O(N__14246),
            .I(N__14234));
    InMux I__2782 (
            .O(N__14245),
            .I(N__14228));
    InMux I__2781 (
            .O(N__14244),
            .I(N__14228));
    LocalMux I__2780 (
            .O(N__14241),
            .I(N__14222));
    LocalMux I__2779 (
            .O(N__14238),
            .I(N__14222));
    CascadeMux I__2778 (
            .O(N__14237),
            .I(N__14218));
    InMux I__2777 (
            .O(N__14234),
            .I(N__14212));
    InMux I__2776 (
            .O(N__14233),
            .I(N__14212));
    LocalMux I__2775 (
            .O(N__14228),
            .I(N__14209));
    InMux I__2774 (
            .O(N__14227),
            .I(N__14206));
    Span12Mux_h I__2773 (
            .O(N__14222),
            .I(N__14203));
    InMux I__2772 (
            .O(N__14221),
            .I(N__14196));
    InMux I__2771 (
            .O(N__14218),
            .I(N__14196));
    InMux I__2770 (
            .O(N__14217),
            .I(N__14196));
    LocalMux I__2769 (
            .O(N__14212),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    Odrv4 I__2768 (
            .O(N__14209),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    LocalMux I__2767 (
            .O(N__14206),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    Odrv12 I__2766 (
            .O(N__14203),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    LocalMux I__2765 (
            .O(N__14196),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    InMux I__2764 (
            .O(N__14185),
            .I(N__14181));
    InMux I__2763 (
            .O(N__14184),
            .I(N__14170));
    LocalMux I__2762 (
            .O(N__14181),
            .I(N__14167));
    InMux I__2761 (
            .O(N__14180),
            .I(N__14164));
    InMux I__2760 (
            .O(N__14179),
            .I(N__14161));
    InMux I__2759 (
            .O(N__14178),
            .I(N__14158));
    InMux I__2758 (
            .O(N__14177),
            .I(N__14153));
    InMux I__2757 (
            .O(N__14176),
            .I(N__14153));
    InMux I__2756 (
            .O(N__14175),
            .I(N__14150));
    InMux I__2755 (
            .O(N__14174),
            .I(N__14145));
    InMux I__2754 (
            .O(N__14173),
            .I(N__14145));
    LocalMux I__2753 (
            .O(N__14170),
            .I(N__14140));
    Span12Mux_h I__2752 (
            .O(N__14167),
            .I(N__14140));
    LocalMux I__2751 (
            .O(N__14164),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2750 (
            .O(N__14161),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2749 (
            .O(N__14158),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2748 (
            .O(N__14153),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2747 (
            .O(N__14150),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2746 (
            .O(N__14145),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    Odrv12 I__2745 (
            .O(N__14140),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    InMux I__2744 (
            .O(N__14125),
            .I(N__14121));
    InMux I__2743 (
            .O(N__14124),
            .I(N__14118));
    LocalMux I__2742 (
            .O(N__14121),
            .I(N__14113));
    LocalMux I__2741 (
            .O(N__14118),
            .I(N__14106));
    InMux I__2740 (
            .O(N__14117),
            .I(N__14100));
    InMux I__2739 (
            .O(N__14116),
            .I(N__14097));
    Span4Mux_v I__2738 (
            .O(N__14113),
            .I(N__14094));
    InMux I__2737 (
            .O(N__14112),
            .I(N__14091));
    InMux I__2736 (
            .O(N__14111),
            .I(N__14086));
    InMux I__2735 (
            .O(N__14110),
            .I(N__14086));
    InMux I__2734 (
            .O(N__14109),
            .I(N__14083));
    Span12Mux_v I__2733 (
            .O(N__14106),
            .I(N__14080));
    InMux I__2732 (
            .O(N__14105),
            .I(N__14073));
    InMux I__2731 (
            .O(N__14104),
            .I(N__14073));
    InMux I__2730 (
            .O(N__14103),
            .I(N__14073));
    LocalMux I__2729 (
            .O(N__14100),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__2728 (
            .O(N__14097),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    Odrv4 I__2727 (
            .O(N__14094),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__2726 (
            .O(N__14091),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__2725 (
            .O(N__14086),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__2724 (
            .O(N__14083),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    Odrv12 I__2723 (
            .O(N__14080),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__2722 (
            .O(N__14073),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    InMux I__2721 (
            .O(N__14056),
            .I(N__14053));
    LocalMux I__2720 (
            .O(N__14053),
            .I(N__14050));
    Span4Mux_h I__2719 (
            .O(N__14050),
            .I(N__14046));
    InMux I__2718 (
            .O(N__14049),
            .I(N__14043));
    Span4Mux_h I__2717 (
            .O(N__14046),
            .I(N__14040));
    LocalMux I__2716 (
            .O(N__14043),
            .I(N__14037));
    Odrv4 I__2715 (
            .O(N__14040),
            .I(\c0.rx.N_335 ));
    Odrv12 I__2714 (
            .O(N__14037),
            .I(\c0.rx.N_335 ));
    InMux I__2713 (
            .O(N__14032),
            .I(N__14029));
    LocalMux I__2712 (
            .O(N__14029),
            .I(\c0.N_121 ));
    InMux I__2711 (
            .O(N__14026),
            .I(N__14023));
    LocalMux I__2710 (
            .O(N__14023),
            .I(\c0.m163_4 ));
    InMux I__2709 (
            .O(N__14020),
            .I(N__14017));
    LocalMux I__2708 (
            .O(N__14017),
            .I(N__14014));
    Odrv4 I__2707 (
            .O(N__14014),
            .I(\c0.un1_data_in_7__1_0_a2_24_a2_7 ));
    InMux I__2706 (
            .O(N__14011),
            .I(N__14008));
    LocalMux I__2705 (
            .O(N__14008),
            .I(N__14005));
    Odrv4 I__2704 (
            .O(N__14005),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_6 ));
    CascadeMux I__2703 (
            .O(N__14002),
            .I(\c0.m163_8_cascade_ ));
    InMux I__2702 (
            .O(N__13999),
            .I(N__13996));
    LocalMux I__2701 (
            .O(N__13996),
            .I(\c0.un1_data_in_7__1_3 ));
    InMux I__2700 (
            .O(N__13993),
            .I(N__13990));
    LocalMux I__2699 (
            .O(N__13990),
            .I(\c0.m163_10 ));
    CascadeMux I__2698 (
            .O(N__13987),
            .I(\c0.m163_1_cascade_ ));
    InMux I__2697 (
            .O(N__13984),
            .I(N__13981));
    LocalMux I__2696 (
            .O(N__13981),
            .I(\c0.un1_data_in_7__0 ));
    CascadeMux I__2695 (
            .O(N__13978),
            .I(\c0.N_164_0_cascade_ ));
    CascadeMux I__2694 (
            .O(N__13975),
            .I(\c0.N_173_0_cascade_ ));
    InMux I__2693 (
            .O(N__13972),
            .I(N__13969));
    LocalMux I__2692 (
            .O(N__13969),
            .I(N__13966));
    Span4Mux_h I__2691 (
            .O(N__13966),
            .I(N__13961));
    CascadeMux I__2690 (
            .O(N__13965),
            .I(N__13958));
    InMux I__2689 (
            .O(N__13964),
            .I(N__13955));
    Span4Mux_v I__2688 (
            .O(N__13961),
            .I(N__13952));
    InMux I__2687 (
            .O(N__13958),
            .I(N__13949));
    LocalMux I__2686 (
            .O(N__13955),
            .I(\c0.data_in_3_Z0Z_7 ));
    Odrv4 I__2685 (
            .O(N__13952),
            .I(\c0.data_in_3_Z0Z_7 ));
    LocalMux I__2684 (
            .O(N__13949),
            .I(\c0.data_in_3_Z0Z_7 ));
    InMux I__2683 (
            .O(N__13942),
            .I(N__13939));
    LocalMux I__2682 (
            .O(N__13939),
            .I(\c0.d_4_RNIB3JJZ0Z_2 ));
    InMux I__2681 (
            .O(N__13936),
            .I(N__13931));
    InMux I__2680 (
            .O(N__13935),
            .I(N__13928));
    CascadeMux I__2679 (
            .O(N__13934),
            .I(N__13924));
    LocalMux I__2678 (
            .O(N__13931),
            .I(N__13921));
    LocalMux I__2677 (
            .O(N__13928),
            .I(N__13918));
    InMux I__2676 (
            .O(N__13927),
            .I(N__13915));
    InMux I__2675 (
            .O(N__13924),
            .I(N__13912));
    Odrv4 I__2674 (
            .O(N__13921),
            .I(\c0.d_4_44 ));
    Odrv4 I__2673 (
            .O(N__13918),
            .I(\c0.d_4_44 ));
    LocalMux I__2672 (
            .O(N__13915),
            .I(\c0.d_4_44 ));
    LocalMux I__2671 (
            .O(N__13912),
            .I(\c0.d_4_44 ));
    InMux I__2670 (
            .O(N__13903),
            .I(N__13897));
    InMux I__2669 (
            .O(N__13902),
            .I(N__13890));
    InMux I__2668 (
            .O(N__13901),
            .I(N__13890));
    InMux I__2667 (
            .O(N__13900),
            .I(N__13890));
    LocalMux I__2666 (
            .O(N__13897),
            .I(\c0.d_4_36 ));
    LocalMux I__2665 (
            .O(N__13890),
            .I(\c0.d_4_36 ));
    InMux I__2664 (
            .O(N__13885),
            .I(N__13878));
    InMux I__2663 (
            .O(N__13884),
            .I(N__13878));
    InMux I__2662 (
            .O(N__13883),
            .I(N__13875));
    LocalMux I__2661 (
            .O(N__13878),
            .I(\c0.N_104 ));
    LocalMux I__2660 (
            .O(N__13875),
            .I(\c0.N_104 ));
    InMux I__2659 (
            .O(N__13870),
            .I(N__13867));
    LocalMux I__2658 (
            .O(N__13867),
            .I(N__13864));
    Span4Mux_h I__2657 (
            .O(N__13864),
            .I(N__13861));
    Odrv4 I__2656 (
            .O(N__13861),
            .I(\c0.un1_data_in_6__3_0_a2_5_a2_2 ));
    CascadeMux I__2655 (
            .O(N__13858),
            .I(\c0.un1_data_in_6__5_cascade_ ));
    InMux I__2654 (
            .O(N__13855),
            .I(N__13852));
    LocalMux I__2653 (
            .O(N__13852),
            .I(\c0.un1_data_in_6__6 ));
    InMux I__2652 (
            .O(N__13849),
            .I(N__13846));
    LocalMux I__2651 (
            .O(N__13846),
            .I(\c0.un1_data_in_6__1_0_a2_4_a2_2 ));
    CascadeMux I__2650 (
            .O(N__13843),
            .I(\c0.m163_2_cascade_ ));
    InMux I__2649 (
            .O(N__13840),
            .I(N__13837));
    LocalMux I__2648 (
            .O(N__13837),
            .I(N__13834));
    Span4Mux_h I__2647 (
            .O(N__13834),
            .I(N__13830));
    InMux I__2646 (
            .O(N__13833),
            .I(N__13827));
    Odrv4 I__2645 (
            .O(N__13830),
            .I(\c0.N_126 ));
    LocalMux I__2644 (
            .O(N__13827),
            .I(\c0.N_126 ));
    CascadeMux I__2643 (
            .O(N__13822),
            .I(\c0.m163_7_cascade_ ));
    InMux I__2642 (
            .O(N__13819),
            .I(N__13816));
    LocalMux I__2641 (
            .O(N__13816),
            .I(N__13813));
    Odrv4 I__2640 (
            .O(N__13813),
            .I(\c0.m163_0 ));
    CascadeMux I__2639 (
            .O(N__13810),
            .I(N__13807));
    InMux I__2638 (
            .O(N__13807),
            .I(N__13804));
    LocalMux I__2637 (
            .O(N__13804),
            .I(\c0.un1_data_in_6__5_0_a2_5_a2_2 ));
    InMux I__2636 (
            .O(N__13801),
            .I(N__13798));
    LocalMux I__2635 (
            .O(N__13798),
            .I(N__13794));
    InMux I__2634 (
            .O(N__13797),
            .I(N__13790));
    Span4Mux_v I__2633 (
            .O(N__13794),
            .I(N__13787));
    InMux I__2632 (
            .O(N__13793),
            .I(N__13784));
    LocalMux I__2631 (
            .O(N__13790),
            .I(\c0.N_120 ));
    Odrv4 I__2630 (
            .O(N__13787),
            .I(\c0.N_120 ));
    LocalMux I__2629 (
            .O(N__13784),
            .I(\c0.N_120 ));
    InMux I__2628 (
            .O(N__13777),
            .I(N__13774));
    LocalMux I__2627 (
            .O(N__13774),
            .I(N__13770));
    InMux I__2626 (
            .O(N__13773),
            .I(N__13767));
    Span4Mux_h I__2625 (
            .O(N__13770),
            .I(N__13763));
    LocalMux I__2624 (
            .O(N__13767),
            .I(N__13760));
    InMux I__2623 (
            .O(N__13766),
            .I(N__13757));
    Odrv4 I__2622 (
            .O(N__13763),
            .I(\c0.data_in_1_Z0Z_4 ));
    Odrv4 I__2621 (
            .O(N__13760),
            .I(\c0.data_in_1_Z0Z_4 ));
    LocalMux I__2620 (
            .O(N__13757),
            .I(\c0.data_in_1_Z0Z_4 ));
    CascadeMux I__2619 (
            .O(N__13750),
            .I(N__13745));
    InMux I__2618 (
            .O(N__13749),
            .I(N__13740));
    InMux I__2617 (
            .O(N__13748),
            .I(N__13740));
    InMux I__2616 (
            .O(N__13745),
            .I(N__13737));
    LocalMux I__2615 (
            .O(N__13740),
            .I(\c0.d_4_6 ));
    LocalMux I__2614 (
            .O(N__13737),
            .I(\c0.d_4_6 ));
    InMux I__2613 (
            .O(N__13732),
            .I(N__13729));
    LocalMux I__2612 (
            .O(N__13729),
            .I(N__13726));
    Odrv4 I__2611 (
            .O(N__13726),
            .I(\c0.N_109 ));
    InMux I__2610 (
            .O(N__13723),
            .I(N__13720));
    LocalMux I__2609 (
            .O(N__13720),
            .I(N__13717));
    Span4Mux_h I__2608 (
            .O(N__13717),
            .I(N__13713));
    InMux I__2607 (
            .O(N__13716),
            .I(N__13710));
    Span4Mux_h I__2606 (
            .O(N__13713),
            .I(N__13704));
    LocalMux I__2605 (
            .O(N__13710),
            .I(N__13704));
    InMux I__2604 (
            .O(N__13709),
            .I(N__13701));
    Odrv4 I__2603 (
            .O(N__13704),
            .I(\c0.data_in_1_Z0Z_6 ));
    LocalMux I__2602 (
            .O(N__13701),
            .I(\c0.data_in_1_Z0Z_6 ));
    InMux I__2601 (
            .O(N__13696),
            .I(N__13693));
    LocalMux I__2600 (
            .O(N__13693),
            .I(N__13690));
    Span4Mux_v I__2599 (
            .O(N__13690),
            .I(N__13685));
    InMux I__2598 (
            .O(N__13689),
            .I(N__13680));
    InMux I__2597 (
            .O(N__13688),
            .I(N__13680));
    Odrv4 I__2596 (
            .O(N__13685),
            .I(\c0.d_4_7 ));
    LocalMux I__2595 (
            .O(N__13680),
            .I(\c0.d_4_7 ));
    InMux I__2594 (
            .O(N__13675),
            .I(N__13672));
    LocalMux I__2593 (
            .O(N__13672),
            .I(N__13669));
    Span4Mux_v I__2592 (
            .O(N__13669),
            .I(N__13666));
    Odrv4 I__2591 (
            .O(N__13666),
            .I(\c0.tx2_data_RNO_3Z0Z_7 ));
    InMux I__2590 (
            .O(N__13663),
            .I(N__13660));
    LocalMux I__2589 (
            .O(N__13660),
            .I(N__13656));
    InMux I__2588 (
            .O(N__13659),
            .I(N__13653));
    Span4Mux_v I__2587 (
            .O(N__13656),
            .I(N__13650));
    LocalMux I__2586 (
            .O(N__13653),
            .I(N__13647));
    Odrv4 I__2585 (
            .O(N__13650),
            .I(\c0.data_in_4_Z0Z_4 ));
    Odrv4 I__2584 (
            .O(N__13647),
            .I(\c0.data_in_4_Z0Z_4 ));
    InMux I__2583 (
            .O(N__13642),
            .I(N__13637));
    InMux I__2582 (
            .O(N__13641),
            .I(N__13634));
    InMux I__2581 (
            .O(N__13640),
            .I(N__13631));
    LocalMux I__2580 (
            .O(N__13637),
            .I(N__13628));
    LocalMux I__2579 (
            .O(N__13634),
            .I(\c0.data_in_6_Z0Z_1 ));
    LocalMux I__2578 (
            .O(N__13631),
            .I(\c0.data_in_6_Z0Z_1 ));
    Odrv4 I__2577 (
            .O(N__13628),
            .I(\c0.data_in_6_Z0Z_1 ));
    CascadeMux I__2576 (
            .O(N__13621),
            .I(\c0.N_34_cascade_ ));
    InMux I__2575 (
            .O(N__13618),
            .I(N__13614));
    CascadeMux I__2574 (
            .O(N__13617),
            .I(N__13610));
    LocalMux I__2573 (
            .O(N__13614),
            .I(N__13607));
    InMux I__2572 (
            .O(N__13613),
            .I(N__13604));
    InMux I__2571 (
            .O(N__13610),
            .I(N__13601));
    Odrv12 I__2570 (
            .O(N__13607),
            .I(\c0.data_in_2_Z0Z_6 ));
    LocalMux I__2569 (
            .O(N__13604),
            .I(\c0.data_in_2_Z0Z_6 ));
    LocalMux I__2568 (
            .O(N__13601),
            .I(\c0.data_in_2_Z0Z_6 ));
    InMux I__2567 (
            .O(N__13594),
            .I(N__13591));
    LocalMux I__2566 (
            .O(N__13591),
            .I(\c0.byte_transmit_counterZ0Z_5 ));
    InMux I__2565 (
            .O(N__13588),
            .I(N__13585));
    LocalMux I__2564 (
            .O(N__13585),
            .I(N__13580));
    InMux I__2563 (
            .O(N__13584),
            .I(N__13577));
    CascadeMux I__2562 (
            .O(N__13583),
            .I(N__13574));
    Span4Mux_v I__2561 (
            .O(N__13580),
            .I(N__13571));
    LocalMux I__2560 (
            .O(N__13577),
            .I(N__13568));
    InMux I__2559 (
            .O(N__13574),
            .I(N__13565));
    Odrv4 I__2558 (
            .O(N__13571),
            .I(\c0.data_in_6_Z0Z_7 ));
    Odrv4 I__2557 (
            .O(N__13568),
            .I(\c0.data_in_6_Z0Z_7 ));
    LocalMux I__2556 (
            .O(N__13565),
            .I(\c0.data_in_6_Z0Z_7 ));
    InMux I__2555 (
            .O(N__13558),
            .I(N__13555));
    LocalMux I__2554 (
            .O(N__13555),
            .I(\c0.data_in_frame_6_Z0Z_7 ));
    InMux I__2553 (
            .O(N__13552),
            .I(N__13549));
    LocalMux I__2552 (
            .O(N__13549),
            .I(N__13545));
    InMux I__2551 (
            .O(N__13548),
            .I(N__13542));
    Span4Mux_h I__2550 (
            .O(N__13545),
            .I(N__13536));
    LocalMux I__2549 (
            .O(N__13542),
            .I(N__13536));
    CascadeMux I__2548 (
            .O(N__13541),
            .I(N__13533));
    Span4Mux_v I__2547 (
            .O(N__13536),
            .I(N__13530));
    InMux I__2546 (
            .O(N__13533),
            .I(N__13527));
    Odrv4 I__2545 (
            .O(N__13530),
            .I(\c0.data_in_7_Z0Z_7 ));
    LocalMux I__2544 (
            .O(N__13527),
            .I(\c0.data_in_7_Z0Z_7 ));
    CascadeMux I__2543 (
            .O(N__13522),
            .I(N__13519));
    InMux I__2542 (
            .O(N__13519),
            .I(N__13516));
    LocalMux I__2541 (
            .O(N__13516),
            .I(\c0.data_in_frame_7_Z0Z_7 ));
    InMux I__2540 (
            .O(N__13513),
            .I(N__13510));
    LocalMux I__2539 (
            .O(N__13510),
            .I(N__13507));
    Span4Mux_h I__2538 (
            .O(N__13507),
            .I(N__13503));
    CascadeMux I__2537 (
            .O(N__13506),
            .I(N__13500));
    Span4Mux_v I__2536 (
            .O(N__13503),
            .I(N__13497));
    InMux I__2535 (
            .O(N__13500),
            .I(N__13494));
    Odrv4 I__2534 (
            .O(N__13497),
            .I(\c0.data_in_0_Z0Z_6 ));
    LocalMux I__2533 (
            .O(N__13494),
            .I(\c0.data_in_0_Z0Z_6 ));
    InMux I__2532 (
            .O(N__13489),
            .I(N__13486));
    LocalMux I__2531 (
            .O(N__13486),
            .I(N__13481));
    InMux I__2530 (
            .O(N__13485),
            .I(N__13478));
    InMux I__2529 (
            .O(N__13484),
            .I(N__13475));
    Span4Mux_h I__2528 (
            .O(N__13481),
            .I(N__13472));
    LocalMux I__2527 (
            .O(N__13478),
            .I(N__13467));
    LocalMux I__2526 (
            .O(N__13475),
            .I(N__13467));
    Span4Mux_h I__2525 (
            .O(N__13472),
            .I(N__13464));
    Odrv12 I__2524 (
            .O(N__13467),
            .I(\c0.d_2_9 ));
    Odrv4 I__2523 (
            .O(N__13464),
            .I(\c0.d_2_9 ));
    InMux I__2522 (
            .O(N__13459),
            .I(N__13456));
    LocalMux I__2521 (
            .O(N__13456),
            .I(\c0.tx_data_RNO_3Z0Z_1 ));
    CascadeMux I__2520 (
            .O(N__13453),
            .I(N__13449));
    InMux I__2519 (
            .O(N__13452),
            .I(N__13445));
    InMux I__2518 (
            .O(N__13449),
            .I(N__13442));
    CascadeMux I__2517 (
            .O(N__13448),
            .I(N__13438));
    LocalMux I__2516 (
            .O(N__13445),
            .I(N__13433));
    LocalMux I__2515 (
            .O(N__13442),
            .I(N__13433));
    InMux I__2514 (
            .O(N__13441),
            .I(N__13428));
    InMux I__2513 (
            .O(N__13438),
            .I(N__13428));
    Odrv4 I__2512 (
            .O(N__13433),
            .I(\c0.d_2_2 ));
    LocalMux I__2511 (
            .O(N__13428),
            .I(\c0.d_2_2 ));
    CascadeMux I__2510 (
            .O(N__13423),
            .I(\c0.tx_data_RNO_3Z0Z_2_cascade_ ));
    InMux I__2509 (
            .O(N__13420),
            .I(N__13417));
    LocalMux I__2508 (
            .O(N__13417),
            .I(\c0.tx_data_RNO_4Z0Z_2 ));
    InMux I__2507 (
            .O(N__13414),
            .I(N__13411));
    LocalMux I__2506 (
            .O(N__13411),
            .I(\c0.tx_data_1_0_i_ns_1_2 ));
    InMux I__2505 (
            .O(N__13408),
            .I(N__13405));
    LocalMux I__2504 (
            .O(N__13405),
            .I(N__13401));
    InMux I__2503 (
            .O(N__13404),
            .I(N__13396));
    Span4Mux_v I__2502 (
            .O(N__13401),
            .I(N__13392));
    InMux I__2501 (
            .O(N__13400),
            .I(N__13389));
    InMux I__2500 (
            .O(N__13399),
            .I(N__13386));
    LocalMux I__2499 (
            .O(N__13396),
            .I(N__13383));
    InMux I__2498 (
            .O(N__13395),
            .I(N__13380));
    Span4Mux_h I__2497 (
            .O(N__13392),
            .I(N__13375));
    LocalMux I__2496 (
            .O(N__13389),
            .I(N__13375));
    LocalMux I__2495 (
            .O(N__13386),
            .I(\c0.d_2_39 ));
    Odrv4 I__2494 (
            .O(N__13383),
            .I(\c0.d_2_39 ));
    LocalMux I__2493 (
            .O(N__13380),
            .I(\c0.d_2_39 ));
    Odrv4 I__2492 (
            .O(N__13375),
            .I(\c0.d_2_39 ));
    CascadeMux I__2491 (
            .O(N__13366),
            .I(N__13362));
    InMux I__2490 (
            .O(N__13365),
            .I(N__13358));
    InMux I__2489 (
            .O(N__13362),
            .I(N__13355));
    CascadeMux I__2488 (
            .O(N__13361),
            .I(N__13352));
    LocalMux I__2487 (
            .O(N__13358),
            .I(N__13347));
    LocalMux I__2486 (
            .O(N__13355),
            .I(N__13347));
    InMux I__2485 (
            .O(N__13352),
            .I(N__13344));
    Odrv12 I__2484 (
            .O(N__13347),
            .I(\c0.d_2_47 ));
    LocalMux I__2483 (
            .O(N__13344),
            .I(\c0.d_2_47 ));
    InMux I__2482 (
            .O(N__13339),
            .I(N__13336));
    LocalMux I__2481 (
            .O(N__13336),
            .I(N__13333));
    Odrv4 I__2480 (
            .O(N__13333),
            .I(\c0.tx_data_RNO_0Z0Z_7 ));
    InMux I__2479 (
            .O(N__13330),
            .I(N__13324));
    InMux I__2478 (
            .O(N__13329),
            .I(N__13321));
    InMux I__2477 (
            .O(N__13328),
            .I(N__13316));
    InMux I__2476 (
            .O(N__13327),
            .I(N__13316));
    LocalMux I__2475 (
            .O(N__13324),
            .I(N__13313));
    LocalMux I__2474 (
            .O(N__13321),
            .I(N__13308));
    LocalMux I__2473 (
            .O(N__13316),
            .I(N__13308));
    Odrv4 I__2472 (
            .O(N__13313),
            .I(\c0.d_2_36 ));
    Odrv4 I__2471 (
            .O(N__13308),
            .I(\c0.d_2_36 ));
    CascadeMux I__2470 (
            .O(N__13303),
            .I(N__13300));
    InMux I__2469 (
            .O(N__13300),
            .I(N__13297));
    LocalMux I__2468 (
            .O(N__13297),
            .I(N__13294));
    Span4Mux_h I__2467 (
            .O(N__13294),
            .I(N__13290));
    InMux I__2466 (
            .O(N__13293),
            .I(N__13287));
    Odrv4 I__2465 (
            .O(N__13290),
            .I(\c0.d_2_44 ));
    LocalMux I__2464 (
            .O(N__13287),
            .I(\c0.d_2_44 ));
    InMux I__2463 (
            .O(N__13282),
            .I(N__13279));
    LocalMux I__2462 (
            .O(N__13279),
            .I(N__13276));
    Span4Mux_h I__2461 (
            .O(N__13276),
            .I(N__13273));
    Odrv4 I__2460 (
            .O(N__13273),
            .I(\c0.tx_data_RNO_0Z0Z_4 ));
    InMux I__2459 (
            .O(N__13270),
            .I(N__13267));
    LocalMux I__2458 (
            .O(N__13267),
            .I(N__13264));
    Odrv4 I__2457 (
            .O(N__13264),
            .I(\c0.data_out_6_Z0Z_1 ));
    CascadeMux I__2456 (
            .O(N__13261),
            .I(N__13258));
    InMux I__2455 (
            .O(N__13258),
            .I(N__13255));
    LocalMux I__2454 (
            .O(N__13255),
            .I(N__13252));
    Span4Mux_v I__2453 (
            .O(N__13252),
            .I(N__13249));
    Odrv4 I__2452 (
            .O(N__13249),
            .I(\c0.data_out_7_Z0Z_1 ));
    InMux I__2451 (
            .O(N__13246),
            .I(N__13243));
    LocalMux I__2450 (
            .O(N__13243),
            .I(N__13240));
    Odrv4 I__2449 (
            .O(N__13240),
            .I(\c0.tx_data_RNO_1Z0Z_1 ));
    CascadeMux I__2448 (
            .O(N__13237),
            .I(\c0.m2_e_1_cascade_ ));
    InMux I__2447 (
            .O(N__13234),
            .I(N__13231));
    LocalMux I__2446 (
            .O(N__13231),
            .I(\c0.data_out_7_Z0Z_3 ));
    InMux I__2445 (
            .O(N__13228),
            .I(N__13225));
    LocalMux I__2444 (
            .O(N__13225),
            .I(N__13222));
    Odrv4 I__2443 (
            .O(N__13222),
            .I(\c0.data_out_6_Z0Z_3 ));
    CascadeMux I__2442 (
            .O(N__13219),
            .I(\c0.N_132_mux_cascade_ ));
    InMux I__2441 (
            .O(N__13216),
            .I(N__13213));
    LocalMux I__2440 (
            .O(N__13213),
            .I(N__13210));
    Span4Mux_v I__2439 (
            .O(N__13210),
            .I(N__13207));
    Odrv4 I__2438 (
            .O(N__13207),
            .I(\c0.tx_data_RNO_1Z0Z_3 ));
    InMux I__2437 (
            .O(N__13204),
            .I(N__13201));
    LocalMux I__2436 (
            .O(N__13201),
            .I(\c0.tx_data_RNO_4Z0Z_5 ));
    InMux I__2435 (
            .O(N__13198),
            .I(N__13195));
    LocalMux I__2434 (
            .O(N__13195),
            .I(N__13192));
    Span4Mux_h I__2433 (
            .O(N__13192),
            .I(N__13189));
    Odrv4 I__2432 (
            .O(N__13189),
            .I(\c0.tx_data_RNO_1Z0Z_0 ));
    InMux I__2431 (
            .O(N__13186),
            .I(N__13183));
    LocalMux I__2430 (
            .O(N__13183),
            .I(\c0.tx_data_RNO_0Z0Z_0 ));
    InMux I__2429 (
            .O(N__13180),
            .I(N__13177));
    LocalMux I__2428 (
            .O(N__13177),
            .I(\c0.tx_data_1_0_i_ns_1_0 ));
    InMux I__2427 (
            .O(N__13174),
            .I(N__13171));
    LocalMux I__2426 (
            .O(N__13171),
            .I(N__13168));
    Span4Mux_h I__2425 (
            .O(N__13168),
            .I(N__13165));
    Odrv4 I__2424 (
            .O(N__13165),
            .I(\c0.tx.r_Tx_DataZ0Z_0 ));
    InMux I__2423 (
            .O(N__13162),
            .I(N__13159));
    LocalMux I__2422 (
            .O(N__13159),
            .I(\c0.tx_data_RNO_0Z0Z_2 ));
    InMux I__2421 (
            .O(N__13156),
            .I(N__13153));
    LocalMux I__2420 (
            .O(N__13153),
            .I(N__13150));
    Span4Mux_h I__2419 (
            .O(N__13150),
            .I(N__13147));
    Odrv4 I__2418 (
            .O(N__13147),
            .I(\c0.tx.r_Tx_DataZ0Z_2 ));
    CascadeMux I__2417 (
            .O(N__13144),
            .I(N__13141));
    InMux I__2416 (
            .O(N__13141),
            .I(N__13137));
    InMux I__2415 (
            .O(N__13140),
            .I(N__13132));
    LocalMux I__2414 (
            .O(N__13137),
            .I(N__13129));
    InMux I__2413 (
            .O(N__13136),
            .I(N__13124));
    InMux I__2412 (
            .O(N__13135),
            .I(N__13124));
    LocalMux I__2411 (
            .O(N__13132),
            .I(N__13121));
    Span4Mux_v I__2410 (
            .O(N__13129),
            .I(N__13118));
    LocalMux I__2409 (
            .O(N__13124),
            .I(N__13115));
    Odrv4 I__2408 (
            .O(N__13121),
            .I(\c0.d_2_25 ));
    Odrv4 I__2407 (
            .O(N__13118),
            .I(\c0.d_2_25 ));
    Odrv4 I__2406 (
            .O(N__13115),
            .I(\c0.d_2_25 ));
    CascadeMux I__2405 (
            .O(N__13108),
            .I(\c0.tx_data_RNO_4Z0Z_1_cascade_ ));
    InMux I__2404 (
            .O(N__13105),
            .I(N__13102));
    LocalMux I__2403 (
            .O(N__13102),
            .I(\c0.tx_data_RNO_0Z0Z_1 ));
    CascadeMux I__2402 (
            .O(N__13099),
            .I(\c0.tx_data_1_0_i_ns_1_1_cascade_ ));
    InMux I__2401 (
            .O(N__13096),
            .I(N__13093));
    LocalMux I__2400 (
            .O(N__13093),
            .I(N__13090));
    Span4Mux_h I__2399 (
            .O(N__13090),
            .I(N__13087));
    Odrv4 I__2398 (
            .O(N__13087),
            .I(\c0.tx.r_Tx_DataZ0Z_1 ));
    InMux I__2397 (
            .O(N__13084),
            .I(N__13081));
    LocalMux I__2396 (
            .O(N__13081),
            .I(N__13078));
    Span4Mux_v I__2395 (
            .O(N__13078),
            .I(N__13075));
    Odrv4 I__2394 (
            .O(N__13075),
            .I(\c0.data_out_7_Z0Z_2 ));
    InMux I__2393 (
            .O(N__13072),
            .I(N__13069));
    LocalMux I__2392 (
            .O(N__13069),
            .I(N__13066));
    Span4Mux_v I__2391 (
            .O(N__13066),
            .I(N__13063));
    Odrv4 I__2390 (
            .O(N__13063),
            .I(\c0.data_out_6_Z0Z_2 ));
    InMux I__2389 (
            .O(N__13060),
            .I(N__13057));
    LocalMux I__2388 (
            .O(N__13057),
            .I(\c0.tx_data_RNO_1Z0Z_2 ));
    InMux I__2387 (
            .O(N__13054),
            .I(N__13051));
    LocalMux I__2386 (
            .O(N__13051),
            .I(N__13046));
    InMux I__2385 (
            .O(N__13050),
            .I(N__13043));
    InMux I__2384 (
            .O(N__13049),
            .I(N__13040));
    Span4Mux_v I__2383 (
            .O(N__13046),
            .I(N__13032));
    LocalMux I__2382 (
            .O(N__13043),
            .I(N__13032));
    LocalMux I__2381 (
            .O(N__13040),
            .I(N__13032));
    InMux I__2380 (
            .O(N__13039),
            .I(N__13029));
    Span4Mux_h I__2379 (
            .O(N__13032),
            .I(N__13026));
    LocalMux I__2378 (
            .O(N__13029),
            .I(\c0.d_2_1 ));
    Odrv4 I__2377 (
            .O(N__13026),
            .I(\c0.d_2_1 ));
    CascadeMux I__2376 (
            .O(N__13021),
            .I(N__13017));
    InMux I__2375 (
            .O(N__13020),
            .I(N__13014));
    InMux I__2374 (
            .O(N__13017),
            .I(N__13010));
    LocalMux I__2373 (
            .O(N__13014),
            .I(N__13006));
    InMux I__2372 (
            .O(N__13013),
            .I(N__13003));
    LocalMux I__2371 (
            .O(N__13010),
            .I(N__13000));
    InMux I__2370 (
            .O(N__13009),
            .I(N__12997));
    Span4Mux_h I__2369 (
            .O(N__13006),
            .I(N__12988));
    LocalMux I__2368 (
            .O(N__13003),
            .I(N__12988));
    Span4Mux_h I__2367 (
            .O(N__13000),
            .I(N__12988));
    LocalMux I__2366 (
            .O(N__12997),
            .I(N__12988));
    Odrv4 I__2365 (
            .O(N__12988),
            .I(\c0.d_2_37 ));
    InMux I__2364 (
            .O(N__12985),
            .I(N__12981));
    InMux I__2363 (
            .O(N__12984),
            .I(N__12978));
    LocalMux I__2362 (
            .O(N__12981),
            .I(N__12975));
    LocalMux I__2361 (
            .O(N__12978),
            .I(N__12972));
    Span4Mux_v I__2360 (
            .O(N__12975),
            .I(N__12969));
    Span4Mux_v I__2359 (
            .O(N__12972),
            .I(N__12966));
    Odrv4 I__2358 (
            .O(N__12969),
            .I(\c0.d_2_45 ));
    Odrv4 I__2357 (
            .O(N__12966),
            .I(\c0.d_2_45 ));
    InMux I__2356 (
            .O(N__12961),
            .I(N__12958));
    LocalMux I__2355 (
            .O(N__12958),
            .I(\c0.tx_data_RNO_0Z0Z_5 ));
    CascadeMux I__2354 (
            .O(N__12955),
            .I(\c0.tx_data_RNO_3Z0Z_6_cascade_ ));
    InMux I__2353 (
            .O(N__12952),
            .I(N__12949));
    LocalMux I__2352 (
            .O(N__12949),
            .I(\c0.tx_data_RNO_4Z0Z_6 ));
    CascadeMux I__2351 (
            .O(N__12946),
            .I(N__12943));
    InMux I__2350 (
            .O(N__12943),
            .I(N__12938));
    CascadeMux I__2349 (
            .O(N__12942),
            .I(N__12935));
    CascadeMux I__2348 (
            .O(N__12941),
            .I(N__12930));
    LocalMux I__2347 (
            .O(N__12938),
            .I(N__12927));
    InMux I__2346 (
            .O(N__12935),
            .I(N__12924));
    InMux I__2345 (
            .O(N__12934),
            .I(N__12921));
    InMux I__2344 (
            .O(N__12933),
            .I(N__12916));
    InMux I__2343 (
            .O(N__12930),
            .I(N__12916));
    Span4Mux_v I__2342 (
            .O(N__12927),
            .I(N__12913));
    LocalMux I__2341 (
            .O(N__12924),
            .I(N__12908));
    LocalMux I__2340 (
            .O(N__12921),
            .I(N__12908));
    LocalMux I__2339 (
            .O(N__12916),
            .I(N__12905));
    Span4Mux_h I__2338 (
            .O(N__12913),
            .I(N__12902));
    Span4Mux_v I__2337 (
            .O(N__12908),
            .I(N__12899));
    Span4Mux_h I__2336 (
            .O(N__12905),
            .I(N__12896));
    Span4Mux_h I__2335 (
            .O(N__12902),
            .I(N__12893));
    Odrv4 I__2334 (
            .O(N__12899),
            .I(\c0.d_2_42 ));
    Odrv4 I__2333 (
            .O(N__12896),
            .I(\c0.d_2_42 ));
    Odrv4 I__2332 (
            .O(N__12893),
            .I(\c0.d_2_42 ));
    InMux I__2331 (
            .O(N__12886),
            .I(N__12883));
    LocalMux I__2330 (
            .O(N__12883),
            .I(\c0.nextCRC16_3_3_1 ));
    InMux I__2329 (
            .O(N__12880),
            .I(N__12875));
    InMux I__2328 (
            .O(N__12879),
            .I(N__12870));
    InMux I__2327 (
            .O(N__12878),
            .I(N__12870));
    LocalMux I__2326 (
            .O(N__12875),
            .I(N__12865));
    LocalMux I__2325 (
            .O(N__12870),
            .I(N__12865));
    Span4Mux_h I__2324 (
            .O(N__12865),
            .I(N__12861));
    InMux I__2323 (
            .O(N__12864),
            .I(N__12858));
    Odrv4 I__2322 (
            .O(N__12861),
            .I(\c0.d_2_4 ));
    LocalMux I__2321 (
            .O(N__12858),
            .I(\c0.d_2_4 ));
    CascadeMux I__2320 (
            .O(N__12853),
            .I(\c0.nextCRC16_3_3_1_cascade_ ));
    CascadeMux I__2319 (
            .O(N__12850),
            .I(N__12847));
    InMux I__2318 (
            .O(N__12847),
            .I(N__12844));
    LocalMux I__2317 (
            .O(N__12844),
            .I(N__12841));
    Span4Mux_h I__2316 (
            .O(N__12841),
            .I(N__12838));
    Span4Mux_h I__2315 (
            .O(N__12838),
            .I(N__12835));
    Odrv4 I__2314 (
            .O(N__12835),
            .I(\c0.nextCRC16_3_0_a2_1_1 ));
    InMux I__2313 (
            .O(N__12832),
            .I(N__12829));
    LocalMux I__2312 (
            .O(N__12829),
            .I(N__12824));
    InMux I__2311 (
            .O(N__12828),
            .I(N__12821));
    InMux I__2310 (
            .O(N__12827),
            .I(N__12818));
    Odrv4 I__2309 (
            .O(N__12824),
            .I(\c0.d_2_28 ));
    LocalMux I__2308 (
            .O(N__12821),
            .I(\c0.d_2_28 ));
    LocalMux I__2307 (
            .O(N__12818),
            .I(\c0.d_2_28 ));
    InMux I__2306 (
            .O(N__12811),
            .I(N__12807));
    InMux I__2305 (
            .O(N__12810),
            .I(N__12804));
    LocalMux I__2304 (
            .O(N__12807),
            .I(N__12800));
    LocalMux I__2303 (
            .O(N__12804),
            .I(N__12797));
    InMux I__2302 (
            .O(N__12803),
            .I(N__12794));
    Span4Mux_h I__2301 (
            .O(N__12800),
            .I(N__12791));
    Span4Mux_v I__2300 (
            .O(N__12797),
            .I(N__12786));
    LocalMux I__2299 (
            .O(N__12794),
            .I(N__12786));
    Span4Mux_h I__2298 (
            .O(N__12791),
            .I(N__12783));
    Span4Mux_h I__2297 (
            .O(N__12786),
            .I(N__12780));
    Odrv4 I__2296 (
            .O(N__12783),
            .I(\c0.d_2_5 ));
    Odrv4 I__2295 (
            .O(N__12780),
            .I(\c0.d_2_5 ));
    InMux I__2294 (
            .O(N__12775),
            .I(N__12771));
    CascadeMux I__2293 (
            .O(N__12774),
            .I(N__12768));
    LocalMux I__2292 (
            .O(N__12771),
            .I(N__12764));
    InMux I__2291 (
            .O(N__12768),
            .I(N__12759));
    InMux I__2290 (
            .O(N__12767),
            .I(N__12759));
    Odrv12 I__2289 (
            .O(N__12764),
            .I(\c0.d_2_13 ));
    LocalMux I__2288 (
            .O(N__12759),
            .I(\c0.d_2_13 ));
    CascadeMux I__2287 (
            .O(N__12754),
            .I(\c0.tx_data_RNO_3Z0Z_5_cascade_ ));
    InMux I__2286 (
            .O(N__12751),
            .I(N__12748));
    LocalMux I__2285 (
            .O(N__12748),
            .I(\c0.tx_data_1_0_i_ns_1_5 ));
    InMux I__2284 (
            .O(N__12745),
            .I(N__12742));
    LocalMux I__2283 (
            .O(N__12742),
            .I(N__12739));
    Span4Mux_v I__2282 (
            .O(N__12739),
            .I(N__12735));
    InMux I__2281 (
            .O(N__12738),
            .I(N__12732));
    Odrv4 I__2280 (
            .O(N__12735),
            .I(\c0.N_108 ));
    LocalMux I__2279 (
            .O(N__12732),
            .I(\c0.N_108 ));
    CascadeMux I__2278 (
            .O(N__12727),
            .I(\c0.un1_data_in_7__6_0_a2_5_a2_2_cascade_ ));
    InMux I__2277 (
            .O(N__12724),
            .I(N__12721));
    LocalMux I__2276 (
            .O(N__12721),
            .I(\c0.un1_data_in_7__4_0_a2_0_a2_4 ));
    InMux I__2275 (
            .O(N__12718),
            .I(N__12715));
    LocalMux I__2274 (
            .O(N__12715),
            .I(N__12712));
    Span4Mux_h I__2273 (
            .O(N__12712),
            .I(N__12708));
    InMux I__2272 (
            .O(N__12711),
            .I(N__12705));
    Odrv4 I__2271 (
            .O(N__12708),
            .I(\c0.data_in_0_Z0Z_3 ));
    LocalMux I__2270 (
            .O(N__12705),
            .I(\c0.data_in_0_Z0Z_3 ));
    InMux I__2269 (
            .O(N__12700),
            .I(N__12697));
    LocalMux I__2268 (
            .O(N__12697),
            .I(N__12694));
    Span4Mux_h I__2267 (
            .O(N__12694),
            .I(N__12690));
    InMux I__2266 (
            .O(N__12693),
            .I(N__12687));
    Odrv4 I__2265 (
            .O(N__12690),
            .I(\c0.data_in_0_Z0Z_5 ));
    LocalMux I__2264 (
            .O(N__12687),
            .I(\c0.data_in_0_Z0Z_5 ));
    InMux I__2263 (
            .O(N__12682),
            .I(N__12679));
    LocalMux I__2262 (
            .O(N__12679),
            .I(N__12676));
    Span4Mux_v I__2261 (
            .O(N__12676),
            .I(N__12671));
    InMux I__2260 (
            .O(N__12675),
            .I(N__12666));
    InMux I__2259 (
            .O(N__12674),
            .I(N__12666));
    Odrv4 I__2258 (
            .O(N__12671),
            .I(\c0.data_in_2_Z0Z_2 ));
    LocalMux I__2257 (
            .O(N__12666),
            .I(\c0.data_in_2_Z0Z_2 ));
    CascadeMux I__2256 (
            .O(N__12661),
            .I(N__12658));
    InMux I__2255 (
            .O(N__12658),
            .I(N__12653));
    InMux I__2254 (
            .O(N__12657),
            .I(N__12648));
    InMux I__2253 (
            .O(N__12656),
            .I(N__12648));
    LocalMux I__2252 (
            .O(N__12653),
            .I(\c0.d_4_18 ));
    LocalMux I__2251 (
            .O(N__12648),
            .I(\c0.d_4_18 ));
    InMux I__2250 (
            .O(N__12643),
            .I(N__12638));
    InMux I__2249 (
            .O(N__12642),
            .I(N__12632));
    InMux I__2248 (
            .O(N__12641),
            .I(N__12632));
    LocalMux I__2247 (
            .O(N__12638),
            .I(N__12629));
    InMux I__2246 (
            .O(N__12637),
            .I(N__12626));
    LocalMux I__2245 (
            .O(N__12632),
            .I(N__12623));
    Span4Mux_h I__2244 (
            .O(N__12629),
            .I(N__12618));
    LocalMux I__2243 (
            .O(N__12626),
            .I(N__12618));
    Odrv4 I__2242 (
            .O(N__12623),
            .I(\c0.d_2_38 ));
    Odrv4 I__2241 (
            .O(N__12618),
            .I(\c0.d_2_38 ));
    CascadeMux I__2240 (
            .O(N__12613),
            .I(N__12610));
    InMux I__2239 (
            .O(N__12610),
            .I(N__12607));
    LocalMux I__2238 (
            .O(N__12607),
            .I(N__12603));
    InMux I__2237 (
            .O(N__12606),
            .I(N__12599));
    Span4Mux_h I__2236 (
            .O(N__12603),
            .I(N__12596));
    InMux I__2235 (
            .O(N__12602),
            .I(N__12593));
    LocalMux I__2234 (
            .O(N__12599),
            .I(\c0.d_2_46 ));
    Odrv4 I__2233 (
            .O(N__12596),
            .I(\c0.d_2_46 ));
    LocalMux I__2232 (
            .O(N__12593),
            .I(\c0.d_2_46 ));
    InMux I__2231 (
            .O(N__12586),
            .I(N__12583));
    LocalMux I__2230 (
            .O(N__12583),
            .I(N__12580));
    Span4Mux_v I__2229 (
            .O(N__12580),
            .I(N__12577));
    Odrv4 I__2228 (
            .O(N__12577),
            .I(\c0.data_out_6_Z0Z_7 ));
    CascadeMux I__2227 (
            .O(N__12574),
            .I(N__12571));
    InMux I__2226 (
            .O(N__12571),
            .I(N__12568));
    LocalMux I__2225 (
            .O(N__12568),
            .I(N__12565));
    Span12Mux_h I__2224 (
            .O(N__12565),
            .I(N__12562));
    Odrv12 I__2223 (
            .O(N__12562),
            .I(\c0.data_out_7_Z0Z_7 ));
    InMux I__2222 (
            .O(N__12559),
            .I(N__12556));
    LocalMux I__2221 (
            .O(N__12556),
            .I(\c0.tx_data_RNO_1Z0Z_7 ));
    CascadeMux I__2220 (
            .O(N__12553),
            .I(\c0.un1_data_in_7__1_0_a2_24_a2_3_cascade_ ));
    InMux I__2219 (
            .O(N__12550),
            .I(N__12547));
    LocalMux I__2218 (
            .O(N__12547),
            .I(\c0.un1_data_in_7__1_0_a2_24_a2_4 ));
    InMux I__2217 (
            .O(N__12544),
            .I(N__12541));
    LocalMux I__2216 (
            .O(N__12541),
            .I(N__12538));
    Span4Mux_v I__2215 (
            .O(N__12538),
            .I(N__12534));
    InMux I__2214 (
            .O(N__12537),
            .I(N__12531));
    Odrv4 I__2213 (
            .O(N__12534),
            .I(\c0.data_in_5_Z0Z_4 ));
    LocalMux I__2212 (
            .O(N__12531),
            .I(\c0.data_in_5_Z0Z_4 ));
    InMux I__2211 (
            .O(N__12526),
            .I(N__12523));
    LocalMux I__2210 (
            .O(N__12523),
            .I(N__12520));
    Span4Mux_h I__2209 (
            .O(N__12520),
            .I(N__12516));
    InMux I__2208 (
            .O(N__12519),
            .I(N__12513));
    Odrv4 I__2207 (
            .O(N__12516),
            .I(\c0.data_in_5_Z0Z_2 ));
    LocalMux I__2206 (
            .O(N__12513),
            .I(\c0.data_in_5_Z0Z_2 ));
    InMux I__2205 (
            .O(N__12508),
            .I(N__12505));
    LocalMux I__2204 (
            .O(N__12505),
            .I(N__12501));
    CascadeMux I__2203 (
            .O(N__12504),
            .I(N__12497));
    Span4Mux_v I__2202 (
            .O(N__12501),
            .I(N__12494));
    InMux I__2201 (
            .O(N__12500),
            .I(N__12491));
    InMux I__2200 (
            .O(N__12497),
            .I(N__12488));
    Odrv4 I__2199 (
            .O(N__12494),
            .I(\c0.data_in_2_Z0Z_0 ));
    LocalMux I__2198 (
            .O(N__12491),
            .I(\c0.data_in_2_Z0Z_0 ));
    LocalMux I__2197 (
            .O(N__12488),
            .I(\c0.data_in_2_Z0Z_0 ));
    CascadeMux I__2196 (
            .O(N__12481),
            .I(N__12476));
    InMux I__2195 (
            .O(N__12480),
            .I(N__12473));
    InMux I__2194 (
            .O(N__12479),
            .I(N__12469));
    InMux I__2193 (
            .O(N__12476),
            .I(N__12466));
    LocalMux I__2192 (
            .O(N__12473),
            .I(N__12463));
    InMux I__2191 (
            .O(N__12472),
            .I(N__12460));
    LocalMux I__2190 (
            .O(N__12469),
            .I(N__12455));
    LocalMux I__2189 (
            .O(N__12466),
            .I(N__12455));
    Odrv4 I__2188 (
            .O(N__12463),
            .I(\c0.d_4_33 ));
    LocalMux I__2187 (
            .O(N__12460),
            .I(\c0.d_4_33 ));
    Odrv4 I__2186 (
            .O(N__12455),
            .I(\c0.d_4_33 ));
    CascadeMux I__2185 (
            .O(N__12448),
            .I(\c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_ ));
    InMux I__2184 (
            .O(N__12445),
            .I(N__12442));
    LocalMux I__2183 (
            .O(N__12442),
            .I(N__12439));
    Odrv4 I__2182 (
            .O(N__12439),
            .I(\c0.N_124 ));
    CascadeMux I__2181 (
            .O(N__12436),
            .I(\c0.N_124_cascade_ ));
    CascadeMux I__2180 (
            .O(N__12433),
            .I(\c0.un1_data_in_7__0_0_a2_1_a2_5_cascade_ ));
    CascadeMux I__2179 (
            .O(N__12430),
            .I(\c0.N_121_cascade_ ));
    InMux I__2178 (
            .O(N__12427),
            .I(N__12423));
    InMux I__2177 (
            .O(N__12426),
            .I(N__12420));
    LocalMux I__2176 (
            .O(N__12423),
            .I(N__12417));
    LocalMux I__2175 (
            .O(N__12420),
            .I(\c0.N_125 ));
    Odrv4 I__2174 (
            .O(N__12417),
            .I(\c0.N_125 ));
    CascadeMux I__2173 (
            .O(N__12412),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_4_3_cascade_ ));
    InMux I__2172 (
            .O(N__12409),
            .I(N__12406));
    LocalMux I__2171 (
            .O(N__12406),
            .I(\c0.N_136 ));
    CascadeMux I__2170 (
            .O(N__12403),
            .I(\c0.N_136_cascade_ ));
    CascadeMux I__2169 (
            .O(N__12400),
            .I(N__12397));
    InMux I__2168 (
            .O(N__12397),
            .I(N__12394));
    LocalMux I__2167 (
            .O(N__12394),
            .I(N__12391));
    Odrv12 I__2166 (
            .O(N__12391),
            .I(\c0.un1_data_in_7__0_0_a2_1_a2_2 ));
    CascadeMux I__2165 (
            .O(N__12388),
            .I(N__12383));
    InMux I__2164 (
            .O(N__12387),
            .I(N__12380));
    InMux I__2163 (
            .O(N__12386),
            .I(N__12377));
    InMux I__2162 (
            .O(N__12383),
            .I(N__12374));
    LocalMux I__2161 (
            .O(N__12380),
            .I(N__12371));
    LocalMux I__2160 (
            .O(N__12377),
            .I(N__12366));
    LocalMux I__2159 (
            .O(N__12374),
            .I(N__12366));
    Odrv4 I__2158 (
            .O(N__12371),
            .I(\c0.data_in_3_Z0Z_3 ));
    Odrv4 I__2157 (
            .O(N__12366),
            .I(\c0.data_in_3_Z0Z_3 ));
    CascadeMux I__2156 (
            .O(N__12361),
            .I(\c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_ ));
    InMux I__2155 (
            .O(N__12358),
            .I(N__12354));
    InMux I__2154 (
            .O(N__12357),
            .I(N__12351));
    LocalMux I__2153 (
            .O(N__12354),
            .I(N__12348));
    LocalMux I__2152 (
            .O(N__12351),
            .I(N__12344));
    Span4Mux_h I__2151 (
            .O(N__12348),
            .I(N__12341));
    InMux I__2150 (
            .O(N__12347),
            .I(N__12338));
    Odrv12 I__2149 (
            .O(N__12344),
            .I(\c0.data_in_3_Z0Z_4 ));
    Odrv4 I__2148 (
            .O(N__12341),
            .I(\c0.data_in_3_Z0Z_4 ));
    LocalMux I__2147 (
            .O(N__12338),
            .I(\c0.data_in_3_Z0Z_4 ));
    InMux I__2146 (
            .O(N__12331),
            .I(N__12328));
    LocalMux I__2145 (
            .O(N__12328),
            .I(N__12325));
    Span4Mux_h I__2144 (
            .O(N__12325),
            .I(N__12320));
    InMux I__2143 (
            .O(N__12324),
            .I(N__12315));
    InMux I__2142 (
            .O(N__12323),
            .I(N__12315));
    Odrv4 I__2141 (
            .O(N__12320),
            .I(\c0.data_in_1_Z0Z_5 ));
    LocalMux I__2140 (
            .O(N__12315),
            .I(\c0.data_in_1_Z0Z_5 ));
    InMux I__2139 (
            .O(N__12310),
            .I(N__12307));
    LocalMux I__2138 (
            .O(N__12307),
            .I(N__12302));
    InMux I__2137 (
            .O(N__12306),
            .I(N__12297));
    InMux I__2136 (
            .O(N__12305),
            .I(N__12297));
    Odrv12 I__2135 (
            .O(N__12302),
            .I(\c0.data_in_3_Z0Z_2 ));
    LocalMux I__2134 (
            .O(N__12297),
            .I(\c0.data_in_3_Z0Z_2 ));
    InMux I__2133 (
            .O(N__12292),
            .I(N__12289));
    LocalMux I__2132 (
            .O(N__12289),
            .I(N__12285));
    InMux I__2131 (
            .O(N__12288),
            .I(N__12282));
    Odrv4 I__2130 (
            .O(N__12285),
            .I(\c0.data_in_5_Z0Z_1 ));
    LocalMux I__2129 (
            .O(N__12282),
            .I(\c0.data_in_5_Z0Z_1 ));
    InMux I__2128 (
            .O(N__12277),
            .I(N__12274));
    LocalMux I__2127 (
            .O(N__12274),
            .I(N__12271));
    Span4Mux_h I__2126 (
            .O(N__12271),
            .I(N__12267));
    InMux I__2125 (
            .O(N__12270),
            .I(N__12264));
    Odrv4 I__2124 (
            .O(N__12267),
            .I(\c0.data_in_5_Z0Z_0 ));
    LocalMux I__2123 (
            .O(N__12264),
            .I(\c0.data_in_5_Z0Z_0 ));
    InMux I__2122 (
            .O(N__12259),
            .I(N__12255));
    InMux I__2121 (
            .O(N__12258),
            .I(N__12252));
    LocalMux I__2120 (
            .O(N__12255),
            .I(N__12246));
    LocalMux I__2119 (
            .O(N__12252),
            .I(N__12246));
    InMux I__2118 (
            .O(N__12251),
            .I(N__12243));
    Odrv4 I__2117 (
            .O(N__12246),
            .I(\c0.N_132 ));
    LocalMux I__2116 (
            .O(N__12243),
            .I(\c0.N_132 ));
    InMux I__2115 (
            .O(N__12238),
            .I(N__12235));
    LocalMux I__2114 (
            .O(N__12235),
            .I(N__12232));
    Span4Mux_h I__2113 (
            .O(N__12232),
            .I(N__12229));
    Span4Mux_h I__2112 (
            .O(N__12229),
            .I(N__12225));
    InMux I__2111 (
            .O(N__12228),
            .I(N__12222));
    Odrv4 I__2110 (
            .O(N__12225),
            .I(\c0.rx_data_4 ));
    LocalMux I__2109 (
            .O(N__12222),
            .I(\c0.rx_data_4 ));
    InMux I__2108 (
            .O(N__12217),
            .I(N__12214));
    LocalMux I__2107 (
            .O(N__12214),
            .I(N__12211));
    Span12Mux_v I__2106 (
            .O(N__12211),
            .I(N__12207));
    InMux I__2105 (
            .O(N__12210),
            .I(N__12204));
    Odrv12 I__2104 (
            .O(N__12207),
            .I(\c0.rx_data_2 ));
    LocalMux I__2103 (
            .O(N__12204),
            .I(\c0.rx_data_2 ));
    InMux I__2102 (
            .O(N__12199),
            .I(N__12195));
    InMux I__2101 (
            .O(N__12198),
            .I(N__12190));
    LocalMux I__2100 (
            .O(N__12195),
            .I(N__12187));
    InMux I__2099 (
            .O(N__12194),
            .I(N__12184));
    InMux I__2098 (
            .O(N__12193),
            .I(N__12181));
    LocalMux I__2097 (
            .O(N__12190),
            .I(N__12178));
    Odrv12 I__2096 (
            .O(N__12187),
            .I(\c0.d_4_34 ));
    LocalMux I__2095 (
            .O(N__12184),
            .I(\c0.d_4_34 ));
    LocalMux I__2094 (
            .O(N__12181),
            .I(\c0.d_4_34 ));
    Odrv4 I__2093 (
            .O(N__12178),
            .I(\c0.d_4_34 ));
    CascadeMux I__2092 (
            .O(N__12169),
            .I(\c0.un1_data_in_7__7_0_a2_0_a2_2_cascade_ ));
    InMux I__2091 (
            .O(N__12166),
            .I(N__12163));
    LocalMux I__2090 (
            .O(N__12163),
            .I(N__12160));
    Odrv4 I__2089 (
            .O(N__12160),
            .I(\c0.un1_data_in_6__0_0_a2_5_a2_2 ));
    CascadeMux I__2088 (
            .O(N__12157),
            .I(\c0.un1_data_in_7__7_i_cascade_ ));
    InMux I__2087 (
            .O(N__12154),
            .I(N__12151));
    LocalMux I__2086 (
            .O(N__12151),
            .I(N__12147));
    InMux I__2085 (
            .O(N__12150),
            .I(N__12144));
    Odrv4 I__2084 (
            .O(N__12147),
            .I(\c0.data_in_5_Z0Z_7 ));
    LocalMux I__2083 (
            .O(N__12144),
            .I(\c0.data_in_5_Z0Z_7 ));
    InMux I__2082 (
            .O(N__12139),
            .I(N__12135));
    InMux I__2081 (
            .O(N__12138),
            .I(N__12132));
    LocalMux I__2080 (
            .O(N__12135),
            .I(N__12129));
    LocalMux I__2079 (
            .O(N__12132),
            .I(N__12126));
    Odrv4 I__2078 (
            .O(N__12129),
            .I(\c0.data_in_4_Z0Z_3 ));
    Odrv4 I__2077 (
            .O(N__12126),
            .I(\c0.data_in_4_Z0Z_3 ));
    InMux I__2076 (
            .O(N__12121),
            .I(N__12115));
    InMux I__2075 (
            .O(N__12120),
            .I(N__12115));
    LocalMux I__2074 (
            .O(N__12115),
            .I(N__12110));
    InMux I__2073 (
            .O(N__12114),
            .I(N__12107));
    InMux I__2072 (
            .O(N__12113),
            .I(N__12104));
    Span4Mux_h I__2071 (
            .O(N__12110),
            .I(N__12101));
    LocalMux I__2070 (
            .O(N__12107),
            .I(N__12098));
    LocalMux I__2069 (
            .O(N__12104),
            .I(\c0.d_2_32 ));
    Odrv4 I__2068 (
            .O(N__12101),
            .I(\c0.d_2_32 ));
    Odrv4 I__2067 (
            .O(N__12098),
            .I(\c0.d_2_32 ));
    CascadeMux I__2066 (
            .O(N__12091),
            .I(N__12087));
    CascadeMux I__2065 (
            .O(N__12090),
            .I(N__12083));
    InMux I__2064 (
            .O(N__12087),
            .I(N__12079));
    InMux I__2063 (
            .O(N__12086),
            .I(N__12074));
    InMux I__2062 (
            .O(N__12083),
            .I(N__12074));
    CascadeMux I__2061 (
            .O(N__12082),
            .I(N__12071));
    LocalMux I__2060 (
            .O(N__12079),
            .I(N__12068));
    LocalMux I__2059 (
            .O(N__12074),
            .I(N__12065));
    InMux I__2058 (
            .O(N__12071),
            .I(N__12062));
    Span4Mux_h I__2057 (
            .O(N__12068),
            .I(N__12059));
    Span4Mux_v I__2056 (
            .O(N__12065),
            .I(N__12056));
    LocalMux I__2055 (
            .O(N__12062),
            .I(\c0.d_2_24 ));
    Odrv4 I__2054 (
            .O(N__12059),
            .I(\c0.d_2_24 ));
    Odrv4 I__2053 (
            .O(N__12056),
            .I(\c0.d_2_24 ));
    InMux I__2052 (
            .O(N__12049),
            .I(N__12046));
    LocalMux I__2051 (
            .O(N__12046),
            .I(\c0.nextCRC16_3_3_12 ));
    CascadeMux I__2050 (
            .O(N__12043),
            .I(\c0.nextCRC16_3_4_12_cascade_ ));
    InMux I__2049 (
            .O(N__12040),
            .I(N__12037));
    LocalMux I__2048 (
            .O(N__12037),
            .I(N__12032));
    InMux I__2047 (
            .O(N__12036),
            .I(N__12029));
    InMux I__2046 (
            .O(N__12035),
            .I(N__12026));
    Span4Mux_v I__2045 (
            .O(N__12032),
            .I(N__12019));
    LocalMux I__2044 (
            .O(N__12029),
            .I(N__12019));
    LocalMux I__2043 (
            .O(N__12026),
            .I(N__12019));
    Span4Mux_h I__2042 (
            .O(N__12019),
            .I(N__12016));
    Odrv4 I__2041 (
            .O(N__12016),
            .I(\c0.d_2_41 ));
    InMux I__2040 (
            .O(N__12013),
            .I(N__12010));
    LocalMux I__2039 (
            .O(N__12010),
            .I(N__12007));
    Span4Mux_h I__2038 (
            .O(N__12007),
            .I(N__12004));
    Odrv4 I__2037 (
            .O(N__12004),
            .I(\c0.N_94 ));
    CascadeMux I__2036 (
            .O(N__12001),
            .I(\c0.N_94_cascade_ ));
    CascadeMux I__2035 (
            .O(N__11998),
            .I(N__11993));
    CascadeMux I__2034 (
            .O(N__11997),
            .I(N__11989));
    InMux I__2033 (
            .O(N__11996),
            .I(N__11986));
    InMux I__2032 (
            .O(N__11993),
            .I(N__11983));
    InMux I__2031 (
            .O(N__11992),
            .I(N__11980));
    InMux I__2030 (
            .O(N__11989),
            .I(N__11977));
    LocalMux I__2029 (
            .O(N__11986),
            .I(N__11974));
    LocalMux I__2028 (
            .O(N__11983),
            .I(N__11969));
    LocalMux I__2027 (
            .O(N__11980),
            .I(N__11969));
    LocalMux I__2026 (
            .O(N__11977),
            .I(N__11964));
    Span4Mux_v I__2025 (
            .O(N__11974),
            .I(N__11964));
    Odrv12 I__2024 (
            .O(N__11969),
            .I(\c0.d_2_23 ));
    Odrv4 I__2023 (
            .O(N__11964),
            .I(\c0.d_2_23 ));
    CascadeMux I__2022 (
            .O(N__11959),
            .I(N__11956));
    InMux I__2021 (
            .O(N__11956),
            .I(N__11951));
    CascadeMux I__2020 (
            .O(N__11955),
            .I(N__11948));
    InMux I__2019 (
            .O(N__11954),
            .I(N__11944));
    LocalMux I__2018 (
            .O(N__11951),
            .I(N__11941));
    InMux I__2017 (
            .O(N__11948),
            .I(N__11935));
    InMux I__2016 (
            .O(N__11947),
            .I(N__11935));
    LocalMux I__2015 (
            .O(N__11944),
            .I(N__11930));
    Span4Mux_v I__2014 (
            .O(N__11941),
            .I(N__11930));
    InMux I__2013 (
            .O(N__11940),
            .I(N__11927));
    LocalMux I__2012 (
            .O(N__11935),
            .I(N__11924));
    Odrv4 I__2011 (
            .O(N__11930),
            .I(\c0.d_2_40 ));
    LocalMux I__2010 (
            .O(N__11927),
            .I(\c0.d_2_40 ));
    Odrv4 I__2009 (
            .O(N__11924),
            .I(\c0.d_2_40 ));
    InMux I__2008 (
            .O(N__11917),
            .I(N__11914));
    LocalMux I__2007 (
            .O(N__11914),
            .I(\c0.nextCRC16_3_0_a2_1_11 ));
    InMux I__2006 (
            .O(N__11911),
            .I(N__11908));
    LocalMux I__2005 (
            .O(N__11908),
            .I(\c0.data_out_6_Z0Z_4 ));
    CascadeMux I__2004 (
            .O(N__11905),
            .I(N__11902));
    InMux I__2003 (
            .O(N__11902),
            .I(N__11899));
    LocalMux I__2002 (
            .O(N__11899),
            .I(N__11896));
    Span4Mux_v I__2001 (
            .O(N__11896),
            .I(N__11893));
    Odrv4 I__2000 (
            .O(N__11893),
            .I(\c0.data_out_7_Z0Z_4 ));
    InMux I__1999 (
            .O(N__11890),
            .I(N__11887));
    LocalMux I__1998 (
            .O(N__11887),
            .I(N__11884));
    Span4Mux_v I__1997 (
            .O(N__11884),
            .I(N__11881));
    Odrv4 I__1996 (
            .O(N__11881),
            .I(\c0.tx_data_RNO_1Z0Z_4 ));
    InMux I__1995 (
            .O(N__11878),
            .I(N__11874));
    InMux I__1994 (
            .O(N__11877),
            .I(N__11871));
    LocalMux I__1993 (
            .O(N__11874),
            .I(\c0.data_in_5_Z0Z_5 ));
    LocalMux I__1992 (
            .O(N__11871),
            .I(\c0.data_in_5_Z0Z_5 ));
    InMux I__1991 (
            .O(N__11866),
            .I(N__11863));
    LocalMux I__1990 (
            .O(N__11863),
            .I(N__11859));
    InMux I__1989 (
            .O(N__11862),
            .I(N__11856));
    Span4Mux_v I__1988 (
            .O(N__11859),
            .I(N__11851));
    LocalMux I__1987 (
            .O(N__11856),
            .I(N__11851));
    Span4Mux_h I__1986 (
            .O(N__11851),
            .I(N__11848));
    Span4Mux_h I__1985 (
            .O(N__11848),
            .I(N__11845));
    Odrv4 I__1984 (
            .O(N__11845),
            .I(\c0.d_2_8 ));
    CascadeMux I__1983 (
            .O(N__11842),
            .I(N__11839));
    InMux I__1982 (
            .O(N__11839),
            .I(N__11836));
    LocalMux I__1981 (
            .O(N__11836),
            .I(N__11832));
    InMux I__1980 (
            .O(N__11835),
            .I(N__11828));
    Span4Mux_h I__1979 (
            .O(N__11832),
            .I(N__11825));
    InMux I__1978 (
            .O(N__11831),
            .I(N__11821));
    LocalMux I__1977 (
            .O(N__11828),
            .I(N__11816));
    Span4Mux_h I__1976 (
            .O(N__11825),
            .I(N__11816));
    InMux I__1975 (
            .O(N__11824),
            .I(N__11813));
    LocalMux I__1974 (
            .O(N__11821),
            .I(\c0.d_2_0 ));
    Odrv4 I__1973 (
            .O(N__11816),
            .I(\c0.d_2_0 ));
    LocalMux I__1972 (
            .O(N__11813),
            .I(\c0.d_2_0 ));
    CascadeMux I__1971 (
            .O(N__11806),
            .I(\c0.tx_data_RNO_3Z0Z_0_cascade_ ));
    InMux I__1970 (
            .O(N__11803),
            .I(N__11800));
    LocalMux I__1969 (
            .O(N__11800),
            .I(\c0.tx_data_RNO_4Z0Z_0 ));
    InMux I__1968 (
            .O(N__11797),
            .I(N__11791));
    InMux I__1967 (
            .O(N__11796),
            .I(N__11791));
    LocalMux I__1966 (
            .O(N__11791),
            .I(N__11787));
    InMux I__1965 (
            .O(N__11790),
            .I(N__11784));
    Odrv4 I__1964 (
            .O(N__11787),
            .I(\c0.d_2_33 ));
    LocalMux I__1963 (
            .O(N__11784),
            .I(\c0.d_2_33 ));
    CascadeMux I__1962 (
            .O(N__11779),
            .I(N__11775));
    InMux I__1961 (
            .O(N__11778),
            .I(N__11772));
    InMux I__1960 (
            .O(N__11775),
            .I(N__11769));
    LocalMux I__1959 (
            .O(N__11772),
            .I(N__11766));
    LocalMux I__1958 (
            .O(N__11769),
            .I(N__11763));
    Span4Mux_v I__1957 (
            .O(N__11766),
            .I(N__11757));
    Span4Mux_h I__1956 (
            .O(N__11763),
            .I(N__11757));
    InMux I__1955 (
            .O(N__11762),
            .I(N__11754));
    Odrv4 I__1954 (
            .O(N__11757),
            .I(\c0.d_2_34 ));
    LocalMux I__1953 (
            .O(N__11754),
            .I(\c0.d_2_34 ));
    CascadeMux I__1952 (
            .O(N__11749),
            .I(N__11745));
    InMux I__1951 (
            .O(N__11748),
            .I(N__11742));
    InMux I__1950 (
            .O(N__11745),
            .I(N__11737));
    LocalMux I__1949 (
            .O(N__11742),
            .I(N__11734));
    InMux I__1948 (
            .O(N__11741),
            .I(N__11731));
    InMux I__1947 (
            .O(N__11740),
            .I(N__11728));
    LocalMux I__1946 (
            .O(N__11737),
            .I(N__11725));
    Span4Mux_h I__1945 (
            .O(N__11734),
            .I(N__11718));
    LocalMux I__1944 (
            .O(N__11731),
            .I(N__11718));
    LocalMux I__1943 (
            .O(N__11728),
            .I(N__11718));
    Odrv12 I__1942 (
            .O(N__11725),
            .I(\c0.d_2_15 ));
    Odrv4 I__1941 (
            .O(N__11718),
            .I(\c0.d_2_15 ));
    InMux I__1940 (
            .O(N__11713),
            .I(N__11707));
    InMux I__1939 (
            .O(N__11712),
            .I(N__11704));
    InMux I__1938 (
            .O(N__11711),
            .I(N__11699));
    InMux I__1937 (
            .O(N__11710),
            .I(N__11699));
    LocalMux I__1936 (
            .O(N__11707),
            .I(N__11696));
    LocalMux I__1935 (
            .O(N__11704),
            .I(N__11693));
    LocalMux I__1934 (
            .O(N__11699),
            .I(N__11690));
    Span4Mux_h I__1933 (
            .O(N__11696),
            .I(N__11687));
    Span4Mux_h I__1932 (
            .O(N__11693),
            .I(N__11684));
    Span4Mux_h I__1931 (
            .O(N__11690),
            .I(N__11681));
    Odrv4 I__1930 (
            .O(N__11687),
            .I(\c0.d_2_43 ));
    Odrv4 I__1929 (
            .O(N__11684),
            .I(\c0.d_2_43 ));
    Odrv4 I__1928 (
            .O(N__11681),
            .I(\c0.d_2_43 ));
    CascadeMux I__1927 (
            .O(N__11674),
            .I(\c0.un105_newcrc_0_a2_0_cascade_ ));
    InMux I__1926 (
            .O(N__11671),
            .I(N__11668));
    LocalMux I__1925 (
            .O(N__11668),
            .I(N__11663));
    InMux I__1924 (
            .O(N__11667),
            .I(N__11660));
    InMux I__1923 (
            .O(N__11666),
            .I(N__11657));
    Odrv4 I__1922 (
            .O(N__11663),
            .I(\c0.N_100 ));
    LocalMux I__1921 (
            .O(N__11660),
            .I(\c0.N_100 ));
    LocalMux I__1920 (
            .O(N__11657),
            .I(\c0.N_100 ));
    InMux I__1919 (
            .O(N__11650),
            .I(N__11646));
    InMux I__1918 (
            .O(N__11649),
            .I(N__11642));
    LocalMux I__1917 (
            .O(N__11646),
            .I(N__11639));
    InMux I__1916 (
            .O(N__11645),
            .I(N__11635));
    LocalMux I__1915 (
            .O(N__11642),
            .I(N__11630));
    Span4Mux_h I__1914 (
            .O(N__11639),
            .I(N__11630));
    InMux I__1913 (
            .O(N__11638),
            .I(N__11627));
    LocalMux I__1912 (
            .O(N__11635),
            .I(\c0.d_2_31 ));
    Odrv4 I__1911 (
            .O(N__11630),
            .I(\c0.d_2_31 ));
    LocalMux I__1910 (
            .O(N__11627),
            .I(\c0.d_2_31 ));
    InMux I__1909 (
            .O(N__11620),
            .I(N__11617));
    LocalMux I__1908 (
            .O(N__11617),
            .I(\c0.un105_newcrc_0_a2_3 ));
    InMux I__1907 (
            .O(N__11614),
            .I(N__11611));
    LocalMux I__1906 (
            .O(N__11611),
            .I(\c0.tx_data_RNO_1Z0Z_5 ));
    CascadeMux I__1905 (
            .O(N__11608),
            .I(N__11605));
    InMux I__1904 (
            .O(N__11605),
            .I(N__11602));
    LocalMux I__1903 (
            .O(N__11602),
            .I(\c0.tx.r_Tx_DataZ0Z_5 ));
    InMux I__1902 (
            .O(N__11599),
            .I(N__11595));
    InMux I__1901 (
            .O(N__11598),
            .I(N__11592));
    LocalMux I__1900 (
            .O(N__11595),
            .I(N__11589));
    LocalMux I__1899 (
            .O(N__11592),
            .I(N__11585));
    Span4Mux_v I__1898 (
            .O(N__11589),
            .I(N__11582));
    InMux I__1897 (
            .O(N__11588),
            .I(N__11579));
    Odrv4 I__1896 (
            .O(N__11585),
            .I(\c0.N_24_0 ));
    Odrv4 I__1895 (
            .O(N__11582),
            .I(\c0.N_24_0 ));
    LocalMux I__1894 (
            .O(N__11579),
            .I(\c0.N_24_0 ));
    InMux I__1893 (
            .O(N__11572),
            .I(N__11569));
    LocalMux I__1892 (
            .O(N__11569),
            .I(N__11566));
    Odrv4 I__1891 (
            .O(N__11566),
            .I(\c0.un144_newcrc_2 ));
    CascadeMux I__1890 (
            .O(N__11563),
            .I(\c0.un144_newcrc_5_cascade_ ));
    CascadeMux I__1889 (
            .O(N__11560),
            .I(N__11557));
    InMux I__1888 (
            .O(N__11557),
            .I(N__11554));
    LocalMux I__1887 (
            .O(N__11554),
            .I(\c0.data_out_7_Z0Z_6 ));
    InMux I__1886 (
            .O(N__11551),
            .I(N__11548));
    LocalMux I__1885 (
            .O(N__11548),
            .I(\c0.N_81 ));
    InMux I__1884 (
            .O(N__11545),
            .I(N__11542));
    LocalMux I__1883 (
            .O(N__11542),
            .I(\c0.data_out_6_Z0Z_6 ));
    CascadeMux I__1882 (
            .O(N__11539),
            .I(\c0.tx_data_RNO_3Z0Z_4_cascade_ ));
    InMux I__1881 (
            .O(N__11536),
            .I(N__11533));
    LocalMux I__1880 (
            .O(N__11533),
            .I(\c0.tx_data_1_0_i_ns_1_4 ));
    CascadeMux I__1879 (
            .O(N__11530),
            .I(N__11526));
    CascadeMux I__1878 (
            .O(N__11529),
            .I(N__11523));
    InMux I__1877 (
            .O(N__11526),
            .I(N__11518));
    InMux I__1876 (
            .O(N__11523),
            .I(N__11518));
    LocalMux I__1875 (
            .O(N__11518),
            .I(N__11514));
    InMux I__1874 (
            .O(N__11517),
            .I(N__11510));
    Span4Mux_h I__1873 (
            .O(N__11514),
            .I(N__11507));
    InMux I__1872 (
            .O(N__11513),
            .I(N__11504));
    LocalMux I__1871 (
            .O(N__11510),
            .I(\c0.d_2_20 ));
    Odrv4 I__1870 (
            .O(N__11507),
            .I(\c0.d_2_20 ));
    LocalMux I__1869 (
            .O(N__11504),
            .I(\c0.d_2_20 ));
    InMux I__1868 (
            .O(N__11497),
            .I(N__11494));
    LocalMux I__1867 (
            .O(N__11494),
            .I(\c0.tx_data_RNO_4Z0Z_4 ));
    InMux I__1866 (
            .O(N__11491),
            .I(N__11488));
    LocalMux I__1865 (
            .O(N__11488),
            .I(\c0.N_95 ));
    CascadeMux I__1864 (
            .O(N__11485),
            .I(\c0.tx2_data_RNO_0Z0Z_2_cascade_ ));
    InMux I__1863 (
            .O(N__11482),
            .I(N__11479));
    LocalMux I__1862 (
            .O(N__11479),
            .I(N__11476));
    Span4Mux_v I__1861 (
            .O(N__11476),
            .I(N__11473));
    Odrv4 I__1860 (
            .O(N__11473),
            .I(\c0.data_in_frame_6_Z0Z_2 ));
    CascadeMux I__1859 (
            .O(N__11470),
            .I(N__11467));
    InMux I__1858 (
            .O(N__11467),
            .I(N__11464));
    LocalMux I__1857 (
            .O(N__11464),
            .I(N__11461));
    Odrv12 I__1856 (
            .O(N__11461),
            .I(\c0.data_in_frame_7_Z0Z_2 ));
    InMux I__1855 (
            .O(N__11458),
            .I(N__11455));
    LocalMux I__1854 (
            .O(N__11455),
            .I(\c0.tx2_data_RNO_1Z0Z_2 ));
    InMux I__1853 (
            .O(N__11452),
            .I(N__11449));
    LocalMux I__1852 (
            .O(N__11449),
            .I(\c0.tx_data_RNO_0Z0Z_3 ));
    InMux I__1851 (
            .O(N__11446),
            .I(N__11443));
    LocalMux I__1850 (
            .O(N__11443),
            .I(\c0.tx_data_1_0_i_ns_1_3 ));
    InMux I__1849 (
            .O(N__11440),
            .I(N__11437));
    LocalMux I__1848 (
            .O(N__11437),
            .I(N__11434));
    Odrv4 I__1847 (
            .O(N__11434),
            .I(\c0.tx.r_Tx_DataZ0Z_3 ));
    InMux I__1846 (
            .O(N__11431),
            .I(N__11428));
    LocalMux I__1845 (
            .O(N__11428),
            .I(N__11424));
    InMux I__1844 (
            .O(N__11427),
            .I(N__11421));
    Odrv12 I__1843 (
            .O(N__11424),
            .I(\c0.d_2_7 ));
    LocalMux I__1842 (
            .O(N__11421),
            .I(\c0.d_2_7 ));
    CascadeMux I__1841 (
            .O(N__11416),
            .I(\c0.tx_data_RNO_3Z0Z_7_cascade_ ));
    InMux I__1840 (
            .O(N__11413),
            .I(N__11410));
    LocalMux I__1839 (
            .O(N__11410),
            .I(\c0.tx_data_RNO_4Z0Z_7 ));
    CascadeMux I__1838 (
            .O(N__11407),
            .I(\c0.tx_data_1_0_i_ns_1_7_cascade_ ));
    InMux I__1837 (
            .O(N__11404),
            .I(N__11401));
    LocalMux I__1836 (
            .O(N__11401),
            .I(\c0.tx.r_Tx_DataZ0Z_7 ));
    CascadeMux I__1835 (
            .O(N__11398),
            .I(N__11395));
    InMux I__1834 (
            .O(N__11395),
            .I(N__11392));
    LocalMux I__1833 (
            .O(N__11392),
            .I(N__11389));
    Odrv4 I__1832 (
            .O(N__11389),
            .I(\c0.tx.r_Tx_DataZ0Z_4 ));
    InMux I__1831 (
            .O(N__11386),
            .I(N__11382));
    CascadeMux I__1830 (
            .O(N__11385),
            .I(N__11378));
    LocalMux I__1829 (
            .O(N__11382),
            .I(N__11375));
    InMux I__1828 (
            .O(N__11381),
            .I(N__11372));
    InMux I__1827 (
            .O(N__11378),
            .I(N__11369));
    Odrv4 I__1826 (
            .O(N__11375),
            .I(\c0.data_in_7_Z0Z_3 ));
    LocalMux I__1825 (
            .O(N__11372),
            .I(\c0.data_in_7_Z0Z_3 ));
    LocalMux I__1824 (
            .O(N__11369),
            .I(\c0.data_in_7_Z0Z_3 ));
    InMux I__1823 (
            .O(N__11362),
            .I(N__11357));
    InMux I__1822 (
            .O(N__11361),
            .I(N__11354));
    InMux I__1821 (
            .O(N__11360),
            .I(N__11351));
    LocalMux I__1820 (
            .O(N__11357),
            .I(\c0.data_in_2_Z0Z_1 ));
    LocalMux I__1819 (
            .O(N__11354),
            .I(\c0.data_in_2_Z0Z_1 ));
    LocalMux I__1818 (
            .O(N__11351),
            .I(\c0.data_in_2_Z0Z_1 ));
    InMux I__1817 (
            .O(N__11344),
            .I(N__11341));
    LocalMux I__1816 (
            .O(N__11341),
            .I(N__11338));
    Span4Mux_h I__1815 (
            .O(N__11338),
            .I(N__11333));
    InMux I__1814 (
            .O(N__11337),
            .I(N__11328));
    InMux I__1813 (
            .O(N__11336),
            .I(N__11328));
    Odrv4 I__1812 (
            .O(N__11333),
            .I(\c0.data_in_3_Z0Z_6 ));
    LocalMux I__1811 (
            .O(N__11328),
            .I(\c0.data_in_3_Z0Z_6 ));
    CascadeMux I__1810 (
            .O(N__11323),
            .I(N__11320));
    InMux I__1809 (
            .O(N__11320),
            .I(N__11317));
    LocalMux I__1808 (
            .O(N__11317),
            .I(N__11314));
    Odrv4 I__1807 (
            .O(N__11314),
            .I(\c0.data_in_frame_7_Z0Z_3 ));
    InMux I__1806 (
            .O(N__11311),
            .I(N__11307));
    InMux I__1805 (
            .O(N__11310),
            .I(N__11304));
    LocalMux I__1804 (
            .O(N__11307),
            .I(N__11298));
    LocalMux I__1803 (
            .O(N__11304),
            .I(N__11298));
    InMux I__1802 (
            .O(N__11303),
            .I(N__11295));
    Odrv4 I__1801 (
            .O(N__11298),
            .I(\c0.data_in_6_Z0Z_3 ));
    LocalMux I__1800 (
            .O(N__11295),
            .I(\c0.data_in_6_Z0Z_3 ));
    InMux I__1799 (
            .O(N__11290),
            .I(N__11287));
    LocalMux I__1798 (
            .O(N__11287),
            .I(\c0.data_in_frame_6_Z0Z_3 ));
    CascadeMux I__1797 (
            .O(N__11284),
            .I(N__11278));
    InMux I__1796 (
            .O(N__11283),
            .I(N__11273));
    InMux I__1795 (
            .O(N__11282),
            .I(N__11273));
    InMux I__1794 (
            .O(N__11281),
            .I(N__11268));
    InMux I__1793 (
            .O(N__11278),
            .I(N__11268));
    LocalMux I__1792 (
            .O(N__11273),
            .I(\c0.d_4_17 ));
    LocalMux I__1791 (
            .O(N__11268),
            .I(\c0.d_4_17 ));
    CascadeMux I__1790 (
            .O(N__11263),
            .I(N__11260));
    InMux I__1789 (
            .O(N__11260),
            .I(N__11257));
    LocalMux I__1788 (
            .O(N__11257),
            .I(\c0.tx2_data_RNO_4Z0Z_1 ));
    CascadeMux I__1787 (
            .O(N__11254),
            .I(\c0.m161_ns_1_cascade_ ));
    InMux I__1786 (
            .O(N__11251),
            .I(N__11248));
    LocalMux I__1785 (
            .O(N__11248),
            .I(\c0.tx2_data_RNO_0Z0Z_1 ));
    InMux I__1784 (
            .O(N__11245),
            .I(N__11242));
    LocalMux I__1783 (
            .O(N__11242),
            .I(N__11238));
    InMux I__1782 (
            .O(N__11241),
            .I(N__11235));
    Odrv4 I__1781 (
            .O(N__11238),
            .I(\c0.data_in_4_Z0Z_7 ));
    LocalMux I__1780 (
            .O(N__11235),
            .I(\c0.data_in_4_Z0Z_7 ));
    InMux I__1779 (
            .O(N__11230),
            .I(N__11227));
    LocalMux I__1778 (
            .O(N__11227),
            .I(N__11223));
    InMux I__1777 (
            .O(N__11226),
            .I(N__11220));
    Odrv12 I__1776 (
            .O(N__11223),
            .I(\c0.data_in_5_Z0Z_3 ));
    LocalMux I__1775 (
            .O(N__11220),
            .I(\c0.data_in_5_Z0Z_3 ));
    CascadeMux I__1774 (
            .O(N__11215),
            .I(\c0.N_108_cascade_ ));
    CascadeMux I__1773 (
            .O(N__11212),
            .I(\c0.N_122_cascade_ ));
    CascadeMux I__1772 (
            .O(N__11209),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_2_cascade_ ));
    CascadeMux I__1771 (
            .O(N__11206),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_4_cascade_ ));
    InMux I__1770 (
            .O(N__11203),
            .I(N__11200));
    LocalMux I__1769 (
            .O(N__11200),
            .I(N__11197));
    Span4Mux_h I__1768 (
            .O(N__11197),
            .I(N__11192));
    InMux I__1767 (
            .O(N__11196),
            .I(N__11187));
    InMux I__1766 (
            .O(N__11195),
            .I(N__11187));
    Odrv4 I__1765 (
            .O(N__11192),
            .I(\c0.data_in_2_Z0Z_4 ));
    LocalMux I__1764 (
            .O(N__11187),
            .I(\c0.data_in_2_Z0Z_4 ));
    InMux I__1763 (
            .O(N__11182),
            .I(N__11178));
    InMux I__1762 (
            .O(N__11181),
            .I(N__11175));
    LocalMux I__1761 (
            .O(N__11178),
            .I(\c0.data_in_4_Z0Z_2 ));
    LocalMux I__1760 (
            .O(N__11175),
            .I(\c0.data_in_4_Z0Z_2 ));
    InMux I__1759 (
            .O(N__11170),
            .I(N__11167));
    LocalMux I__1758 (
            .O(N__11167),
            .I(N__11163));
    InMux I__1757 (
            .O(N__11166),
            .I(N__11160));
    Span4Mux_h I__1756 (
            .O(N__11163),
            .I(N__11157));
    LocalMux I__1755 (
            .O(N__11160),
            .I(N__11154));
    Odrv4 I__1754 (
            .O(N__11157),
            .I(\c0.data_in_4_Z0Z_5 ));
    Odrv4 I__1753 (
            .O(N__11154),
            .I(\c0.data_in_4_Z0Z_5 ));
    InMux I__1752 (
            .O(N__11149),
            .I(N__11146));
    LocalMux I__1751 (
            .O(N__11146),
            .I(N__11143));
    Span4Mux_h I__1750 (
            .O(N__11143),
            .I(N__11139));
    InMux I__1749 (
            .O(N__11142),
            .I(N__11136));
    Odrv4 I__1748 (
            .O(N__11139),
            .I(\c0.data_in_0_Z0Z_0 ));
    LocalMux I__1747 (
            .O(N__11136),
            .I(\c0.data_in_0_Z0Z_0 ));
    InMux I__1746 (
            .O(N__11131),
            .I(N__11128));
    LocalMux I__1745 (
            .O(N__11128),
            .I(N__11124));
    CascadeMux I__1744 (
            .O(N__11127),
            .I(N__11120));
    Span4Mux_h I__1743 (
            .O(N__11124),
            .I(N__11117));
    InMux I__1742 (
            .O(N__11123),
            .I(N__11114));
    InMux I__1741 (
            .O(N__11120),
            .I(N__11111));
    Odrv4 I__1740 (
            .O(N__11117),
            .I(\c0.data_in_1_Z0Z_3 ));
    LocalMux I__1739 (
            .O(N__11114),
            .I(\c0.data_in_1_Z0Z_3 ));
    LocalMux I__1738 (
            .O(N__11111),
            .I(\c0.data_in_1_Z0Z_3 ));
    InMux I__1737 (
            .O(N__11104),
            .I(N__11101));
    LocalMux I__1736 (
            .O(N__11101),
            .I(N__11096));
    InMux I__1735 (
            .O(N__11100),
            .I(N__11093));
    InMux I__1734 (
            .O(N__11099),
            .I(N__11090));
    Odrv4 I__1733 (
            .O(N__11096),
            .I(\c0.data_in_1_Z0Z_7 ));
    LocalMux I__1732 (
            .O(N__11093),
            .I(\c0.data_in_1_Z0Z_7 ));
    LocalMux I__1731 (
            .O(N__11090),
            .I(\c0.data_in_1_Z0Z_7 ));
    InMux I__1730 (
            .O(N__11083),
            .I(N__11080));
    LocalMux I__1729 (
            .O(N__11080),
            .I(N__11076));
    InMux I__1728 (
            .O(N__11079),
            .I(N__11073));
    Span4Mux_h I__1727 (
            .O(N__11076),
            .I(N__11069));
    LocalMux I__1726 (
            .O(N__11073),
            .I(N__11066));
    InMux I__1725 (
            .O(N__11072),
            .I(N__11063));
    Odrv4 I__1724 (
            .O(N__11069),
            .I(\c0.data_in_3_Z0Z_0 ));
    Odrv4 I__1723 (
            .O(N__11066),
            .I(\c0.data_in_3_Z0Z_0 ));
    LocalMux I__1722 (
            .O(N__11063),
            .I(\c0.data_in_3_Z0Z_0 ));
    InMux I__1721 (
            .O(N__11056),
            .I(N__11053));
    LocalMux I__1720 (
            .O(N__11053),
            .I(N__11050));
    Span4Mux_h I__1719 (
            .O(N__11050),
            .I(N__11045));
    InMux I__1718 (
            .O(N__11049),
            .I(N__11042));
    InMux I__1717 (
            .O(N__11048),
            .I(N__11039));
    Odrv4 I__1716 (
            .O(N__11045),
            .I(\c0.data_in_3_Z0Z_5 ));
    LocalMux I__1715 (
            .O(N__11042),
            .I(\c0.data_in_3_Z0Z_5 ));
    LocalMux I__1714 (
            .O(N__11039),
            .I(\c0.data_in_3_Z0Z_5 ));
    InMux I__1713 (
            .O(N__11032),
            .I(N__11028));
    InMux I__1712 (
            .O(N__11031),
            .I(N__11025));
    LocalMux I__1711 (
            .O(N__11028),
            .I(\c0.data_in_4_Z0Z_1 ));
    LocalMux I__1710 (
            .O(N__11025),
            .I(\c0.data_in_4_Z0Z_1 ));
    InMux I__1709 (
            .O(N__11020),
            .I(N__11017));
    LocalMux I__1708 (
            .O(N__11017),
            .I(N__11014));
    Span4Mux_h I__1707 (
            .O(N__11014),
            .I(N__11009));
    InMux I__1706 (
            .O(N__11013),
            .I(N__11006));
    InMux I__1705 (
            .O(N__11012),
            .I(N__11003));
    Odrv4 I__1704 (
            .O(N__11009),
            .I(\c0.data_in_2_Z0Z_5 ));
    LocalMux I__1703 (
            .O(N__11006),
            .I(\c0.data_in_2_Z0Z_5 ));
    LocalMux I__1702 (
            .O(N__11003),
            .I(\c0.data_in_2_Z0Z_5 ));
    InMux I__1701 (
            .O(N__10996),
            .I(N__10993));
    LocalMux I__1700 (
            .O(N__10993),
            .I(N__10988));
    InMux I__1699 (
            .O(N__10992),
            .I(N__10985));
    InMux I__1698 (
            .O(N__10991),
            .I(N__10982));
    Odrv4 I__1697 (
            .O(N__10988),
            .I(\c0.data_in_2_Z0Z_3 ));
    LocalMux I__1696 (
            .O(N__10985),
            .I(\c0.data_in_2_Z0Z_3 ));
    LocalMux I__1695 (
            .O(N__10982),
            .I(\c0.data_in_2_Z0Z_3 ));
    InMux I__1694 (
            .O(N__10975),
            .I(N__10972));
    LocalMux I__1693 (
            .O(N__10972),
            .I(N__10969));
    Span4Mux_h I__1692 (
            .O(N__10969),
            .I(N__10965));
    InMux I__1691 (
            .O(N__10968),
            .I(N__10962));
    Odrv4 I__1690 (
            .O(N__10965),
            .I(\c0.data_in_0_Z0Z_7 ));
    LocalMux I__1689 (
            .O(N__10962),
            .I(\c0.data_in_0_Z0Z_7 ));
    InMux I__1688 (
            .O(N__10957),
            .I(N__10953));
    CascadeMux I__1687 (
            .O(N__10956),
            .I(N__10949));
    LocalMux I__1686 (
            .O(N__10953),
            .I(N__10946));
    InMux I__1685 (
            .O(N__10952),
            .I(N__10943));
    InMux I__1684 (
            .O(N__10949),
            .I(N__10940));
    Odrv4 I__1683 (
            .O(N__10946),
            .I(\c0.data_in_2_Z0Z_7 ));
    LocalMux I__1682 (
            .O(N__10943),
            .I(\c0.data_in_2_Z0Z_7 ));
    LocalMux I__1681 (
            .O(N__10940),
            .I(\c0.data_in_2_Z0Z_7 ));
    CascadeMux I__1680 (
            .O(N__10933),
            .I(N__10928));
    InMux I__1679 (
            .O(N__10932),
            .I(N__10925));
    InMux I__1678 (
            .O(N__10931),
            .I(N__10922));
    InMux I__1677 (
            .O(N__10928),
            .I(N__10919));
    LocalMux I__1676 (
            .O(N__10925),
            .I(\c0.data_in_6_Z0Z_0 ));
    LocalMux I__1675 (
            .O(N__10922),
            .I(\c0.data_in_6_Z0Z_0 ));
    LocalMux I__1674 (
            .O(N__10919),
            .I(\c0.data_in_6_Z0Z_0 ));
    CascadeMux I__1673 (
            .O(N__10912),
            .I(\c0.N_75_cascade_ ));
    CascadeMux I__1672 (
            .O(N__10909),
            .I(N__10906));
    InMux I__1671 (
            .O(N__10906),
            .I(N__10903));
    LocalMux I__1670 (
            .O(N__10903),
            .I(\c0.N_93 ));
    InMux I__1669 (
            .O(N__10900),
            .I(N__10897));
    LocalMux I__1668 (
            .O(N__10897),
            .I(N__10891));
    InMux I__1667 (
            .O(N__10896),
            .I(N__10888));
    InMux I__1666 (
            .O(N__10895),
            .I(N__10885));
    InMux I__1665 (
            .O(N__10894),
            .I(N__10882));
    Span4Mux_h I__1664 (
            .O(N__10891),
            .I(N__10875));
    LocalMux I__1663 (
            .O(N__10888),
            .I(N__10875));
    LocalMux I__1662 (
            .O(N__10885),
            .I(N__10875));
    LocalMux I__1661 (
            .O(N__10882),
            .I(\c0.d_2_35 ));
    Odrv4 I__1660 (
            .O(N__10875),
            .I(\c0.d_2_35 ));
    InMux I__1659 (
            .O(N__10870),
            .I(N__10867));
    LocalMux I__1658 (
            .O(N__10867),
            .I(N__10863));
    CascadeMux I__1657 (
            .O(N__10866),
            .I(N__10860));
    Span12Mux_v I__1656 (
            .O(N__10863),
            .I(N__10857));
    InMux I__1655 (
            .O(N__10860),
            .I(N__10854));
    Odrv12 I__1654 (
            .O(N__10857),
            .I(\c0.rx_data_7 ));
    LocalMux I__1653 (
            .O(N__10854),
            .I(\c0.rx_data_7 ));
    CascadeMux I__1652 (
            .O(N__10849),
            .I(\c0.N_105_cascade_ ));
    InMux I__1651 (
            .O(N__10846),
            .I(N__10843));
    LocalMux I__1650 (
            .O(N__10843),
            .I(N__10840));
    Odrv4 I__1649 (
            .O(N__10840),
            .I(\c0.data_out_6_Z0Z_5 ));
    CascadeMux I__1648 (
            .O(N__10837),
            .I(\c0.nextCRC16_3_0_a2_1_15_cascade_ ));
    InMux I__1647 (
            .O(N__10834),
            .I(N__10830));
    InMux I__1646 (
            .O(N__10833),
            .I(N__10827));
    LocalMux I__1645 (
            .O(N__10830),
            .I(\c0.N_99 ));
    LocalMux I__1644 (
            .O(N__10827),
            .I(\c0.N_99 ));
    InMux I__1643 (
            .O(N__10822),
            .I(N__10819));
    LocalMux I__1642 (
            .O(N__10819),
            .I(\c0.nextCRC16_3_0_a2_5_15 ));
    InMux I__1641 (
            .O(N__10816),
            .I(N__10813));
    LocalMux I__1640 (
            .O(N__10813),
            .I(\c0.nextCRC16_3_0_a2_2_15 ));
    CascadeMux I__1639 (
            .O(N__10810),
            .I(\c0.N_95_cascade_ ));
    InMux I__1638 (
            .O(N__10807),
            .I(N__10804));
    LocalMux I__1637 (
            .O(N__10804),
            .I(N__10799));
    InMux I__1636 (
            .O(N__10803),
            .I(N__10794));
    InMux I__1635 (
            .O(N__10802),
            .I(N__10794));
    Odrv4 I__1634 (
            .O(N__10799),
            .I(\c0.N_85 ));
    LocalMux I__1633 (
            .O(N__10794),
            .I(\c0.N_85 ));
    InMux I__1632 (
            .O(N__10789),
            .I(N__10783));
    InMux I__1631 (
            .O(N__10788),
            .I(N__10783));
    LocalMux I__1630 (
            .O(N__10783),
            .I(\c0.nextCRC16_3_2_1 ));
    InMux I__1629 (
            .O(N__10780),
            .I(N__10777));
    LocalMux I__1628 (
            .O(N__10777),
            .I(N__10773));
    InMux I__1627 (
            .O(N__10776),
            .I(N__10770));
    Odrv12 I__1626 (
            .O(N__10773),
            .I(\c0.d_2_3 ));
    LocalMux I__1625 (
            .O(N__10770),
            .I(\c0.d_2_3 ));
    InMux I__1624 (
            .O(N__10765),
            .I(N__10762));
    LocalMux I__1623 (
            .O(N__10762),
            .I(N__10758));
    InMux I__1622 (
            .O(N__10761),
            .I(N__10755));
    Odrv4 I__1621 (
            .O(N__10758),
            .I(\c0.N_75 ));
    LocalMux I__1620 (
            .O(N__10755),
            .I(\c0.N_75 ));
    CascadeMux I__1619 (
            .O(N__10750),
            .I(\c0.nextCRC16_3_0_a2_1_2_cascade_ ));
    InMux I__1618 (
            .O(N__10747),
            .I(N__10744));
    LocalMux I__1617 (
            .O(N__10744),
            .I(N__10741));
    Span4Mux_h I__1616 (
            .O(N__10741),
            .I(N__10737));
    InMux I__1615 (
            .O(N__10740),
            .I(N__10734));
    Odrv4 I__1614 (
            .O(N__10737),
            .I(\c0.dataZ0Z_6 ));
    LocalMux I__1613 (
            .O(N__10734),
            .I(\c0.dataZ0Z_6 ));
    CascadeMux I__1612 (
            .O(N__10729),
            .I(\c0.N_99_cascade_ ));
    InMux I__1611 (
            .O(N__10726),
            .I(N__10723));
    LocalMux I__1610 (
            .O(N__10723),
            .I(\c0.nextCRC16_3_0_a2_0_0 ));
    CascadeMux I__1609 (
            .O(N__10720),
            .I(\c0.nextCRC16_3_0_a2_3_0_cascade_ ));
    InMux I__1608 (
            .O(N__10717),
            .I(N__10714));
    LocalMux I__1607 (
            .O(N__10714),
            .I(\c0.nextCRC16_3_0_a2_4_0 ));
    CascadeMux I__1606 (
            .O(N__10711),
            .I(N__10707));
    InMux I__1605 (
            .O(N__10710),
            .I(N__10704));
    InMux I__1604 (
            .O(N__10707),
            .I(N__10701));
    LocalMux I__1603 (
            .O(N__10704),
            .I(N__10698));
    LocalMux I__1602 (
            .O(N__10701),
            .I(N__10695));
    Span4Mux_h I__1601 (
            .O(N__10698),
            .I(N__10692));
    Span4Mux_h I__1600 (
            .O(N__10695),
            .I(N__10689));
    Span4Mux_h I__1599 (
            .O(N__10692),
            .I(N__10686));
    Span4Mux_h I__1598 (
            .O(N__10689),
            .I(N__10683));
    Odrv4 I__1597 (
            .O(N__10686),
            .I(\c0.d_2_27 ));
    Odrv4 I__1596 (
            .O(N__10683),
            .I(\c0.d_2_27 ));
    CascadeMux I__1595 (
            .O(N__10678),
            .I(\c0.N_81_cascade_ ));
    InMux I__1594 (
            .O(N__10675),
            .I(N__10669));
    InMux I__1593 (
            .O(N__10674),
            .I(N__10669));
    LocalMux I__1592 (
            .O(N__10669),
            .I(\c0.N_105 ));
    SRMux I__1591 (
            .O(N__10666),
            .I(N__10663));
    LocalMux I__1590 (
            .O(N__10663),
            .I(N__10660));
    Span4Mux_h I__1589 (
            .O(N__10660),
            .I(N__10657));
    Odrv4 I__1588 (
            .O(N__10657),
            .I(\c0.tx.N_390_i ));
    InMux I__1587 (
            .O(N__10654),
            .I(N__10642));
    InMux I__1586 (
            .O(N__10653),
            .I(N__10642));
    InMux I__1585 (
            .O(N__10652),
            .I(N__10635));
    InMux I__1584 (
            .O(N__10651),
            .I(N__10635));
    InMux I__1583 (
            .O(N__10650),
            .I(N__10635));
    InMux I__1582 (
            .O(N__10649),
            .I(N__10628));
    InMux I__1581 (
            .O(N__10648),
            .I(N__10628));
    InMux I__1580 (
            .O(N__10647),
            .I(N__10628));
    LocalMux I__1579 (
            .O(N__10642),
            .I(N__10623));
    LocalMux I__1578 (
            .O(N__10635),
            .I(N__10623));
    LocalMux I__1577 (
            .O(N__10628),
            .I(\c0.tx.r_SM_Main_dup_2 ));
    Odrv4 I__1576 (
            .O(N__10623),
            .I(\c0.tx.r_SM_Main_dup_2 ));
    CascadeMux I__1575 (
            .O(N__10618),
            .I(N__10615));
    InMux I__1574 (
            .O(N__10615),
            .I(N__10612));
    LocalMux I__1573 (
            .O(N__10612),
            .I(N__10609));
    Odrv4 I__1572 (
            .O(N__10609),
            .I(\c0.tx.r_SM_Main_recr_i_0_a2_0_2_0_1_3 ));
    InMux I__1571 (
            .O(N__10606),
            .I(N__10596));
    InMux I__1570 (
            .O(N__10605),
            .I(N__10593));
    InMux I__1569 (
            .O(N__10604),
            .I(N__10584));
    InMux I__1568 (
            .O(N__10603),
            .I(N__10584));
    InMux I__1567 (
            .O(N__10602),
            .I(N__10584));
    InMux I__1566 (
            .O(N__10601),
            .I(N__10584));
    InMux I__1565 (
            .O(N__10600),
            .I(N__10579));
    InMux I__1564 (
            .O(N__10599),
            .I(N__10579));
    LocalMux I__1563 (
            .O(N__10596),
            .I(\c0.tx.r_Bit_IndexZ0Z_1 ));
    LocalMux I__1562 (
            .O(N__10593),
            .I(\c0.tx.r_Bit_IndexZ0Z_1 ));
    LocalMux I__1561 (
            .O(N__10584),
            .I(\c0.tx.r_Bit_IndexZ0Z_1 ));
    LocalMux I__1560 (
            .O(N__10579),
            .I(\c0.tx.r_Bit_IndexZ0Z_1 ));
    InMux I__1559 (
            .O(N__10570),
            .I(N__10563));
    InMux I__1558 (
            .O(N__10569),
            .I(N__10556));
    InMux I__1557 (
            .O(N__10568),
            .I(N__10556));
    InMux I__1556 (
            .O(N__10567),
            .I(N__10556));
    InMux I__1555 (
            .O(N__10566),
            .I(N__10553));
    LocalMux I__1554 (
            .O(N__10563),
            .I(\c0.tx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__1553 (
            .O(N__10556),
            .I(\c0.tx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__1552 (
            .O(N__10553),
            .I(\c0.tx.r_Bit_IndexZ0Z_2 ));
    CascadeMux I__1551 (
            .O(N__10546),
            .I(N__10543));
    InMux I__1550 (
            .O(N__10543),
            .I(N__10540));
    LocalMux I__1549 (
            .O(N__10540),
            .I(N__10534));
    InMux I__1548 (
            .O(N__10539),
            .I(N__10531));
    InMux I__1547 (
            .O(N__10538),
            .I(N__10524));
    InMux I__1546 (
            .O(N__10537),
            .I(N__10524));
    Span4Mux_h I__1545 (
            .O(N__10534),
            .I(N__10521));
    LocalMux I__1544 (
            .O(N__10531),
            .I(N__10518));
    InMux I__1543 (
            .O(N__10530),
            .I(N__10513));
    InMux I__1542 (
            .O(N__10529),
            .I(N__10513));
    LocalMux I__1541 (
            .O(N__10524),
            .I(\c0.tx.r_SM_Main_dup_1 ));
    Odrv4 I__1540 (
            .O(N__10521),
            .I(\c0.tx.r_SM_Main_dup_1 ));
    Odrv12 I__1539 (
            .O(N__10518),
            .I(\c0.tx.r_SM_Main_dup_1 ));
    LocalMux I__1538 (
            .O(N__10513),
            .I(\c0.tx.r_SM_Main_dup_1 ));
    CascadeMux I__1537 (
            .O(N__10504),
            .I(N__10499));
    CascadeMux I__1536 (
            .O(N__10503),
            .I(N__10495));
    InMux I__1535 (
            .O(N__10502),
            .I(N__10487));
    InMux I__1534 (
            .O(N__10499),
            .I(N__10487));
    InMux I__1533 (
            .O(N__10498),
            .I(N__10487));
    InMux I__1532 (
            .O(N__10495),
            .I(N__10481));
    InMux I__1531 (
            .O(N__10494),
            .I(N__10481));
    LocalMux I__1530 (
            .O(N__10487),
            .I(N__10478));
    InMux I__1529 (
            .O(N__10486),
            .I(N__10475));
    LocalMux I__1528 (
            .O(N__10481),
            .I(\c0.tx.r_Bit_IndexZ0Z_0 ));
    Odrv4 I__1527 (
            .O(N__10478),
            .I(\c0.tx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__1526 (
            .O(N__10475),
            .I(\c0.tx.r_Bit_IndexZ0Z_0 ));
    InMux I__1525 (
            .O(N__10468),
            .I(N__10465));
    LocalMux I__1524 (
            .O(N__10465),
            .I(N__10462));
    Odrv4 I__1523 (
            .O(N__10462),
            .I(\c0.tx.r_SM_Main_recr_i_i_a2_0_1_2 ));
    InMux I__1522 (
            .O(N__10459),
            .I(N__10456));
    LocalMux I__1521 (
            .O(N__10456),
            .I(\c0.data_out_7_Z0Z_5 ));
    CascadeMux I__1520 (
            .O(N__10453),
            .I(\c0.tx_data_RNO_3Z0Z_3_cascade_ ));
    CascadeMux I__1519 (
            .O(N__10450),
            .I(N__10447));
    InMux I__1518 (
            .O(N__10447),
            .I(N__10441));
    InMux I__1517 (
            .O(N__10446),
            .I(N__10441));
    LocalMux I__1516 (
            .O(N__10441),
            .I(N__10437));
    InMux I__1515 (
            .O(N__10440),
            .I(N__10434));
    Span4Mux_v I__1514 (
            .O(N__10437),
            .I(N__10429));
    LocalMux I__1513 (
            .O(N__10434),
            .I(N__10429));
    Odrv4 I__1512 (
            .O(N__10429),
            .I(\c0.d_2_19 ));
    InMux I__1511 (
            .O(N__10426),
            .I(N__10423));
    LocalMux I__1510 (
            .O(N__10423),
            .I(\c0.tx_data_RNO_4Z0Z_3 ));
    InMux I__1509 (
            .O(N__10420),
            .I(N__10417));
    LocalMux I__1508 (
            .O(N__10417),
            .I(N__10414));
    Span4Mux_h I__1507 (
            .O(N__10414),
            .I(N__10410));
    InMux I__1506 (
            .O(N__10413),
            .I(N__10407));
    Odrv4 I__1505 (
            .O(N__10410),
            .I(\c0.rx_data_0 ));
    LocalMux I__1504 (
            .O(N__10407),
            .I(\c0.rx_data_0 ));
    CascadeMux I__1503 (
            .O(N__10402),
            .I(\c0.tx.o_Tx_Serial_2_3_i_m2_ns_1_cascade_ ));
    InMux I__1502 (
            .O(N__10399),
            .I(N__10394));
    InMux I__1501 (
            .O(N__10398),
            .I(N__10391));
    InMux I__1500 (
            .O(N__10397),
            .I(N__10388));
    LocalMux I__1499 (
            .O(N__10394),
            .I(\c0.tx.N_90_ip_RNI1U1EZ0 ));
    LocalMux I__1498 (
            .O(N__10391),
            .I(\c0.tx.N_90_ip_RNI1U1EZ0 ));
    LocalMux I__1497 (
            .O(N__10388),
            .I(\c0.tx.N_90_ip_RNI1U1EZ0 ));
    CascadeMux I__1496 (
            .O(N__10381),
            .I(\c0.tx.o_Tx_Serial_2_6_i_m2_ns_1_cascade_ ));
    InMux I__1495 (
            .O(N__10378),
            .I(N__10375));
    LocalMux I__1494 (
            .O(N__10375),
            .I(\c0.tx.o_Tx_Serial_RNO_3_0 ));
    CascadeMux I__1493 (
            .O(N__10372),
            .I(\c0.tx.o_Tx_Serial_RNO_2_0_cascade_ ));
    CascadeMux I__1492 (
            .O(N__10369),
            .I(N__10364));
    CascadeMux I__1491 (
            .O(N__10368),
            .I(N__10361));
    CascadeMux I__1490 (
            .O(N__10367),
            .I(N__10357));
    InMux I__1489 (
            .O(N__10364),
            .I(N__10347));
    InMux I__1488 (
            .O(N__10361),
            .I(N__10347));
    InMux I__1487 (
            .O(N__10360),
            .I(N__10347));
    InMux I__1486 (
            .O(N__10357),
            .I(N__10347));
    InMux I__1485 (
            .O(N__10356),
            .I(N__10344));
    LocalMux I__1484 (
            .O(N__10347),
            .I(N__10341));
    LocalMux I__1483 (
            .O(N__10344),
            .I(N__10338));
    Span4Mux_h I__1482 (
            .O(N__10341),
            .I(N__10335));
    Span4Mux_h I__1481 (
            .O(N__10338),
            .I(N__10332));
    Odrv4 I__1480 (
            .O(N__10335),
            .I(\c0.tx.r_SM_Main_RNI522EZ0Z_4 ));
    Odrv4 I__1479 (
            .O(N__10332),
            .I(\c0.tx.r_SM_Main_RNI522EZ0Z_4 ));
    CascadeMux I__1478 (
            .O(N__10327),
            .I(\c0.tx.o_Tx_Serial_RNOZ0Z_1_cascade_ ));
    InMux I__1477 (
            .O(N__10324),
            .I(N__10320));
    InMux I__1476 (
            .O(N__10323),
            .I(N__10313));
    LocalMux I__1475 (
            .O(N__10320),
            .I(N__10310));
    InMux I__1474 (
            .O(N__10319),
            .I(N__10307));
    InMux I__1473 (
            .O(N__10318),
            .I(N__10304));
    InMux I__1472 (
            .O(N__10317),
            .I(N__10299));
    InMux I__1471 (
            .O(N__10316),
            .I(N__10299));
    LocalMux I__1470 (
            .O(N__10313),
            .I(\c0.tx.r_SM_Main_dup_3 ));
    Odrv4 I__1469 (
            .O(N__10310),
            .I(\c0.tx.r_SM_Main_dup_3 ));
    LocalMux I__1468 (
            .O(N__10307),
            .I(\c0.tx.r_SM_Main_dup_3 ));
    LocalMux I__1467 (
            .O(N__10304),
            .I(\c0.tx.r_SM_Main_dup_3 ));
    LocalMux I__1466 (
            .O(N__10299),
            .I(\c0.tx.r_SM_Main_dup_3 ));
    IoInMux I__1465 (
            .O(N__10288),
            .I(N__10285));
    LocalMux I__1464 (
            .O(N__10285),
            .I(N__10282));
    IoSpan4Mux I__1463 (
            .O(N__10282),
            .I(N__10279));
    IoSpan4Mux I__1462 (
            .O(N__10279),
            .I(N__10276));
    Span4Mux_s3_h I__1461 (
            .O(N__10276),
            .I(N__10273));
    Span4Mux_h I__1460 (
            .O(N__10273),
            .I(N__10269));
    InMux I__1459 (
            .O(N__10272),
            .I(N__10266));
    Odrv4 I__1458 (
            .O(N__10269),
            .I(PIN_1_c));
    LocalMux I__1457 (
            .O(N__10266),
            .I(PIN_1_c));
    InMux I__1456 (
            .O(N__10261),
            .I(N__10258));
    LocalMux I__1455 (
            .O(N__10258),
            .I(N__10255));
    Span4Mux_h I__1454 (
            .O(N__10255),
            .I(N__10251));
    InMux I__1453 (
            .O(N__10254),
            .I(N__10248));
    Odrv4 I__1452 (
            .O(N__10251),
            .I(\c0.data_in_0_Z0Z_4 ));
    LocalMux I__1451 (
            .O(N__10248),
            .I(\c0.data_in_0_Z0Z_4 ));
    InMux I__1450 (
            .O(N__10243),
            .I(N__10238));
    InMux I__1449 (
            .O(N__10242),
            .I(N__10235));
    InMux I__1448 (
            .O(N__10241),
            .I(N__10232));
    LocalMux I__1447 (
            .O(N__10238),
            .I(\c0.data_in_1_Z0Z_0 ));
    LocalMux I__1446 (
            .O(N__10235),
            .I(\c0.data_in_1_Z0Z_0 ));
    LocalMux I__1445 (
            .O(N__10232),
            .I(\c0.data_in_1_Z0Z_0 ));
    InMux I__1444 (
            .O(N__10225),
            .I(N__10222));
    LocalMux I__1443 (
            .O(N__10222),
            .I(N__10219));
    Span12Mux_v I__1442 (
            .O(N__10219),
            .I(N__10215));
    InMux I__1441 (
            .O(N__10218),
            .I(N__10212));
    Odrv12 I__1440 (
            .O(N__10215),
            .I(\c0.rx_data_3 ));
    LocalMux I__1439 (
            .O(N__10212),
            .I(\c0.rx_data_3 ));
    InMux I__1438 (
            .O(N__10207),
            .I(N__10204));
    LocalMux I__1437 (
            .O(N__10204),
            .I(N__10200));
    CascadeMux I__1436 (
            .O(N__10203),
            .I(N__10197));
    Span12Mux_v I__1435 (
            .O(N__10200),
            .I(N__10194));
    InMux I__1434 (
            .O(N__10197),
            .I(N__10191));
    Odrv12 I__1433 (
            .O(N__10194),
            .I(\c0.rx_data_1 ));
    LocalMux I__1432 (
            .O(N__10191),
            .I(\c0.rx_data_1 ));
    InMux I__1431 (
            .O(N__10186),
            .I(N__10182));
    InMux I__1430 (
            .O(N__10185),
            .I(N__10179));
    LocalMux I__1429 (
            .O(N__10182),
            .I(\c0.dataZ0Z_0 ));
    LocalMux I__1428 (
            .O(N__10179),
            .I(\c0.dataZ0Z_0 ));
    InMux I__1427 (
            .O(N__10174),
            .I(N__10170));
    InMux I__1426 (
            .O(N__10173),
            .I(N__10167));
    LocalMux I__1425 (
            .O(N__10170),
            .I(\c0.dataZ0Z_14 ));
    LocalMux I__1424 (
            .O(N__10167),
            .I(\c0.dataZ0Z_14 ));
    InMux I__1423 (
            .O(N__10162),
            .I(N__10158));
    InMux I__1422 (
            .O(N__10161),
            .I(N__10155));
    LocalMux I__1421 (
            .O(N__10158),
            .I(\c0.dataZ0Z_11 ));
    LocalMux I__1420 (
            .O(N__10155),
            .I(\c0.dataZ0Z_11 ));
    InMux I__1419 (
            .O(N__10150),
            .I(N__10146));
    InMux I__1418 (
            .O(N__10149),
            .I(N__10143));
    LocalMux I__1417 (
            .O(N__10146),
            .I(\c0.dataZ0Z_2 ));
    LocalMux I__1416 (
            .O(N__10143),
            .I(\c0.dataZ0Z_2 ));
    InMux I__1415 (
            .O(N__10138),
            .I(N__10134));
    InMux I__1414 (
            .O(N__10137),
            .I(N__10131));
    LocalMux I__1413 (
            .O(N__10134),
            .I(\c0.dataZ0Z_15 ));
    LocalMux I__1412 (
            .O(N__10131),
            .I(\c0.dataZ0Z_15 ));
    InMux I__1411 (
            .O(N__10126),
            .I(N__10122));
    InMux I__1410 (
            .O(N__10125),
            .I(N__10119));
    LocalMux I__1409 (
            .O(N__10122),
            .I(\c0.dataZ0Z_4 ));
    LocalMux I__1408 (
            .O(N__10119),
            .I(\c0.dataZ0Z_4 ));
    InMux I__1407 (
            .O(N__10114),
            .I(N__10110));
    InMux I__1406 (
            .O(N__10113),
            .I(N__10107));
    LocalMux I__1405 (
            .O(N__10110),
            .I(\c0.dataZ0Z_8 ));
    LocalMux I__1404 (
            .O(N__10107),
            .I(\c0.dataZ0Z_8 ));
    InMux I__1403 (
            .O(N__10102),
            .I(N__10099));
    LocalMux I__1402 (
            .O(N__10099),
            .I(\c0.nextCRC16_3_0_a2_6_0_15 ));
    CascadeMux I__1401 (
            .O(N__10096),
            .I(\c0.nextCRC16_3_9_cascade_ ));
    CascadeMux I__1400 (
            .O(N__10093),
            .I(\c0.N_106_cascade_ ));
    InMux I__1399 (
            .O(N__10090),
            .I(N__10087));
    LocalMux I__1398 (
            .O(N__10087),
            .I(N__10084));
    Span12Mux_v I__1397 (
            .O(N__10084),
            .I(N__10080));
    InMux I__1396 (
            .O(N__10083),
            .I(N__10077));
    Odrv12 I__1395 (
            .O(N__10080),
            .I(\c0.N_92 ));
    LocalMux I__1394 (
            .O(N__10077),
            .I(\c0.N_92 ));
    InMux I__1393 (
            .O(N__10072),
            .I(N__10066));
    InMux I__1392 (
            .O(N__10071),
            .I(N__10066));
    LocalMux I__1391 (
            .O(N__10066),
            .I(\c0.N_106 ));
    CascadeMux I__1390 (
            .O(N__10063),
            .I(N__10060));
    InMux I__1389 (
            .O(N__10060),
            .I(N__10057));
    LocalMux I__1388 (
            .O(N__10057),
            .I(\c0.data_out_7_Z0Z_0 ));
    CascadeMux I__1387 (
            .O(N__10054),
            .I(N__10051));
    InMux I__1386 (
            .O(N__10051),
            .I(N__10048));
    LocalMux I__1385 (
            .O(N__10048),
            .I(N__10045));
    Odrv4 I__1384 (
            .O(N__10045),
            .I(\c0.nextCRC16_3_0_a2_0_10 ));
    InMux I__1383 (
            .O(N__10042),
            .I(N__10039));
    LocalMux I__1382 (
            .O(N__10039),
            .I(N__10035));
    InMux I__1381 (
            .O(N__10038),
            .I(N__10032));
    Odrv4 I__1380 (
            .O(N__10035),
            .I(\c0.dataZ0Z_12 ));
    LocalMux I__1379 (
            .O(N__10032),
            .I(\c0.dataZ0Z_12 ));
    InMux I__1378 (
            .O(N__10027),
            .I(N__10024));
    LocalMux I__1377 (
            .O(N__10024),
            .I(N__10019));
    InMux I__1376 (
            .O(N__10023),
            .I(N__10016));
    InMux I__1375 (
            .O(N__10022),
            .I(N__10013));
    Odrv4 I__1374 (
            .O(N__10019),
            .I(\c0.N_77 ));
    LocalMux I__1373 (
            .O(N__10016),
            .I(\c0.N_77 ));
    LocalMux I__1372 (
            .O(N__10013),
            .I(\c0.N_77 ));
    InMux I__1371 (
            .O(N__10006),
            .I(N__10002));
    InMux I__1370 (
            .O(N__10005),
            .I(N__9999));
    LocalMux I__1369 (
            .O(N__10002),
            .I(N__9993));
    LocalMux I__1368 (
            .O(N__9999),
            .I(N__9993));
    InMux I__1367 (
            .O(N__9998),
            .I(N__9990));
    Odrv4 I__1366 (
            .O(N__9993),
            .I(\c0.N_76 ));
    LocalMux I__1365 (
            .O(N__9990),
            .I(\c0.N_76 ));
    InMux I__1364 (
            .O(N__9985),
            .I(N__9981));
    CascadeMux I__1363 (
            .O(N__9984),
            .I(N__9976));
    LocalMux I__1362 (
            .O(N__9981),
            .I(N__9973));
    InMux I__1361 (
            .O(N__9980),
            .I(N__9970));
    InMux I__1360 (
            .O(N__9979),
            .I(N__9965));
    InMux I__1359 (
            .O(N__9976),
            .I(N__9965));
    Odrv4 I__1358 (
            .O(N__9973),
            .I(\c0.tx.r_SM_Main_dup_4 ));
    LocalMux I__1357 (
            .O(N__9970),
            .I(\c0.tx.r_SM_Main_dup_4 ));
    LocalMux I__1356 (
            .O(N__9965),
            .I(\c0.tx.r_SM_Main_dup_4 ));
    InMux I__1355 (
            .O(N__9958),
            .I(N__9954));
    CascadeMux I__1354 (
            .O(N__9957),
            .I(N__9951));
    LocalMux I__1353 (
            .O(N__9954),
            .I(N__9948));
    InMux I__1352 (
            .O(N__9951),
            .I(N__9944));
    Span4Mux_h I__1351 (
            .O(N__9948),
            .I(N__9941));
    CascadeMux I__1350 (
            .O(N__9947),
            .I(N__9937));
    LocalMux I__1349 (
            .O(N__9944),
            .I(N__9933));
    Span4Mux_h I__1348 (
            .O(N__9941),
            .I(N__9930));
    InMux I__1347 (
            .O(N__9940),
            .I(N__9927));
    InMux I__1346 (
            .O(N__9937),
            .I(N__9922));
    InMux I__1345 (
            .O(N__9936),
            .I(N__9922));
    Odrv4 I__1344 (
            .O(N__9933),
            .I(\c0.tx_transmitZ0 ));
    Odrv4 I__1343 (
            .O(N__9930),
            .I(\c0.tx_transmitZ0 ));
    LocalMux I__1342 (
            .O(N__9927),
            .I(\c0.tx_transmitZ0 ));
    LocalMux I__1341 (
            .O(N__9922),
            .I(\c0.tx_transmitZ0 ));
    CascadeMux I__1340 (
            .O(N__9913),
            .I(N__9910));
    InMux I__1339 (
            .O(N__9910),
            .I(N__9907));
    LocalMux I__1338 (
            .O(N__9907),
            .I(\c0.tx.r_SM_Main_RNO_0Z0Z_0 ));
    InMux I__1337 (
            .O(N__9904),
            .I(N__9898));
    InMux I__1336 (
            .O(N__9903),
            .I(N__9891));
    InMux I__1335 (
            .O(N__9902),
            .I(N__9891));
    InMux I__1334 (
            .O(N__9901),
            .I(N__9891));
    LocalMux I__1333 (
            .O(N__9898),
            .I(\c0.tx.N_171_0 ));
    LocalMux I__1332 (
            .O(N__9891),
            .I(\c0.tx.N_171_0 ));
    CascadeMux I__1331 (
            .O(N__9886),
            .I(\c0.tx.r_SM_Main_RNO_0Z0Z_2_cascade_ ));
    CascadeMux I__1330 (
            .O(N__9883),
            .I(N__9880));
    InMux I__1329 (
            .O(N__9880),
            .I(N__9873));
    InMux I__1328 (
            .O(N__9879),
            .I(N__9864));
    InMux I__1327 (
            .O(N__9878),
            .I(N__9864));
    InMux I__1326 (
            .O(N__9877),
            .I(N__9864));
    InMux I__1325 (
            .O(N__9876),
            .I(N__9864));
    LocalMux I__1324 (
            .O(N__9873),
            .I(N__9858));
    LocalMux I__1323 (
            .O(N__9864),
            .I(N__9858));
    InMux I__1322 (
            .O(N__9863),
            .I(N__9849));
    Span4Mux_h I__1321 (
            .O(N__9858),
            .I(N__9846));
    InMux I__1320 (
            .O(N__9857),
            .I(N__9841));
    InMux I__1319 (
            .O(N__9856),
            .I(N__9841));
    InMux I__1318 (
            .O(N__9855),
            .I(N__9832));
    InMux I__1317 (
            .O(N__9854),
            .I(N__9832));
    InMux I__1316 (
            .O(N__9853),
            .I(N__9832));
    InMux I__1315 (
            .O(N__9852),
            .I(N__9832));
    LocalMux I__1314 (
            .O(N__9849),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    Odrv4 I__1313 (
            .O(N__9846),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    LocalMux I__1312 (
            .O(N__9841),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    LocalMux I__1311 (
            .O(N__9832),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    CascadeMux I__1310 (
            .O(N__9823),
            .I(N__9811));
    InMux I__1309 (
            .O(N__9822),
            .I(N__9808));
    InMux I__1308 (
            .O(N__9821),
            .I(N__9803));
    InMux I__1307 (
            .O(N__9820),
            .I(N__9803));
    InMux I__1306 (
            .O(N__9819),
            .I(N__9796));
    InMux I__1305 (
            .O(N__9818),
            .I(N__9796));
    InMux I__1304 (
            .O(N__9817),
            .I(N__9796));
    InMux I__1303 (
            .O(N__9816),
            .I(N__9787));
    InMux I__1302 (
            .O(N__9815),
            .I(N__9787));
    InMux I__1301 (
            .O(N__9814),
            .I(N__9787));
    InMux I__1300 (
            .O(N__9811),
            .I(N__9787));
    LocalMux I__1299 (
            .O(N__9808),
            .I(\c0.tx.N_90_dup ));
    LocalMux I__1298 (
            .O(N__9803),
            .I(\c0.tx.N_90_dup ));
    LocalMux I__1297 (
            .O(N__9796),
            .I(\c0.tx.N_90_dup ));
    LocalMux I__1296 (
            .O(N__9787),
            .I(\c0.tx.N_90_dup ));
    InMux I__1295 (
            .O(N__9778),
            .I(N__9775));
    LocalMux I__1294 (
            .O(N__9775),
            .I(N__9772));
    Span4Mux_v I__1293 (
            .O(N__9772),
            .I(N__9763));
    InMux I__1292 (
            .O(N__9771),
            .I(N__9760));
    InMux I__1291 (
            .O(N__9770),
            .I(N__9757));
    InMux I__1290 (
            .O(N__9769),
            .I(N__9748));
    InMux I__1289 (
            .O(N__9768),
            .I(N__9748));
    InMux I__1288 (
            .O(N__9767),
            .I(N__9748));
    InMux I__1287 (
            .O(N__9766),
            .I(N__9748));
    Sp12to4 I__1286 (
            .O(N__9763),
            .I(N__9741));
    LocalMux I__1285 (
            .O(N__9760),
            .I(N__9741));
    LocalMux I__1284 (
            .O(N__9757),
            .I(N__9741));
    LocalMux I__1283 (
            .O(N__9748),
            .I(\c0.tx.r_Clock_Count12_THRU_CO ));
    Odrv12 I__1282 (
            .O(N__9741),
            .I(\c0.tx.r_Clock_Count12_THRU_CO ));
    InMux I__1281 (
            .O(N__9736),
            .I(N__9729));
    InMux I__1280 (
            .O(N__9735),
            .I(N__9729));
    InMux I__1279 (
            .O(N__9734),
            .I(N__9726));
    LocalMux I__1278 (
            .O(N__9729),
            .I(\c0.tx.r_SM_Main_RNIVDI71Z0Z_2 ));
    LocalMux I__1277 (
            .O(N__9726),
            .I(\c0.tx.r_SM_Main_RNIVDI71Z0Z_2 ));
    InMux I__1276 (
            .O(N__9721),
            .I(N__9718));
    LocalMux I__1275 (
            .O(N__9718),
            .I(\c0.i12_4_and ));
    CascadeMux I__1274 (
            .O(N__9715),
            .I(\c0.tx.r_Bit_Index_RNO_0Z0Z_2_cascade_ ));
    CascadeMux I__1273 (
            .O(N__9712),
            .I(\c0.tx.r_Tx_Active_1_sqmuxa_cascade_ ));
    InMux I__1272 (
            .O(N__9709),
            .I(N__9706));
    LocalMux I__1271 (
            .O(N__9706),
            .I(\c0.tx.N_90_ip_RNIVJLQZ0 ));
    InMux I__1270 (
            .O(N__9703),
            .I(N__9694));
    InMux I__1269 (
            .O(N__9702),
            .I(N__9694));
    InMux I__1268 (
            .O(N__9701),
            .I(N__9694));
    LocalMux I__1267 (
            .O(N__9694),
            .I(\c0.tx_active ));
    CascadeMux I__1266 (
            .O(N__9691),
            .I(\c0.tx.N_90_ip_RNI1U1EZ0_cascade_ ));
    InMux I__1265 (
            .O(N__9688),
            .I(N__9685));
    LocalMux I__1264 (
            .O(N__9685),
            .I(\c0.i12_5_and ));
    InMux I__1263 (
            .O(N__9682),
            .I(N__9679));
    LocalMux I__1262 (
            .O(N__9679),
            .I(\c0.i12_6_and ));
    InMux I__1261 (
            .O(N__9676),
            .I(N__9673));
    LocalMux I__1260 (
            .O(N__9673),
            .I(\c0.i12_2_and ));
    InMux I__1259 (
            .O(N__9670),
            .I(\c0.data_cry_10 ));
    InMux I__1258 (
            .O(N__9667),
            .I(\c0.data_cry_11 ));
    InMux I__1257 (
            .O(N__9664),
            .I(N__9661));
    LocalMux I__1256 (
            .O(N__9661),
            .I(N__9657));
    InMux I__1255 (
            .O(N__9660),
            .I(N__9654));
    Odrv4 I__1254 (
            .O(N__9657),
            .I(\c0.dataZ0Z_13 ));
    LocalMux I__1253 (
            .O(N__9654),
            .I(\c0.dataZ0Z_13 ));
    InMux I__1252 (
            .O(N__9649),
            .I(\c0.data_cry_12 ));
    InMux I__1251 (
            .O(N__9646),
            .I(\c0.data_cry_13 ));
    InMux I__1250 (
            .O(N__9643),
            .I(\c0.data_cry_14 ));
    InMux I__1249 (
            .O(N__9640),
            .I(N__9637));
    LocalMux I__1248 (
            .O(N__9637),
            .I(\c0.i12_3_and ));
    InMux I__1247 (
            .O(N__9634),
            .I(\c0.data_cry_1 ));
    InMux I__1246 (
            .O(N__9631),
            .I(N__9628));
    LocalMux I__1245 (
            .O(N__9628),
            .I(N__9624));
    InMux I__1244 (
            .O(N__9627),
            .I(N__9621));
    Odrv4 I__1243 (
            .O(N__9624),
            .I(\c0.dataZ0Z_3 ));
    LocalMux I__1242 (
            .O(N__9621),
            .I(\c0.dataZ0Z_3 ));
    InMux I__1241 (
            .O(N__9616),
            .I(\c0.data_cry_2 ));
    InMux I__1240 (
            .O(N__9613),
            .I(\c0.data_cry_3 ));
    InMux I__1239 (
            .O(N__9610),
            .I(N__9607));
    LocalMux I__1238 (
            .O(N__9607),
            .I(N__9603));
    InMux I__1237 (
            .O(N__9606),
            .I(N__9600));
    Odrv4 I__1236 (
            .O(N__9603),
            .I(\c0.dataZ0Z_5 ));
    LocalMux I__1235 (
            .O(N__9600),
            .I(\c0.dataZ0Z_5 ));
    InMux I__1234 (
            .O(N__9595),
            .I(\c0.data_cry_4 ));
    InMux I__1233 (
            .O(N__9592),
            .I(\c0.data_cry_5 ));
    InMux I__1232 (
            .O(N__9589),
            .I(N__9585));
    InMux I__1231 (
            .O(N__9588),
            .I(N__9582));
    LocalMux I__1230 (
            .O(N__9585),
            .I(\c0.dataZ0Z_7 ));
    LocalMux I__1229 (
            .O(N__9582),
            .I(\c0.dataZ0Z_7 ));
    InMux I__1228 (
            .O(N__9577),
            .I(\c0.data_cry_6 ));
    InMux I__1227 (
            .O(N__9574),
            .I(bfn_9_28_0_));
    InMux I__1226 (
            .O(N__9571),
            .I(N__9568));
    LocalMux I__1225 (
            .O(N__9568),
            .I(N__9564));
    InMux I__1224 (
            .O(N__9567),
            .I(N__9561));
    Odrv4 I__1223 (
            .O(N__9564),
            .I(\c0.dataZ0Z_9 ));
    LocalMux I__1222 (
            .O(N__9561),
            .I(\c0.dataZ0Z_9 ));
    InMux I__1221 (
            .O(N__9556),
            .I(\c0.data_cry_8 ));
    InMux I__1220 (
            .O(N__9553),
            .I(N__9550));
    LocalMux I__1219 (
            .O(N__9550),
            .I(N__9546));
    InMux I__1218 (
            .O(N__9549),
            .I(N__9543));
    Odrv4 I__1217 (
            .O(N__9546),
            .I(\c0.dataZ0Z_10 ));
    LocalMux I__1216 (
            .O(N__9543),
            .I(\c0.dataZ0Z_10 ));
    InMux I__1215 (
            .O(N__9538),
            .I(\c0.data_cry_9 ));
    InMux I__1214 (
            .O(N__9535),
            .I(bfn_9_27_0_));
    InMux I__1213 (
            .O(N__9532),
            .I(N__9528));
    InMux I__1212 (
            .O(N__9531),
            .I(N__9525));
    LocalMux I__1211 (
            .O(N__9528),
            .I(\c0.dataZ0Z_1 ));
    LocalMux I__1210 (
            .O(N__9525),
            .I(\c0.dataZ0Z_1 ));
    InMux I__1209 (
            .O(N__9520),
            .I(\c0.data_cry_0 ));
    InMux I__1208 (
            .O(N__9517),
            .I(N__9514));
    LocalMux I__1207 (
            .O(N__9514),
            .I(N__9511));
    Odrv12 I__1206 (
            .O(N__9511),
            .I(\c0.tx.r_Clock_Count_RNO_0Z0Z_2 ));
    InMux I__1205 (
            .O(N__9508),
            .I(\c0.tx.un1_r_Clock_Count_cry_1 ));
    InMux I__1204 (
            .O(N__9505),
            .I(\c0.tx.un1_r_Clock_Count_cry_2 ));
    InMux I__1203 (
            .O(N__9502),
            .I(N__9499));
    LocalMux I__1202 (
            .O(N__9499),
            .I(N__9496));
    Odrv12 I__1201 (
            .O(N__9496),
            .I(\c0.tx.r_Clock_Count_RNO_0Z0Z_3 ));
    InMux I__1200 (
            .O(N__9493),
            .I(N__9489));
    InMux I__1199 (
            .O(N__9492),
            .I(N__9486));
    LocalMux I__1198 (
            .O(N__9489),
            .I(N__9480));
    LocalMux I__1197 (
            .O(N__9486),
            .I(N__9480));
    InMux I__1196 (
            .O(N__9485),
            .I(N__9477));
    Odrv12 I__1195 (
            .O(N__9480),
            .I(\c0.tx.r_Clock_CountZ0Z_2 ));
    LocalMux I__1194 (
            .O(N__9477),
            .I(\c0.tx.r_Clock_CountZ0Z_2 ));
    InMux I__1193 (
            .O(N__9472),
            .I(N__9468));
    InMux I__1192 (
            .O(N__9471),
            .I(N__9465));
    LocalMux I__1191 (
            .O(N__9468),
            .I(N__9459));
    LocalMux I__1190 (
            .O(N__9465),
            .I(N__9459));
    InMux I__1189 (
            .O(N__9464),
            .I(N__9456));
    Odrv12 I__1188 (
            .O(N__9459),
            .I(\c0.tx.r_Clock_CountZ0Z_1 ));
    LocalMux I__1187 (
            .O(N__9456),
            .I(\c0.tx.r_Clock_CountZ0Z_1 ));
    CascadeMux I__1186 (
            .O(N__9451),
            .I(N__9447));
    InMux I__1185 (
            .O(N__9450),
            .I(N__9442));
    InMux I__1184 (
            .O(N__9447),
            .I(N__9442));
    LocalMux I__1183 (
            .O(N__9442),
            .I(N__9439));
    Span4Mux_h I__1182 (
            .O(N__9439),
            .I(N__9435));
    InMux I__1181 (
            .O(N__9438),
            .I(N__9432));
    Odrv4 I__1180 (
            .O(N__9435),
            .I(\c0.tx.r_Clock_CountZ0Z_3 ));
    LocalMux I__1179 (
            .O(N__9432),
            .I(\c0.tx.r_Clock_CountZ0Z_3 ));
    InMux I__1178 (
            .O(N__9427),
            .I(N__9421));
    InMux I__1177 (
            .O(N__9426),
            .I(N__9421));
    LocalMux I__1176 (
            .O(N__9421),
            .I(N__9417));
    InMux I__1175 (
            .O(N__9420),
            .I(N__9414));
    Odrv12 I__1174 (
            .O(N__9417),
            .I(\c0.tx.r_Clock_CountZ0Z_0 ));
    LocalMux I__1173 (
            .O(N__9414),
            .I(\c0.tx.r_Clock_CountZ0Z_0 ));
    InMux I__1172 (
            .O(N__9409),
            .I(N__9406));
    LocalMux I__1171 (
            .O(N__9406),
            .I(N__9403));
    Span4Mux_h I__1170 (
            .O(N__9403),
            .I(N__9400));
    Odrv4 I__1169 (
            .O(N__9400),
            .I(\c0.tx.r_SM_Main_RNO_0Z0Z_1 ));
    CascadeMux I__1168 (
            .O(N__9397),
            .I(\c0.tx.N_171_0_cascade_ ));
    CascadeMux I__1167 (
            .O(N__9394),
            .I(\c0.nextCRC16_3_0_a2_1_8_cascade_ ));
    InMux I__1166 (
            .O(N__9391),
            .I(N__9388));
    LocalMux I__1165 (
            .O(N__9388),
            .I(\c0.data_out_6_Z0Z_0 ));
    CascadeMux I__1164 (
            .O(N__9385),
            .I(N__9382));
    InMux I__1163 (
            .O(N__9382),
            .I(N__9379));
    LocalMux I__1162 (
            .O(N__9379),
            .I(N__9376));
    Span12Mux_v I__1161 (
            .O(N__9376),
            .I(N__9373));
    Odrv12 I__1160 (
            .O(N__9373),
            .I(\c0.N_71 ));
    CascadeMux I__1159 (
            .O(N__9370),
            .I(\c0.tx.N_90_ip_RNIVJLQZ0_cascade_ ));
    InMux I__1158 (
            .O(N__9367),
            .I(N__9364));
    LocalMux I__1157 (
            .O(N__9364),
            .I(\c0.tx.r_SM_Main_illegal_0 ));
    CascadeMux I__1156 (
            .O(N__9361),
            .I(\c0.tx.N_90_dup_cascade_ ));
    InMux I__1155 (
            .O(N__9358),
            .I(N__9355));
    LocalMux I__1154 (
            .O(N__9355),
            .I(\c0.tx.N_83_0 ));
    InMux I__1153 (
            .O(N__9352),
            .I(N__9348));
    CascadeMux I__1152 (
            .O(N__9351),
            .I(N__9345));
    LocalMux I__1151 (
            .O(N__9348),
            .I(N__9342));
    InMux I__1150 (
            .O(N__9345),
            .I(N__9339));
    Odrv4 I__1149 (
            .O(N__9342),
            .I(\c0.tx.r_Clock_Count_0_sqmuxa ));
    LocalMux I__1148 (
            .O(N__9339),
            .I(\c0.tx.r_Clock_Count_0_sqmuxa ));
    InMux I__1147 (
            .O(N__9334),
            .I(N__9331));
    LocalMux I__1146 (
            .O(N__9331),
            .I(N__9328));
    Span4Mux_h I__1145 (
            .O(N__9328),
            .I(N__9325));
    Odrv4 I__1144 (
            .O(N__9325),
            .I(\c0.tx.r_Clock_Count_RNO_0Z0Z_0 ));
    InMux I__1143 (
            .O(N__9322),
            .I(N__9319));
    LocalMux I__1142 (
            .O(N__9319),
            .I(N__9316));
    Span4Mux_h I__1141 (
            .O(N__9316),
            .I(N__9313));
    Odrv4 I__1140 (
            .O(N__9313),
            .I(\c0.tx.r_Clock_Count_RNO_0Z0Z_1 ));
    InMux I__1139 (
            .O(N__9310),
            .I(\c0.tx.un1_r_Clock_Count_cry_0 ));
    InMux I__1138 (
            .O(N__9307),
            .I(N__9304));
    LocalMux I__1137 (
            .O(N__9304),
            .I(\c0.i12_1_and ));
    InMux I__1136 (
            .O(N__9301),
            .I(N__9298));
    LocalMux I__1135 (
            .O(N__9298),
            .I(N__9295));
    Span4Mux_v I__1134 (
            .O(N__9295),
            .I(N__9291));
    InMux I__1133 (
            .O(N__9294),
            .I(N__9288));
    Odrv4 I__1132 (
            .O(N__9291),
            .I(blink_counterZ0Z_21));
    LocalMux I__1131 (
            .O(N__9288),
            .I(blink_counterZ0Z_21));
    InMux I__1130 (
            .O(N__9283),
            .I(N__9277));
    InMux I__1129 (
            .O(N__9282),
            .I(N__9277));
    LocalMux I__1128 (
            .O(N__9277),
            .I(N__9274));
    Span4Mux_v I__1127 (
            .O(N__9274),
            .I(N__9270));
    InMux I__1126 (
            .O(N__9273),
            .I(N__9267));
    Odrv4 I__1125 (
            .O(N__9270),
            .I(blink_counterZ0Z_22));
    LocalMux I__1124 (
            .O(N__9267),
            .I(blink_counterZ0Z_22));
    CascadeMux I__1123 (
            .O(N__9262),
            .I(N__9259));
    InMux I__1122 (
            .O(N__9259),
            .I(N__9253));
    InMux I__1121 (
            .O(N__9258),
            .I(N__9253));
    LocalMux I__1120 (
            .O(N__9253),
            .I(N__9250));
    Span4Mux_v I__1119 (
            .O(N__9250),
            .I(N__9246));
    InMux I__1118 (
            .O(N__9249),
            .I(N__9243));
    Odrv4 I__1117 (
            .O(N__9246),
            .I(blink_counterZ0Z_24));
    LocalMux I__1116 (
            .O(N__9243),
            .I(blink_counterZ0Z_24));
    InMux I__1115 (
            .O(N__9238),
            .I(N__9235));
    LocalMux I__1114 (
            .O(N__9235),
            .I(N_12));
    InMux I__1113 (
            .O(N__9232),
            .I(N__9226));
    InMux I__1112 (
            .O(N__9231),
            .I(N__9226));
    LocalMux I__1111 (
            .O(N__9226),
            .I(N__9223));
    Span4Mux_v I__1110 (
            .O(N__9223),
            .I(N__9219));
    InMux I__1109 (
            .O(N__9222),
            .I(N__9216));
    Odrv4 I__1108 (
            .O(N__9219),
            .I(blink_counterZ0Z_25));
    LocalMux I__1107 (
            .O(N__9216),
            .I(blink_counterZ0Z_25));
    CascadeMux I__1106 (
            .O(N__9211),
            .I(N_8_0_cascade_));
    InMux I__1105 (
            .O(N__9208),
            .I(N__9205));
    LocalMux I__1104 (
            .O(N__9205),
            .I(N__9202));
    Span4Mux_h I__1103 (
            .O(N__9202),
            .I(N__9198));
    InMux I__1102 (
            .O(N__9201),
            .I(N__9195));
    Odrv4 I__1101 (
            .O(N__9198),
            .I(blink_counterZ0Z_23));
    LocalMux I__1100 (
            .O(N__9195),
            .I(blink_counterZ0Z_23));
    IoInMux I__1099 (
            .O(N__9190),
            .I(N__9187));
    LocalMux I__1098 (
            .O(N__9187),
            .I(N__9184));
    Span4Mux_s1_h I__1097 (
            .O(N__9184),
            .I(N__9181));
    Sp12to4 I__1096 (
            .O(N__9181),
            .I(N__9178));
    Span12Mux_s11_v I__1095 (
            .O(N__9178),
            .I(N__9175));
    Odrv12 I__1094 (
            .O(N__9175),
            .I(LED_c));
    CascadeMux I__1093 (
            .O(N__9172),
            .I(N__9169));
    InMux I__1092 (
            .O(N__9169),
            .I(N__9166));
    LocalMux I__1091 (
            .O(N__9166),
            .I(\c0.i12_7_and ));
    InMux I__1090 (
            .O(N__9163),
            .I(bfn_9_20_0_));
    InMux I__1089 (
            .O(N__9160),
            .I(N__9157));
    LocalMux I__1088 (
            .O(N__9157),
            .I(\c0.i12_0_and ));
    CascadeMux I__1087 (
            .O(N__9154),
            .I(N__9151));
    InMux I__1086 (
            .O(N__9151),
            .I(N__9148));
    LocalMux I__1085 (
            .O(N__9148),
            .I(\c0.rx.r_SM_Main_ns_0_i_a2_1_0_2 ));
    InMux I__1084 (
            .O(N__9145),
            .I(N__9137));
    InMux I__1083 (
            .O(N__9144),
            .I(N__9132));
    InMux I__1082 (
            .O(N__9143),
            .I(N__9132));
    InMux I__1081 (
            .O(N__9142),
            .I(N__9125));
    InMux I__1080 (
            .O(N__9141),
            .I(N__9125));
    InMux I__1079 (
            .O(N__9140),
            .I(N__9125));
    LocalMux I__1078 (
            .O(N__9137),
            .I(\c0.rx.r_SM_Main_dup_1 ));
    LocalMux I__1077 (
            .O(N__9132),
            .I(\c0.rx.r_SM_Main_dup_1 ));
    LocalMux I__1076 (
            .O(N__9125),
            .I(\c0.rx.r_SM_Main_dup_1 ));
    CascadeMux I__1075 (
            .O(N__9118),
            .I(\c0.rx.un1_r_Rx_DV7_i_0_cascade_ ));
    InMux I__1074 (
            .O(N__9115),
            .I(N__9112));
    LocalMux I__1073 (
            .O(N__9112),
            .I(N__9109));
    Span4Mux_h I__1072 (
            .O(N__9109),
            .I(N__9106));
    Odrv4 I__1071 (
            .O(N__9106),
            .I(\c0.rx.r_Rx_DV_RNOZ0Z_0 ));
    InMux I__1070 (
            .O(N__9103),
            .I(N__9097));
    InMux I__1069 (
            .O(N__9102),
            .I(N__9097));
    LocalMux I__1068 (
            .O(N__9097),
            .I(N__9088));
    InMux I__1067 (
            .O(N__9096),
            .I(N__9081));
    InMux I__1066 (
            .O(N__9095),
            .I(N__9081));
    InMux I__1065 (
            .O(N__9094),
            .I(N__9081));
    InMux I__1064 (
            .O(N__9093),
            .I(N__9074));
    InMux I__1063 (
            .O(N__9092),
            .I(N__9074));
    InMux I__1062 (
            .O(N__9091),
            .I(N__9074));
    Odrv12 I__1061 (
            .O(N__9088),
            .I(\c0.rx.r_SM_Main_dup_2 ));
    LocalMux I__1060 (
            .O(N__9081),
            .I(\c0.rx.r_SM_Main_dup_2 ));
    LocalMux I__1059 (
            .O(N__9074),
            .I(\c0.rx.r_SM_Main_dup_2 ));
    InMux I__1058 (
            .O(N__9067),
            .I(N__9064));
    LocalMux I__1057 (
            .O(N__9064),
            .I(\c0.rx.r_SM_Main_ns_0_i_0_0_2 ));
    InMux I__1056 (
            .O(N__9061),
            .I(N__9057));
    InMux I__1055 (
            .O(N__9060),
            .I(N__9054));
    LocalMux I__1054 (
            .O(N__9057),
            .I(N__9039));
    LocalMux I__1053 (
            .O(N__9054),
            .I(N__9039));
    InMux I__1052 (
            .O(N__9053),
            .I(N__9036));
    InMux I__1051 (
            .O(N__9052),
            .I(N__9033));
    InMux I__1050 (
            .O(N__9051),
            .I(N__9028));
    InMux I__1049 (
            .O(N__9050),
            .I(N__9028));
    InMux I__1048 (
            .O(N__9049),
            .I(N__9025));
    InMux I__1047 (
            .O(N__9048),
            .I(N__9022));
    InMux I__1046 (
            .O(N__9047),
            .I(N__9019));
    InMux I__1045 (
            .O(N__9046),
            .I(N__9016));
    InMux I__1044 (
            .O(N__9045),
            .I(N__9013));
    InMux I__1043 (
            .O(N__9044),
            .I(N__9010));
    Span4Mux_v I__1042 (
            .O(N__9039),
            .I(N__9005));
    LocalMux I__1041 (
            .O(N__9036),
            .I(N__9005));
    LocalMux I__1040 (
            .O(N__9033),
            .I(N__8990));
    LocalMux I__1039 (
            .O(N__9028),
            .I(N__8990));
    LocalMux I__1038 (
            .O(N__9025),
            .I(N__8990));
    LocalMux I__1037 (
            .O(N__9022),
            .I(N__8990));
    LocalMux I__1036 (
            .O(N__9019),
            .I(N__8990));
    LocalMux I__1035 (
            .O(N__9016),
            .I(N__8990));
    LocalMux I__1034 (
            .O(N__9013),
            .I(N__8990));
    LocalMux I__1033 (
            .O(N__9010),
            .I(N__8987));
    Span4Mux_h I__1032 (
            .O(N__9005),
            .I(N__8984));
    Span4Mux_v I__1031 (
            .O(N__8990),
            .I(N__8981));
    Span4Mux_h I__1030 (
            .O(N__8987),
            .I(N__8976));
    Span4Mux_v I__1029 (
            .O(N__8984),
            .I(N__8976));
    Odrv4 I__1028 (
            .O(N__8981),
            .I(\c0.rx.r_Rx_DataZ0 ));
    Odrv4 I__1027 (
            .O(N__8976),
            .I(\c0.rx.r_Rx_DataZ0 ));
    InMux I__1026 (
            .O(N__8971),
            .I(N__8966));
    InMux I__1025 (
            .O(N__8970),
            .I(N__8963));
    InMux I__1024 (
            .O(N__8969),
            .I(N__8960));
    LocalMux I__1023 (
            .O(N__8966),
            .I(N__8957));
    LocalMux I__1022 (
            .O(N__8963),
            .I(\c0.rx.N_383 ));
    LocalMux I__1021 (
            .O(N__8960),
            .I(\c0.rx.N_383 ));
    Odrv4 I__1020 (
            .O(N__8957),
            .I(\c0.rx.N_383 ));
    InMux I__1019 (
            .O(N__8950),
            .I(N__8947));
    LocalMux I__1018 (
            .O(N__8947),
            .I(N__8940));
    InMux I__1017 (
            .O(N__8946),
            .I(N__8937));
    InMux I__1016 (
            .O(N__8945),
            .I(N__8930));
    InMux I__1015 (
            .O(N__8944),
            .I(N__8930));
    InMux I__1014 (
            .O(N__8943),
            .I(N__8930));
    Odrv4 I__1013 (
            .O(N__8940),
            .I(\c0.rx.N_321 ));
    LocalMux I__1012 (
            .O(N__8937),
            .I(\c0.rx.N_321 ));
    LocalMux I__1011 (
            .O(N__8930),
            .I(\c0.rx.N_321 ));
    CascadeMux I__1010 (
            .O(N__8923),
            .I(\c0.rx.r_Clock_Count_8_f0_0_a2_0_0_2_cascade_ ));
    CascadeMux I__1009 (
            .O(N__8920),
            .I(N__8916));
    CascadeMux I__1008 (
            .O(N__8919),
            .I(N__8913));
    InMux I__1007 (
            .O(N__8916),
            .I(N__8909));
    InMux I__1006 (
            .O(N__8913),
            .I(N__8906));
    InMux I__1005 (
            .O(N__8912),
            .I(N__8903));
    LocalMux I__1004 (
            .O(N__8909),
            .I(N__8898));
    LocalMux I__1003 (
            .O(N__8906),
            .I(N__8898));
    LocalMux I__1002 (
            .O(N__8903),
            .I(N__8893));
    Span4Mux_h I__1001 (
            .O(N__8898),
            .I(N__8893));
    Odrv4 I__1000 (
            .O(N__8893),
            .I(\c0.rx.N_371 ));
    InMux I__999 (
            .O(N__8890),
            .I(N__8887));
    LocalMux I__998 (
            .O(N__8887),
            .I(N__8878));
    InMux I__997 (
            .O(N__8886),
            .I(N__8869));
    InMux I__996 (
            .O(N__8885),
            .I(N__8869));
    InMux I__995 (
            .O(N__8884),
            .I(N__8869));
    InMux I__994 (
            .O(N__8883),
            .I(N__8869));
    InMux I__993 (
            .O(N__8882),
            .I(N__8866));
    InMux I__992 (
            .O(N__8881),
            .I(N__8863));
    Odrv4 I__991 (
            .O(N__8878),
            .I(\c0.rx.N_332 ));
    LocalMux I__990 (
            .O(N__8869),
            .I(\c0.rx.N_332 ));
    LocalMux I__989 (
            .O(N__8866),
            .I(\c0.rx.N_332 ));
    LocalMux I__988 (
            .O(N__8863),
            .I(\c0.rx.N_332 ));
    InMux I__987 (
            .O(N__8854),
            .I(N__8851));
    LocalMux I__986 (
            .O(N__8851),
            .I(N__8844));
    InMux I__985 (
            .O(N__8850),
            .I(N__8841));
    InMux I__984 (
            .O(N__8849),
            .I(N__8838));
    InMux I__983 (
            .O(N__8848),
            .I(N__8835));
    InMux I__982 (
            .O(N__8847),
            .I(N__8826));
    Span4Mux_v I__981 (
            .O(N__8844),
            .I(N__8821));
    LocalMux I__980 (
            .O(N__8841),
            .I(N__8821));
    LocalMux I__979 (
            .O(N__8838),
            .I(N__8818));
    LocalMux I__978 (
            .O(N__8835),
            .I(N__8815));
    InMux I__977 (
            .O(N__8834),
            .I(N__8810));
    InMux I__976 (
            .O(N__8833),
            .I(N__8810));
    InMux I__975 (
            .O(N__8832),
            .I(N__8801));
    InMux I__974 (
            .O(N__8831),
            .I(N__8801));
    InMux I__973 (
            .O(N__8830),
            .I(N__8801));
    InMux I__972 (
            .O(N__8829),
            .I(N__8801));
    LocalMux I__971 (
            .O(N__8826),
            .I(\c0.rx.r_SM_Main_RNI58REZ0Z_0 ));
    Odrv4 I__970 (
            .O(N__8821),
            .I(\c0.rx.r_SM_Main_RNI58REZ0Z_0 ));
    Odrv4 I__969 (
            .O(N__8818),
            .I(\c0.rx.r_SM_Main_RNI58REZ0Z_0 ));
    Odrv4 I__968 (
            .O(N__8815),
            .I(\c0.rx.r_SM_Main_RNI58REZ0Z_0 ));
    LocalMux I__967 (
            .O(N__8810),
            .I(\c0.rx.r_SM_Main_RNI58REZ0Z_0 ));
    LocalMux I__966 (
            .O(N__8801),
            .I(\c0.rx.r_SM_Main_RNI58REZ0Z_0 ));
    CascadeMux I__965 (
            .O(N__8788),
            .I(N__8783));
    CascadeMux I__964 (
            .O(N__8787),
            .I(N__8780));
    CascadeMux I__963 (
            .O(N__8786),
            .I(N__8776));
    InMux I__962 (
            .O(N__8783),
            .I(N__8770));
    InMux I__961 (
            .O(N__8780),
            .I(N__8770));
    InMux I__960 (
            .O(N__8779),
            .I(N__8767));
    InMux I__959 (
            .O(N__8776),
            .I(N__8764));
    CascadeMux I__958 (
            .O(N__8775),
            .I(N__8761));
    LocalMux I__957 (
            .O(N__8770),
            .I(N__8754));
    LocalMux I__956 (
            .O(N__8767),
            .I(N__8754));
    LocalMux I__955 (
            .O(N__8764),
            .I(N__8754));
    InMux I__954 (
            .O(N__8761),
            .I(N__8751));
    Odrv4 I__953 (
            .O(N__8754),
            .I(\c0.rx.N_361 ));
    LocalMux I__952 (
            .O(N__8751),
            .I(\c0.rx.N_361 ));
    InMux I__951 (
            .O(N__8746),
            .I(N__8743));
    LocalMux I__950 (
            .O(N__8743),
            .I(N__8740));
    Odrv12 I__949 (
            .O(N__8740),
            .I(\c0.rx.r_Clock_Count_RNO_0_0_3 ));
    InMux I__948 (
            .O(N__8737),
            .I(N__8731));
    InMux I__947 (
            .O(N__8736),
            .I(N__8728));
    InMux I__946 (
            .O(N__8735),
            .I(N__8723));
    InMux I__945 (
            .O(N__8734),
            .I(N__8723));
    LocalMux I__944 (
            .O(N__8731),
            .I(N__8720));
    LocalMux I__943 (
            .O(N__8728),
            .I(N__8715));
    LocalMux I__942 (
            .O(N__8723),
            .I(N__8715));
    Odrv12 I__941 (
            .O(N__8720),
            .I(\c0.rx.r_Clock_CountZ1Z_3 ));
    Odrv4 I__940 (
            .O(N__8715),
            .I(\c0.rx.r_Clock_CountZ1Z_3 ));
    InMux I__939 (
            .O(N__8710),
            .I(N__8700));
    InMux I__938 (
            .O(N__8709),
            .I(N__8700));
    InMux I__937 (
            .O(N__8708),
            .I(N__8697));
    InMux I__936 (
            .O(N__8707),
            .I(N__8690));
    InMux I__935 (
            .O(N__8706),
            .I(N__8690));
    InMux I__934 (
            .O(N__8705),
            .I(N__8690));
    LocalMux I__933 (
            .O(N__8700),
            .I(N__8687));
    LocalMux I__932 (
            .O(N__8697),
            .I(N__8682));
    LocalMux I__931 (
            .O(N__8690),
            .I(N__8682));
    Odrv4 I__930 (
            .O(N__8687),
            .I(\c0.rx.N_386 ));
    Odrv4 I__929 (
            .O(N__8682),
            .I(\c0.rx.N_386 ));
    InMux I__928 (
            .O(N__8677),
            .I(N__8669));
    InMux I__927 (
            .O(N__8676),
            .I(N__8662));
    InMux I__926 (
            .O(N__8675),
            .I(N__8662));
    InMux I__925 (
            .O(N__8674),
            .I(N__8662));
    InMux I__924 (
            .O(N__8673),
            .I(N__8657));
    InMux I__923 (
            .O(N__8672),
            .I(N__8657));
    LocalMux I__922 (
            .O(N__8669),
            .I(\c0.rx.r_SM_Main_dup_3 ));
    LocalMux I__921 (
            .O(N__8662),
            .I(\c0.rx.r_SM_Main_dup_3 ));
    LocalMux I__920 (
            .O(N__8657),
            .I(\c0.rx.r_SM_Main_dup_3 ));
    CascadeMux I__919 (
            .O(N__8650),
            .I(N__8641));
    InMux I__918 (
            .O(N__8649),
            .I(N__8636));
    InMux I__917 (
            .O(N__8648),
            .I(N__8636));
    InMux I__916 (
            .O(N__8647),
            .I(N__8627));
    InMux I__915 (
            .O(N__8646),
            .I(N__8627));
    InMux I__914 (
            .O(N__8645),
            .I(N__8620));
    InMux I__913 (
            .O(N__8644),
            .I(N__8620));
    InMux I__912 (
            .O(N__8641),
            .I(N__8617));
    LocalMux I__911 (
            .O(N__8636),
            .I(N__8614));
    InMux I__910 (
            .O(N__8635),
            .I(N__8607));
    InMux I__909 (
            .O(N__8634),
            .I(N__8607));
    InMux I__908 (
            .O(N__8633),
            .I(N__8607));
    InMux I__907 (
            .O(N__8632),
            .I(N__8604));
    LocalMux I__906 (
            .O(N__8627),
            .I(N__8601));
    InMux I__905 (
            .O(N__8626),
            .I(N__8596));
    InMux I__904 (
            .O(N__8625),
            .I(N__8596));
    LocalMux I__903 (
            .O(N__8620),
            .I(\c0.rx.N_98_dup ));
    LocalMux I__902 (
            .O(N__8617),
            .I(\c0.rx.N_98_dup ));
    Odrv12 I__901 (
            .O(N__8614),
            .I(\c0.rx.N_98_dup ));
    LocalMux I__900 (
            .O(N__8607),
            .I(\c0.rx.N_98_dup ));
    LocalMux I__899 (
            .O(N__8604),
            .I(\c0.rx.N_98_dup ));
    Odrv4 I__898 (
            .O(N__8601),
            .I(\c0.rx.N_98_dup ));
    LocalMux I__897 (
            .O(N__8596),
            .I(\c0.rx.N_98_dup ));
    InMux I__896 (
            .O(N__8581),
            .I(N__8576));
    InMux I__895 (
            .O(N__8580),
            .I(N__8571));
    InMux I__894 (
            .O(N__8579),
            .I(N__8571));
    LocalMux I__893 (
            .O(N__8576),
            .I(N__8561));
    LocalMux I__892 (
            .O(N__8571),
            .I(N__8561));
    InMux I__891 (
            .O(N__8570),
            .I(N__8556));
    InMux I__890 (
            .O(N__8569),
            .I(N__8556));
    InMux I__889 (
            .O(N__8568),
            .I(N__8553));
    InMux I__888 (
            .O(N__8567),
            .I(N__8548));
    InMux I__887 (
            .O(N__8566),
            .I(N__8548));
    Span4Mux_v I__886 (
            .O(N__8561),
            .I(N__8545));
    LocalMux I__885 (
            .O(N__8556),
            .I(N__8542));
    LocalMux I__884 (
            .O(N__8553),
            .I(\c0.rx.r_SM_Main_dup_4 ));
    LocalMux I__883 (
            .O(N__8548),
            .I(\c0.rx.r_SM_Main_dup_4 ));
    Odrv4 I__882 (
            .O(N__8545),
            .I(\c0.rx.r_SM_Main_dup_4 ));
    Odrv4 I__881 (
            .O(N__8542),
            .I(\c0.rx.r_SM_Main_dup_4 ));
    CascadeMux I__880 (
            .O(N__8533),
            .I(\c0.rx.N_138r_0_i_1_cascade_ ));
    CascadeMux I__879 (
            .O(N__8530),
            .I(N__8527));
    InMux I__878 (
            .O(N__8527),
            .I(N__8521));
    CascadeMux I__877 (
            .O(N__8526),
            .I(N__8516));
    CascadeMux I__876 (
            .O(N__8525),
            .I(N__8513));
    InMux I__875 (
            .O(N__8524),
            .I(N__8509));
    LocalMux I__874 (
            .O(N__8521),
            .I(N__8506));
    InMux I__873 (
            .O(N__8520),
            .I(N__8501));
    InMux I__872 (
            .O(N__8519),
            .I(N__8501));
    InMux I__871 (
            .O(N__8516),
            .I(N__8494));
    InMux I__870 (
            .O(N__8513),
            .I(N__8494));
    InMux I__869 (
            .O(N__8512),
            .I(N__8494));
    LocalMux I__868 (
            .O(N__8509),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    Odrv4 I__867 (
            .O(N__8506),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    LocalMux I__866 (
            .O(N__8501),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    LocalMux I__865 (
            .O(N__8494),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    CascadeMux I__864 (
            .O(N__8485),
            .I(\c0.rx.N_91_0_cascade_ ));
    InMux I__863 (
            .O(N__8482),
            .I(N__8479));
    LocalMux I__862 (
            .O(N__8479),
            .I(\c0.rx.r_SM_Main_illegal_0 ));
    CascadeMux I__861 (
            .O(N__8476),
            .I(\c0.rx.r_SM_Main_ns_0_i_a2_0_3_cascade_ ));
    CascadeMux I__860 (
            .O(N__8473),
            .I(\c0.rx.N_320_cascade_ ));
    CascadeMux I__859 (
            .O(N__8470),
            .I(\c0.rx.r_Clock_Count_8_f0_0_o2_0_2_cascade_ ));
    CascadeMux I__858 (
            .O(N__8467),
            .I(N__8463));
    InMux I__857 (
            .O(N__8466),
            .I(N__8460));
    InMux I__856 (
            .O(N__8463),
            .I(N__8457));
    LocalMux I__855 (
            .O(N__8460),
            .I(\c0.rx.un1_r_Clock_Count_2_sqmuxa_0_i ));
    LocalMux I__854 (
            .O(N__8457),
            .I(\c0.rx.un1_r_Clock_Count_2_sqmuxa_0_i ));
    CascadeMux I__853 (
            .O(N__8452),
            .I(N__8449));
    InMux I__852 (
            .O(N__8449),
            .I(N__8446));
    LocalMux I__851 (
            .O(N__8446),
            .I(\c0.rx.r_Clock_Count_8_f0_0_o2_0_2 ));
    InMux I__850 (
            .O(N__8443),
            .I(N__8440));
    LocalMux I__849 (
            .O(N__8440),
            .I(\c0.rx.r_Clock_Count_RNO_0_0_2 ));
    CascadeMux I__848 (
            .O(N__8437),
            .I(\c0.rx.N_332_cascade_ ));
    InMux I__847 (
            .O(N__8434),
            .I(N__8430));
    InMux I__846 (
            .O(N__8433),
            .I(N__8427));
    LocalMux I__845 (
            .O(N__8430),
            .I(\c0.rx.r_Clock_CountZ1Z_2 ));
    LocalMux I__844 (
            .O(N__8427),
            .I(\c0.rx.r_Clock_CountZ1Z_2 ));
    InMux I__843 (
            .O(N__8422),
            .I(N__8418));
    InMux I__842 (
            .O(N__8421),
            .I(N__8415));
    LocalMux I__841 (
            .O(N__8418),
            .I(\c0.rx.r_Clock_CountZ1Z_6 ));
    LocalMux I__840 (
            .O(N__8415),
            .I(\c0.rx.r_Clock_CountZ1Z_6 ));
    CascadeMux I__839 (
            .O(N__8410),
            .I(N__8406));
    InMux I__838 (
            .O(N__8409),
            .I(N__8403));
    InMux I__837 (
            .O(N__8406),
            .I(N__8400));
    LocalMux I__836 (
            .O(N__8403),
            .I(\c0.rx.r_Clock_CountZ0Z_7 ));
    LocalMux I__835 (
            .O(N__8400),
            .I(\c0.rx.r_Clock_CountZ0Z_7 ));
    InMux I__834 (
            .O(N__8395),
            .I(N__8391));
    InMux I__833 (
            .O(N__8394),
            .I(N__8388));
    LocalMux I__832 (
            .O(N__8391),
            .I(\c0.rx.r_Clock_CountZ1Z_4 ));
    LocalMux I__831 (
            .O(N__8388),
            .I(\c0.rx.r_Clock_CountZ1Z_4 ));
    InMux I__830 (
            .O(N__8383),
            .I(N__8380));
    LocalMux I__829 (
            .O(N__8380),
            .I(\c0.rx.r_Clock_Count_RNO_0Z0Z_5 ));
    InMux I__828 (
            .O(N__8377),
            .I(N__8373));
    InMux I__827 (
            .O(N__8376),
            .I(N__8370));
    LocalMux I__826 (
            .O(N__8373),
            .I(\c0.rx.r_Clock_CountZ1Z_5 ));
    LocalMux I__825 (
            .O(N__8370),
            .I(\c0.rx.r_Clock_CountZ1Z_5 ));
    InMux I__824 (
            .O(N__8365),
            .I(N__8361));
    InMux I__823 (
            .O(N__8364),
            .I(N__8358));
    LocalMux I__822 (
            .O(N__8361),
            .I(\c0.rx.N_320 ));
    LocalMux I__821 (
            .O(N__8358),
            .I(\c0.rx.N_320 ));
    InMux I__820 (
            .O(N__8353),
            .I(N__8348));
    InMux I__819 (
            .O(N__8352),
            .I(N__8343));
    InMux I__818 (
            .O(N__8351),
            .I(N__8343));
    LocalMux I__817 (
            .O(N__8348),
            .I(\c0.rx.N_317 ));
    LocalMux I__816 (
            .O(N__8343),
            .I(\c0.rx.N_317 ));
    InMux I__815 (
            .O(N__8338),
            .I(N__8335));
    LocalMux I__814 (
            .O(N__8335),
            .I(\c0.rx.N_337 ));
    CascadeMux I__813 (
            .O(N__8332),
            .I(\c0.rx.N_383_cascade_ ));
    InMux I__812 (
            .O(N__8329),
            .I(N__8326));
    LocalMux I__811 (
            .O(N__8326),
            .I(\c0.rx.r_Clock_Count_RNO_0_0_1 ));
    InMux I__810 (
            .O(N__8323),
            .I(\c0.rx.un1_r_Clock_Count_5_cry_0 ));
    InMux I__809 (
            .O(N__8320),
            .I(\c0.rx.un1_r_Clock_Count_5_cry_1 ));
    InMux I__808 (
            .O(N__8317),
            .I(\c0.rx.un1_r_Clock_Count_5_cry_2 ));
    InMux I__807 (
            .O(N__8314),
            .I(N__8311));
    LocalMux I__806 (
            .O(N__8311),
            .I(\c0.rx.r_Clock_Count_RNO_0Z0Z_4 ));
    InMux I__805 (
            .O(N__8308),
            .I(\c0.rx.un1_r_Clock_Count_5_cry_3 ));
    InMux I__804 (
            .O(N__8305),
            .I(\c0.rx.un1_r_Clock_Count_5_cry_4 ));
    InMux I__803 (
            .O(N__8302),
            .I(N__8299));
    LocalMux I__802 (
            .O(N__8299),
            .I(\c0.rx.r_Clock_Count_RNO_0Z0Z_6 ));
    InMux I__801 (
            .O(N__8296),
            .I(\c0.rx.un1_r_Clock_Count_5_cry_5 ));
    InMux I__800 (
            .O(N__8293),
            .I(\c0.rx.un1_r_Clock_Count_5_cry_6 ));
    InMux I__799 (
            .O(N__8290),
            .I(N__8287));
    LocalMux I__798 (
            .O(N__8287),
            .I(\c0.rx.r_Clock_Count_RNO_0Z0Z_7 ));
    InMux I__797 (
            .O(N__8284),
            .I(N__8280));
    InMux I__796 (
            .O(N__8283),
            .I(N__8277));
    LocalMux I__795 (
            .O(N__8280),
            .I(\c0.rx.r_Clock_CountZ1Z_1 ));
    LocalMux I__794 (
            .O(N__8277),
            .I(\c0.rx.r_Clock_CountZ1Z_1 ));
    InMux I__793 (
            .O(N__8272),
            .I(N__8268));
    InMux I__792 (
            .O(N__8271),
            .I(N__8265));
    LocalMux I__791 (
            .O(N__8268),
            .I(\c0.rx.r_Clock_CountZ1Z_0 ));
    LocalMux I__790 (
            .O(N__8265),
            .I(\c0.rx.r_Clock_CountZ1Z_0 ));
    CascadeMux I__789 (
            .O(N__8260),
            .I(\c0.rx.r_Rx_Bytece_0_5_cascade_ ));
    InMux I__788 (
            .O(N__8257),
            .I(N__8252));
    InMux I__787 (
            .O(N__8256),
            .I(N__8249));
    InMux I__786 (
            .O(N__8255),
            .I(N__8246));
    LocalMux I__785 (
            .O(N__8252),
            .I(\c0.rx.N_388 ));
    LocalMux I__784 (
            .O(N__8249),
            .I(\c0.rx.N_388 ));
    LocalMux I__783 (
            .O(N__8246),
            .I(\c0.rx.N_388 ));
    CascadeMux I__782 (
            .O(N__8239),
            .I(\c0.rx.r_Rx_Bytece_0_6_cascade_ ));
    InMux I__781 (
            .O(N__8236),
            .I(N__8227));
    InMux I__780 (
            .O(N__8235),
            .I(N__8224));
    InMux I__779 (
            .O(N__8234),
            .I(N__8221));
    InMux I__778 (
            .O(N__8233),
            .I(N__8216));
    InMux I__777 (
            .O(N__8232),
            .I(N__8216));
    InMux I__776 (
            .O(N__8231),
            .I(N__8211));
    InMux I__775 (
            .O(N__8230),
            .I(N__8211));
    LocalMux I__774 (
            .O(N__8227),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    LocalMux I__773 (
            .O(N__8224),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    LocalMux I__772 (
            .O(N__8221),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    LocalMux I__771 (
            .O(N__8216),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    LocalMux I__770 (
            .O(N__8211),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    InMux I__769 (
            .O(N__8200),
            .I(N__8197));
    LocalMux I__768 (
            .O(N__8197),
            .I(\c0.rx.r_Rx_Bytece_0_0 ));
    CascadeMux I__767 (
            .O(N__8194),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa_cascade_ ));
    InMux I__766 (
            .O(N__8191),
            .I(N__8188));
    LocalMux I__765 (
            .O(N__8188),
            .I(\c0.rx.r_Clock_Count_RNO_0_0_0 ));
    InMux I__764 (
            .O(N__8185),
            .I(blink_counter_cry_20));
    InMux I__763 (
            .O(N__8182),
            .I(blink_counter_cry_21));
    InMux I__762 (
            .O(N__8179),
            .I(blink_counter_cry_22));
    InMux I__761 (
            .O(N__8176),
            .I(bfn_6_24_0_));
    InMux I__760 (
            .O(N__8173),
            .I(blink_counter_cry_24));
    CascadeMux I__759 (
            .O(N__8170),
            .I(\c0.rx.r_Rx_Bytece_0_2_cascade_ ));
    InMux I__758 (
            .O(N__8167),
            .I(N__8164));
    LocalMux I__757 (
            .O(N__8164),
            .I(\c0.rx.N_325 ));
    CascadeMux I__756 (
            .O(N__8161),
            .I(\c0.rx.N_325_cascade_ ));
    InMux I__755 (
            .O(N__8158),
            .I(N__8155));
    LocalMux I__754 (
            .O(N__8155),
            .I(blink_counterZ0Z_13));
    InMux I__753 (
            .O(N__8152),
            .I(blink_counter_cry_12));
    InMux I__752 (
            .O(N__8149),
            .I(N__8146));
    LocalMux I__751 (
            .O(N__8146),
            .I(blink_counterZ0Z_14));
    InMux I__750 (
            .O(N__8143),
            .I(blink_counter_cry_13));
    InMux I__749 (
            .O(N__8140),
            .I(N__8137));
    LocalMux I__748 (
            .O(N__8137),
            .I(blink_counterZ0Z_15));
    InMux I__747 (
            .O(N__8134),
            .I(blink_counter_cry_14));
    InMux I__746 (
            .O(N__8131),
            .I(N__8128));
    LocalMux I__745 (
            .O(N__8128),
            .I(blink_counterZ0Z_16));
    InMux I__744 (
            .O(N__8125),
            .I(bfn_6_23_0_));
    InMux I__743 (
            .O(N__8122),
            .I(N__8119));
    LocalMux I__742 (
            .O(N__8119),
            .I(blink_counterZ0Z_17));
    InMux I__741 (
            .O(N__8116),
            .I(blink_counter_cry_16));
    InMux I__740 (
            .O(N__8113),
            .I(N__8110));
    LocalMux I__739 (
            .O(N__8110),
            .I(blink_counterZ0Z_18));
    InMux I__738 (
            .O(N__8107),
            .I(blink_counter_cry_17));
    InMux I__737 (
            .O(N__8104),
            .I(N__8101));
    LocalMux I__736 (
            .O(N__8101),
            .I(blink_counterZ0Z_19));
    InMux I__735 (
            .O(N__8098),
            .I(blink_counter_cry_18));
    InMux I__734 (
            .O(N__8095),
            .I(N__8092));
    LocalMux I__733 (
            .O(N__8092),
            .I(blink_counterZ0Z_20));
    InMux I__732 (
            .O(N__8089),
            .I(blink_counter_cry_19));
    InMux I__731 (
            .O(N__8086),
            .I(N__8083));
    LocalMux I__730 (
            .O(N__8083),
            .I(blink_counterZ0Z_4));
    InMux I__729 (
            .O(N__8080),
            .I(blink_counter_cry_3));
    InMux I__728 (
            .O(N__8077),
            .I(N__8074));
    LocalMux I__727 (
            .O(N__8074),
            .I(blink_counterZ0Z_5));
    InMux I__726 (
            .O(N__8071),
            .I(blink_counter_cry_4));
    InMux I__725 (
            .O(N__8068),
            .I(N__8065));
    LocalMux I__724 (
            .O(N__8065),
            .I(blink_counterZ0Z_6));
    InMux I__723 (
            .O(N__8062),
            .I(blink_counter_cry_5));
    InMux I__722 (
            .O(N__8059),
            .I(N__8056));
    LocalMux I__721 (
            .O(N__8056),
            .I(blink_counterZ0Z_7));
    InMux I__720 (
            .O(N__8053),
            .I(blink_counter_cry_6));
    InMux I__719 (
            .O(N__8050),
            .I(N__8047));
    LocalMux I__718 (
            .O(N__8047),
            .I(blink_counterZ0Z_8));
    InMux I__717 (
            .O(N__8044),
            .I(bfn_6_22_0_));
    InMux I__716 (
            .O(N__8041),
            .I(N__8038));
    LocalMux I__715 (
            .O(N__8038),
            .I(blink_counterZ0Z_9));
    InMux I__714 (
            .O(N__8035),
            .I(blink_counter_cry_8));
    InMux I__713 (
            .O(N__8032),
            .I(N__8029));
    LocalMux I__712 (
            .O(N__8029),
            .I(blink_counterZ0Z_10));
    InMux I__711 (
            .O(N__8026),
            .I(blink_counter_cry_9));
    InMux I__710 (
            .O(N__8023),
            .I(N__8020));
    LocalMux I__709 (
            .O(N__8020),
            .I(blink_counterZ0Z_11));
    InMux I__708 (
            .O(N__8017),
            .I(blink_counter_cry_10));
    InMux I__707 (
            .O(N__8014),
            .I(N__8011));
    LocalMux I__706 (
            .O(N__8011),
            .I(blink_counterZ0Z_12));
    InMux I__705 (
            .O(N__8008),
            .I(blink_counter_cry_11));
    CascadeMux I__704 (
            .O(N__8005),
            .I(\c0.rx.r_SM_Main_RNI58REZ0Z_0_cascade_ ));
    IoInMux I__703 (
            .O(N__8002),
            .I(N__7999));
    LocalMux I__702 (
            .O(N__7999),
            .I(N__7996));
    Span4Mux_s1_h I__701 (
            .O(N__7996),
            .I(N__7993));
    Span4Mux_h I__700 (
            .O(N__7993),
            .I(N__7990));
    Odrv4 I__699 (
            .O(N__7990),
            .I(\c0.rx.rx_data_ready ));
    InMux I__698 (
            .O(N__7987),
            .I(N__7984));
    LocalMux I__697 (
            .O(N__7984),
            .I(blink_counterZ0Z_0));
    InMux I__696 (
            .O(N__7981),
            .I(bfn_6_21_0_));
    InMux I__695 (
            .O(N__7978),
            .I(N__7975));
    LocalMux I__694 (
            .O(N__7975),
            .I(blink_counterZ0Z_1));
    InMux I__693 (
            .O(N__7972),
            .I(blink_counter_cry_0));
    InMux I__692 (
            .O(N__7969),
            .I(N__7966));
    LocalMux I__691 (
            .O(N__7966),
            .I(blink_counterZ0Z_2));
    InMux I__690 (
            .O(N__7963),
            .I(blink_counter_cry_1));
    InMux I__689 (
            .O(N__7960),
            .I(N__7957));
    LocalMux I__688 (
            .O(N__7957),
            .I(blink_counterZ0Z_3));
    InMux I__687 (
            .O(N__7954),
            .I(blink_counter_cry_2));
    CascadeMux I__686 (
            .O(N__7951),
            .I(\c0.rx.N_336_cascade_ ));
    InMux I__685 (
            .O(N__7948),
            .I(N__7945));
    LocalMux I__684 (
            .O(N__7945),
            .I(\c0.rx.r_Rx_Bytece_0_1 ));
    InMux I__683 (
            .O(N__7942),
            .I(N__7938));
    InMux I__682 (
            .O(N__7941),
            .I(N__7935));
    LocalMux I__681 (
            .O(N__7938),
            .I(\c0.tx.r_Clock_Count_i_0 ));
    LocalMux I__680 (
            .O(N__7935),
            .I(\c0.tx.r_Clock_Count_i_0 ));
    CascadeMux I__679 (
            .O(N__7930),
            .I(\c0.rx.r_Rx_Bytece_0_4_cascade_ ));
    InMux I__678 (
            .O(N__7927),
            .I(N__7924));
    LocalMux I__677 (
            .O(N__7924),
            .I(N__7921));
    Span4Mux_v I__676 (
            .O(N__7921),
            .I(N__7918));
    Span4Mux_v I__675 (
            .O(N__7918),
            .I(N__7915));
    Span4Mux_v I__674 (
            .O(N__7915),
            .I(N__7912));
    Odrv4 I__673 (
            .O(N__7912),
            .I(PIN_2_c));
    InMux I__672 (
            .O(N__7909),
            .I(N__7906));
    LocalMux I__671 (
            .O(N__7906),
            .I(N__7903));
    Span4Mux_h I__670 (
            .O(N__7903),
            .I(N__7900));
    Odrv4 I__669 (
            .O(N__7900),
            .I(\c0.rx.r_Rx_Data_RZ0 ));
    InMux I__668 (
            .O(N__7897),
            .I(N__7894));
    LocalMux I__667 (
            .O(N__7894),
            .I(\c0.tx.r_Clock_Count_i_1 ));
    InMux I__666 (
            .O(N__7891),
            .I(N__7888));
    LocalMux I__665 (
            .O(N__7888),
            .I(\c0.tx.r_Clock_Count_i_2 ));
    InMux I__664 (
            .O(N__7885),
            .I(N__7882));
    LocalMux I__663 (
            .O(N__7882),
            .I(\c0.tx.r_Clock_Count_i_3 ));
    InMux I__662 (
            .O(N__7879),
            .I(\c0.tx.r_Clock_Count12 ));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_5_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_22_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\c0.i12 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\c0.data_cry_7 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_6_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_21_0_));
    defparam IN_MUX_bfv_6_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_22_0_ (
            .carryinitin(blink_counter_cry_7),
            .carryinitout(bfn_6_22_0_));
    defparam IN_MUX_bfv_6_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_23_0_ (
            .carryinitin(blink_counter_cry_15),
            .carryinitout(bfn_6_23_0_));
    defparam IN_MUX_bfv_6_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_24_0_ (
            .carryinitin(blink_counter_cry_23),
            .carryinitout(bfn_6_24_0_));
    ICE_GB \c0.rx.r_Rx_DV_RNID002  (
            .USERSIGNALTOGLOBALBUFFER(N__8002),
            .GLOBALBUFFEROUTPUT(\c0.rx_data_ready_g ));
    ICE_GB \c0.byte_transmit_counter_RNI4QES5_0_2  (
            .USERSIGNALTOGLOBALBUFFER(N__15046),
            .GLOBALBUFFEROUTPUT(\c0.data_out_0__1_sqmuxa_g ));
    ICE_GB \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_0  (
            .USERSIGNALTOGLOBALBUFFER(N__19270),
            .GLOBALBUFFEROUTPUT(\c0.data_in_frame_0__0_sqmuxa_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_R_LC_1_13_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_R_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_R_LC_1_13_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.rx.r_Rx_Data_R_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__7927),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.rx.r_Rx_Data_RZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19578),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_LC_4_16_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_LC_4_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_LC_4_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7909),
            .lcout(\c0.rx.r_Rx_DataZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_0_c_LC_5_22_0 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count12_cry_0_c_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_0_c_LC_5_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_0_c_LC_5_22_0  (
            .in0(_gnd_net_),
            .in1(N__7941),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_22_0_),
            .carryout(\c0.tx.r_Clock_Count12_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_5_22_1 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_5_22_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_5_22_1  (
            .in0(N__9464),
            .in1(N__7897),
            .in2(N__17115),
            .in3(_gnd_net_),
            .lcout(\c0.tx.r_Clock_Count_i_1 ),
            .ltout(),
            .carryin(\c0.tx.r_Clock_Count12_cry_0 ),
            .carryout(\c0.tx.r_Clock_Count12_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_5_22_2 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_5_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_5_22_2  (
            .in0(_gnd_net_),
            .in1(N__7891),
            .in2(N__17092),
            .in3(N__9485),
            .lcout(\c0.tx.r_Clock_Count_i_2 ),
            .ltout(),
            .carryin(\c0.tx.r_Clock_Count12_cry_1 ),
            .carryout(\c0.tx.r_Clock_Count12_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_5_22_3 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_5_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(N__7885),
            .in2(N__17116),
            .in3(N__9438),
            .lcout(\c0.tx.r_Clock_Count_i_3 ),
            .ltout(),
            .carryin(\c0.tx.r_Clock_Count12_cry_2 ),
            .carryout(\c0.tx.r_Clock_Count12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_5_22_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_5_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_5_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7879),
            .lcout(\c0.tx.r_Clock_Count12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__0_LC_5_22_6 .C_ON=1'b0;
    defparam \c0.data_out_1__0_LC_5_22_6 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__0_LC_5_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_1__0_LC_5_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17104),
            .lcout(\c0.d_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19587),
            .ce(),
            .sr(N__16882));
    defparam \c0.data_out_3__3_LC_5_22_7 .C_ON=1'b0;
    defparam \c0.data_out_3__3_LC_5_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__3_LC_5_22_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_3__3_LC_5_22_7  (
            .in0(N__17105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19587),
            .ce(),
            .sr(N__16882));
    defparam \c0.tx.r_SM_Main_RNO_0_1_LC_5_23_1 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNO_0_1_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNO_0_1_LC_5_23_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \c0.tx.r_SM_Main_RNO_0_1_LC_5_23_1  (
            .in0(N__9958),
            .in1(N__9876),
            .in2(_gnd_net_),
            .in3(N__10539),
            .lcout(\c0.tx.r_SM_Main_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_0_LC_5_23_2 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_0_LC_5_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count_0_LC_5_23_2 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \c0.tx.r_Clock_Count_0_LC_5_23_2  (
            .in0(N__9877),
            .in1(N__9334),
            .in2(N__10368),
            .in3(N__9768),
            .lcout(\c0.tx.r_Clock_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_23_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_23_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_23_3  (
            .in0(N__17056),
            .in1(N__9420),
            .in2(_gnd_net_),
            .in3(N__7942),
            .lcout(\c0.tx.r_Clock_Count_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_1_LC_5_23_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_1_LC_5_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count_1_LC_5_23_4 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \c0.tx.r_Clock_Count_1_LC_5_23_4  (
            .in0(N__9878),
            .in1(N__9322),
            .in2(N__10369),
            .in3(N__9769),
            .lcout(\c0.tx.r_Clock_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_2_LC_5_23_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_2_LC_5_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count_2_LC_5_23_5 .LUT_INIT=16'b1100111000000000;
    LogicCell40 \c0.tx.r_Clock_Count_2_LC_5_23_5  (
            .in0(N__9766),
            .in1(N__10360),
            .in2(N__9883),
            .in3(N__9517),
            .lcout(\c0.tx.r_Clock_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_3_LC_5_23_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_3_LC_5_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count_3_LC_5_23_6 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \c0.tx.r_Clock_Count_3_LC_5_23_6  (
            .in0(N__9879),
            .in1(N__9767),
            .in2(N__10367),
            .in3(N__9502),
            .lcout(\c0.tx.r_Clock_CountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_4_LC_6_17_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_4_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_4_LC_6_17_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_4_LC_6_17_3  (
            .in0(N__14233),
            .in1(N__14112),
            .in2(_gnd_net_),
            .in3(N__14178),
            .lcout(),
            .ltout(\c0.rx.r_Rx_Bytece_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_4_LC_6_17_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_4_LC_6_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_4_LC_6_17_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \c0.rx.r_Rx_Byte_4_LC_6_17_4  (
            .in0(N__9046),
            .in1(N__12228),
            .in2(N__7930),
            .in3(N__8235),
            .lcout(\c0.rx_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_1_LC_6_17_5 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_1_LC_6_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_1_LC_6_17_5 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \c0.rx.r_Bit_Index_1_LC_6_17_5  (
            .in0(N__14117),
            .in1(N__8256),
            .in2(N__14246),
            .in3(N__8849),
            .lcout(\c0.rx.r_Bit_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_0_LC_6_18_0 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_0_LC_6_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_0_LC_6_18_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \c0.rx.r_Bit_Index_0_LC_6_18_0  (
            .in0(N__14116),
            .in1(N__8255),
            .in2(_gnd_net_),
            .in3(N__8848),
            .lcout(\c0.rx.r_Bit_IndexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19582),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_3_LC_6_18_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_3_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_3_LC_6_18_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_3_LC_6_18_2  (
            .in0(_gnd_net_),
            .in1(N__14173),
            .in2(_gnd_net_),
            .in3(N__8167),
            .lcout(),
            .ltout(\c0.rx.N_336_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_3_LC_6_18_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_3_LC_6_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_3_LC_6_18_3 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.rx.r_Rx_Byte_3_LC_6_18_3  (
            .in0(N__10218),
            .in1(N__9048),
            .in2(N__7951),
            .in3(N__8236),
            .lcout(\c0.rx_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19582),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_1_LC_6_18_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_1_LC_6_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_1_LC_6_18_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_1_LC_6_18_4  (
            .in0(N__14227),
            .in1(N__14174),
            .in2(_gnd_net_),
            .in3(N__14109),
            .lcout(\c0.rx.r_Rx_Bytece_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_6_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_6_LC_6_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_6_LC_6_19_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.rx.r_Clock_Count_6_LC_6_19_0  (
            .in0(N__8886),
            .in1(N__8832),
            .in2(N__8788),
            .in3(N__8302),
            .lcout(\c0.rx.r_Clock_CountZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_1_LC_6_19_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_1_LC_6_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_1_LC_6_19_1 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \c0.rx.r_Clock_Count_1_LC_6_19_1  (
            .in0(N__8830),
            .in1(N__8884),
            .in2(N__8919),
            .in3(N__8329),
            .lcout(\c0.rx.r_Clock_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_1_LC_6_19_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_1_LC_6_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_1_LC_6_19_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_1_LC_6_19_3  (
            .in0(N__7948),
            .in1(N__9044),
            .in2(N__10203),
            .in3(N__8234),
            .lcout(\c0.rx_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_4_LC_6_19_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_4_LC_6_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_4_LC_6_19_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.rx.r_Clock_Count_4_LC_6_19_4  (
            .in0(N__8885),
            .in1(N__8831),
            .in2(N__8787),
            .in3(N__8314),
            .lcout(\c0.rx.r_Clock_CountZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_0_LC_6_19_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_0_LC_6_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_0_LC_6_19_6 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \c0.rx.r_Clock_Count_0_LC_6_19_6  (
            .in0(N__8883),
            .in1(N__8829),
            .in2(N__8920),
            .in3(N__8191),
            .lcout(\c0.rx.r_Clock_CountZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNO_0_1_LC_6_20_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNO_0_1_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNO_0_1_LC_6_20_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \c0.rx.r_SM_Main_RNO_0_1_LC_6_20_0  (
            .in0(N__8520),
            .in1(N__9045),
            .in2(_gnd_net_),
            .in3(N__9145),
            .lcout(\c0.rx.N_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNI58RE_0_LC_6_20_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNI58RE_0_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNI58RE_0_LC_6_20_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.r_SM_Main_RNI58RE_0_LC_6_20_1  (
            .in0(_gnd_net_),
            .in1(N__8632),
            .in2(_gnd_net_),
            .in3(N__8519),
            .lcout(\c0.rx.r_SM_Main_RNI58REZ0Z_0 ),
            .ltout(\c0.rx.r_SM_Main_RNI58REZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_7_LC_6_20_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_7_LC_6_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_7_LC_6_20_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.rx.r_Clock_Count_7_LC_6_20_2  (
            .in0(N__8779),
            .in1(N__8882),
            .in2(N__8005),
            .in3(N__8290),
            .lcout(\c0.rx.r_Clock_CountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19585),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_LC_6_20_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_LC_6_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_LC_6_20_7 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \c0.rx.r_Rx_DV_LC_6_20_7  (
            .in0(N__8847),
            .in1(N__9115),
            .in2(N__17734),
            .in3(N__8581),
            .lcout(\c0.rx.rx_data_ready ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19585),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_0_LC_6_21_0.C_ON=1'b1;
    defparam blink_counter_0_LC_6_21_0.SEQ_MODE=4'b1000;
    defparam blink_counter_0_LC_6_21_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_0_LC_6_21_0 (
            .in0(_gnd_net_),
            .in1(N__7987),
            .in2(_gnd_net_),
            .in3(N__7981),
            .lcout(blink_counterZ0Z_0),
            .ltout(),
            .carryin(bfn_6_21_0_),
            .carryout(blink_counter_cry_0),
            .clk(N__19588),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1_LC_6_21_1.C_ON=1'b1;
    defparam blink_counter_1_LC_6_21_1.SEQ_MODE=4'b1000;
    defparam blink_counter_1_LC_6_21_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_1_LC_6_21_1 (
            .in0(_gnd_net_),
            .in1(N__7978),
            .in2(_gnd_net_),
            .in3(N__7972),
            .lcout(blink_counterZ0Z_1),
            .ltout(),
            .carryin(blink_counter_cry_0),
            .carryout(blink_counter_cry_1),
            .clk(N__19588),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2_LC_6_21_2.C_ON=1'b1;
    defparam blink_counter_2_LC_6_21_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2_LC_6_21_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_2_LC_6_21_2 (
            .in0(_gnd_net_),
            .in1(N__7969),
            .in2(_gnd_net_),
            .in3(N__7963),
            .lcout(blink_counterZ0Z_2),
            .ltout(),
            .carryin(blink_counter_cry_1),
            .carryout(blink_counter_cry_2),
            .clk(N__19588),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_3_LC_6_21_3.C_ON=1'b1;
    defparam blink_counter_3_LC_6_21_3.SEQ_MODE=4'b1000;
    defparam blink_counter_3_LC_6_21_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_3_LC_6_21_3 (
            .in0(_gnd_net_),
            .in1(N__7960),
            .in2(_gnd_net_),
            .in3(N__7954),
            .lcout(blink_counterZ0Z_3),
            .ltout(),
            .carryin(blink_counter_cry_2),
            .carryout(blink_counter_cry_3),
            .clk(N__19588),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_4_LC_6_21_4.C_ON=1'b1;
    defparam blink_counter_4_LC_6_21_4.SEQ_MODE=4'b1000;
    defparam blink_counter_4_LC_6_21_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_4_LC_6_21_4 (
            .in0(_gnd_net_),
            .in1(N__8086),
            .in2(_gnd_net_),
            .in3(N__8080),
            .lcout(blink_counterZ0Z_4),
            .ltout(),
            .carryin(blink_counter_cry_3),
            .carryout(blink_counter_cry_4),
            .clk(N__19588),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_5_LC_6_21_5.C_ON=1'b1;
    defparam blink_counter_5_LC_6_21_5.SEQ_MODE=4'b1000;
    defparam blink_counter_5_LC_6_21_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_5_LC_6_21_5 (
            .in0(_gnd_net_),
            .in1(N__8077),
            .in2(_gnd_net_),
            .in3(N__8071),
            .lcout(blink_counterZ0Z_5),
            .ltout(),
            .carryin(blink_counter_cry_4),
            .carryout(blink_counter_cry_5),
            .clk(N__19588),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_6_LC_6_21_6.C_ON=1'b1;
    defparam blink_counter_6_LC_6_21_6.SEQ_MODE=4'b1000;
    defparam blink_counter_6_LC_6_21_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_6_LC_6_21_6 (
            .in0(_gnd_net_),
            .in1(N__8068),
            .in2(_gnd_net_),
            .in3(N__8062),
            .lcout(blink_counterZ0Z_6),
            .ltout(),
            .carryin(blink_counter_cry_5),
            .carryout(blink_counter_cry_6),
            .clk(N__19588),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_7_LC_6_21_7.C_ON=1'b1;
    defparam blink_counter_7_LC_6_21_7.SEQ_MODE=4'b1000;
    defparam blink_counter_7_LC_6_21_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_7_LC_6_21_7 (
            .in0(_gnd_net_),
            .in1(N__8059),
            .in2(_gnd_net_),
            .in3(N__8053),
            .lcout(blink_counterZ0Z_7),
            .ltout(),
            .carryin(blink_counter_cry_6),
            .carryout(blink_counter_cry_7),
            .clk(N__19588),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_8_LC_6_22_0.C_ON=1'b1;
    defparam blink_counter_8_LC_6_22_0.SEQ_MODE=4'b1000;
    defparam blink_counter_8_LC_6_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_8_LC_6_22_0 (
            .in0(_gnd_net_),
            .in1(N__8050),
            .in2(_gnd_net_),
            .in3(N__8044),
            .lcout(blink_counterZ0Z_8),
            .ltout(),
            .carryin(bfn_6_22_0_),
            .carryout(blink_counter_cry_8),
            .clk(N__19595),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_9_LC_6_22_1.C_ON=1'b1;
    defparam blink_counter_9_LC_6_22_1.SEQ_MODE=4'b1000;
    defparam blink_counter_9_LC_6_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_9_LC_6_22_1 (
            .in0(_gnd_net_),
            .in1(N__8041),
            .in2(_gnd_net_),
            .in3(N__8035),
            .lcout(blink_counterZ0Z_9),
            .ltout(),
            .carryin(blink_counter_cry_8),
            .carryout(blink_counter_cry_9),
            .clk(N__19595),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_10_LC_6_22_2.C_ON=1'b1;
    defparam blink_counter_10_LC_6_22_2.SEQ_MODE=4'b1000;
    defparam blink_counter_10_LC_6_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_10_LC_6_22_2 (
            .in0(_gnd_net_),
            .in1(N__8032),
            .in2(_gnd_net_),
            .in3(N__8026),
            .lcout(blink_counterZ0Z_10),
            .ltout(),
            .carryin(blink_counter_cry_9),
            .carryout(blink_counter_cry_10),
            .clk(N__19595),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_11_LC_6_22_3.C_ON=1'b1;
    defparam blink_counter_11_LC_6_22_3.SEQ_MODE=4'b1000;
    defparam blink_counter_11_LC_6_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_11_LC_6_22_3 (
            .in0(_gnd_net_),
            .in1(N__8023),
            .in2(_gnd_net_),
            .in3(N__8017),
            .lcout(blink_counterZ0Z_11),
            .ltout(),
            .carryin(blink_counter_cry_10),
            .carryout(blink_counter_cry_11),
            .clk(N__19595),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_12_LC_6_22_4.C_ON=1'b1;
    defparam blink_counter_12_LC_6_22_4.SEQ_MODE=4'b1000;
    defparam blink_counter_12_LC_6_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_12_LC_6_22_4 (
            .in0(_gnd_net_),
            .in1(N__8014),
            .in2(_gnd_net_),
            .in3(N__8008),
            .lcout(blink_counterZ0Z_12),
            .ltout(),
            .carryin(blink_counter_cry_11),
            .carryout(blink_counter_cry_12),
            .clk(N__19595),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_13_LC_6_22_5.C_ON=1'b1;
    defparam blink_counter_13_LC_6_22_5.SEQ_MODE=4'b1000;
    defparam blink_counter_13_LC_6_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_13_LC_6_22_5 (
            .in0(_gnd_net_),
            .in1(N__8158),
            .in2(_gnd_net_),
            .in3(N__8152),
            .lcout(blink_counterZ0Z_13),
            .ltout(),
            .carryin(blink_counter_cry_12),
            .carryout(blink_counter_cry_13),
            .clk(N__19595),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_14_LC_6_22_6.C_ON=1'b1;
    defparam blink_counter_14_LC_6_22_6.SEQ_MODE=4'b1000;
    defparam blink_counter_14_LC_6_22_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_14_LC_6_22_6 (
            .in0(_gnd_net_),
            .in1(N__8149),
            .in2(_gnd_net_),
            .in3(N__8143),
            .lcout(blink_counterZ0Z_14),
            .ltout(),
            .carryin(blink_counter_cry_13),
            .carryout(blink_counter_cry_14),
            .clk(N__19595),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_15_LC_6_22_7.C_ON=1'b1;
    defparam blink_counter_15_LC_6_22_7.SEQ_MODE=4'b1000;
    defparam blink_counter_15_LC_6_22_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_15_LC_6_22_7 (
            .in0(_gnd_net_),
            .in1(N__8140),
            .in2(_gnd_net_),
            .in3(N__8134),
            .lcout(blink_counterZ0Z_15),
            .ltout(),
            .carryin(blink_counter_cry_14),
            .carryout(blink_counter_cry_15),
            .clk(N__19595),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_16_LC_6_23_0.C_ON=1'b1;
    defparam blink_counter_16_LC_6_23_0.SEQ_MODE=4'b1000;
    defparam blink_counter_16_LC_6_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_16_LC_6_23_0 (
            .in0(_gnd_net_),
            .in1(N__8131),
            .in2(_gnd_net_),
            .in3(N__8125),
            .lcout(blink_counterZ0Z_16),
            .ltout(),
            .carryin(bfn_6_23_0_),
            .carryout(blink_counter_cry_16),
            .clk(N__19600),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_17_LC_6_23_1.C_ON=1'b1;
    defparam blink_counter_17_LC_6_23_1.SEQ_MODE=4'b1000;
    defparam blink_counter_17_LC_6_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_17_LC_6_23_1 (
            .in0(_gnd_net_),
            .in1(N__8122),
            .in2(_gnd_net_),
            .in3(N__8116),
            .lcout(blink_counterZ0Z_17),
            .ltout(),
            .carryin(blink_counter_cry_16),
            .carryout(blink_counter_cry_17),
            .clk(N__19600),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_18_LC_6_23_2.C_ON=1'b1;
    defparam blink_counter_18_LC_6_23_2.SEQ_MODE=4'b1000;
    defparam blink_counter_18_LC_6_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_18_LC_6_23_2 (
            .in0(_gnd_net_),
            .in1(N__8113),
            .in2(_gnd_net_),
            .in3(N__8107),
            .lcout(blink_counterZ0Z_18),
            .ltout(),
            .carryin(blink_counter_cry_17),
            .carryout(blink_counter_cry_18),
            .clk(N__19600),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_19_LC_6_23_3.C_ON=1'b1;
    defparam blink_counter_19_LC_6_23_3.SEQ_MODE=4'b1000;
    defparam blink_counter_19_LC_6_23_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_19_LC_6_23_3 (
            .in0(_gnd_net_),
            .in1(N__8104),
            .in2(_gnd_net_),
            .in3(N__8098),
            .lcout(blink_counterZ0Z_19),
            .ltout(),
            .carryin(blink_counter_cry_18),
            .carryout(blink_counter_cry_19),
            .clk(N__19600),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_20_LC_6_23_4.C_ON=1'b1;
    defparam blink_counter_20_LC_6_23_4.SEQ_MODE=4'b1000;
    defparam blink_counter_20_LC_6_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_20_LC_6_23_4 (
            .in0(_gnd_net_),
            .in1(N__8095),
            .in2(_gnd_net_),
            .in3(N__8089),
            .lcout(blink_counterZ0Z_20),
            .ltout(),
            .carryin(blink_counter_cry_19),
            .carryout(blink_counter_cry_20),
            .clk(N__19600),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_21_LC_6_23_5.C_ON=1'b1;
    defparam blink_counter_21_LC_6_23_5.SEQ_MODE=4'b1000;
    defparam blink_counter_21_LC_6_23_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_21_LC_6_23_5 (
            .in0(_gnd_net_),
            .in1(N__9294),
            .in2(_gnd_net_),
            .in3(N__8185),
            .lcout(blink_counterZ0Z_21),
            .ltout(),
            .carryin(blink_counter_cry_20),
            .carryout(blink_counter_cry_21),
            .clk(N__19600),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_22_LC_6_23_6.C_ON=1'b1;
    defparam blink_counter_22_LC_6_23_6.SEQ_MODE=4'b1000;
    defparam blink_counter_22_LC_6_23_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_22_LC_6_23_6 (
            .in0(_gnd_net_),
            .in1(N__9273),
            .in2(_gnd_net_),
            .in3(N__8182),
            .lcout(blink_counterZ0Z_22),
            .ltout(),
            .carryin(blink_counter_cry_21),
            .carryout(blink_counter_cry_22),
            .clk(N__19600),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_23_LC_6_23_7.C_ON=1'b1;
    defparam blink_counter_23_LC_6_23_7.SEQ_MODE=4'b1000;
    defparam blink_counter_23_LC_6_23_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_23_LC_6_23_7 (
            .in0(_gnd_net_),
            .in1(N__9201),
            .in2(_gnd_net_),
            .in3(N__8179),
            .lcout(blink_counterZ0Z_23),
            .ltout(),
            .carryin(blink_counter_cry_22),
            .carryout(blink_counter_cry_23),
            .clk(N__19600),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_24_LC_6_24_0.C_ON=1'b1;
    defparam blink_counter_24_LC_6_24_0.SEQ_MODE=4'b1000;
    defparam blink_counter_24_LC_6_24_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_24_LC_6_24_0 (
            .in0(_gnd_net_),
            .in1(N__9249),
            .in2(_gnd_net_),
            .in3(N__8176),
            .lcout(blink_counterZ0Z_24),
            .ltout(),
            .carryin(bfn_6_24_0_),
            .carryout(blink_counter_cry_24),
            .clk(N__19607),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_25_LC_6_24_1.C_ON=1'b0;
    defparam blink_counter_25_LC_6_24_1.SEQ_MODE=4'b1000;
    defparam blink_counter_25_LC_6_24_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 blink_counter_25_LC_6_24_1 (
            .in0(_gnd_net_),
            .in1(N__9222),
            .in2(_gnd_net_),
            .in3(N__8173),
            .lcout(blink_counterZ0Z_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19607),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_2_LC_7_17_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_2_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_2_LC_7_17_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_2_LC_7_17_1  (
            .in0(N__14104),
            .in1(_gnd_net_),
            .in2(N__14237),
            .in3(N__14176),
            .lcout(),
            .ltout(\c0.rx.r_Rx_Bytece_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_2_LC_7_17_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_2_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_2_LC_7_17_2 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \c0.rx.r_Rx_Byte_2_LC_7_17_2  (
            .in0(N__12210),
            .in1(N__9047),
            .in2(N__8170),
            .in3(N__8232),
            .lcout(\c0.rx_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_RNIHTCD_1_LC_7_17_4 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_RNIHTCD_1_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Bit_Index_RNIHTCD_1_LC_7_17_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \c0.rx.r_Bit_Index_RNIHTCD_1_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__14217),
            .in2(_gnd_net_),
            .in3(N__14103),
            .lcout(\c0.rx.N_325 ),
            .ltout(\c0.rx.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_2_LC_7_17_5 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_2_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_2_LC_7_17_5 .LUT_INIT=16'b1010011000000000;
    LogicCell40 \c0.rx.r_Bit_Index_2_LC_7_17_5  (
            .in0(N__14180),
            .in1(N__8257),
            .in2(N__8161),
            .in3(N__8850),
            .lcout(\c0.rx.r_Bit_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_5_LC_7_17_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_5_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_5_LC_7_17_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_5_LC_7_17_6  (
            .in0(N__14177),
            .in1(N__14221),
            .in2(_gnd_net_),
            .in3(N__14105),
            .lcout(),
            .ltout(\c0.rx.r_Rx_Bytece_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_5_LC_7_17_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_5_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_5_LC_7_17_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \c0.rx.r_Rx_Byte_5_LC_7_17_7  (
            .in0(N__8233),
            .in1(N__15717),
            .in2(N__8260),
            .in3(N__9049),
            .lcout(\c0.rx_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNI91B33_0_LC_7_18_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNI91B33_0_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNI91B33_0_LC_7_18_0 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \c0.rx.r_SM_Main_RNI91B33_0_LC_7_18_0  (
            .in0(N__8710),
            .in1(N__8649),
            .in2(N__8530),
            .in3(N__9103),
            .lcout(\c0.rx.N_388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_0_LC_7_18_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_0_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_0_LC_7_18_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_0_LC_7_18_1  (
            .in0(N__14244),
            .in1(N__14110),
            .in2(_gnd_net_),
            .in3(N__14175),
            .lcout(\c0.rx.r_Rx_Bytece_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_7_LC_7_18_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_7_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_7_LC_7_18_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_7_LC_7_18_3  (
            .in0(N__9052),
            .in1(N__14056),
            .in2(N__10866),
            .in3(N__8231),
            .lcout(\c0.rx_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19584),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_6_LC_7_18_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_6_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_6_LC_7_18_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_6_LC_7_18_4  (
            .in0(N__14111),
            .in1(N__14245),
            .in2(_gnd_net_),
            .in3(N__14179),
            .lcout(),
            .ltout(\c0.rx.r_Rx_Bytece_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_6_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_6_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_6_LC_7_18_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \c0.rx.r_Rx_Byte_6_LC_7_18_5  (
            .in0(N__16068),
            .in1(N__9051),
            .in2(N__8239),
            .in3(N__8230),
            .lcout(\c0.rx_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19584),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNIJ0FM2_2_LC_7_18_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNIJ0FM2_2_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNIJ0FM2_2_LC_7_18_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.rx.r_SM_Main_RNIJ0FM2_2_LC_7_18_6  (
            .in0(N__8709),
            .in1(N__9102),
            .in2(_gnd_net_),
            .in3(N__8648),
            .lcout(\c0.rx.r_Rx_Byte_1_sqmuxa ),
            .ltout(\c0.rx.r_Rx_Byte_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_0_LC_7_18_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_0_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_0_LC_7_18_7 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.rx.r_Rx_Byte_0_LC_7_18_7  (
            .in0(N__10413),
            .in1(N__8200),
            .in2(N__8194),
            .in3(N__9050),
            .lcout(\c0.rx_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19584),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_0_LC_7_19_0 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count_RNO_0_0_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_0_LC_7_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_0_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__8272),
            .in2(N__8467),
            .in3(N__8466),
            .lcout(\c0.rx.r_Clock_Count_RNO_0_0_0 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\c0.rx.un1_r_Clock_Count_5_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_1_LC_7_19_1 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count_RNO_0_1_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_1_LC_7_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_1_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__8284),
            .in2(_gnd_net_),
            .in3(N__8323),
            .lcout(\c0.rx.r_Clock_Count_RNO_0_0_1 ),
            .ltout(),
            .carryin(\c0.rx.un1_r_Clock_Count_5_cry_0 ),
            .carryout(\c0.rx.un1_r_Clock_Count_5_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_2_LC_7_19_2 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count_RNO_0_2_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_2_LC_7_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_2_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__8434),
            .in2(_gnd_net_),
            .in3(N__8320),
            .lcout(\c0.rx.r_Clock_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\c0.rx.un1_r_Clock_Count_5_cry_1 ),
            .carryout(\c0.rx.un1_r_Clock_Count_5_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_3_LC_7_19_3 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count_RNO_0_3_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_3_LC_7_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_3_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__8737),
            .in2(_gnd_net_),
            .in3(N__8317),
            .lcout(\c0.rx.r_Clock_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\c0.rx.un1_r_Clock_Count_5_cry_2 ),
            .carryout(\c0.rx.un1_r_Clock_Count_5_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_4_LC_7_19_4 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count_RNO_0_4_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_4_LC_7_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_4_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__8395),
            .in2(_gnd_net_),
            .in3(N__8308),
            .lcout(\c0.rx.r_Clock_Count_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\c0.rx.un1_r_Clock_Count_5_cry_3 ),
            .carryout(\c0.rx.un1_r_Clock_Count_5_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_5_LC_7_19_5 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count_RNO_0_5_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_5_LC_7_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_5_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__8377),
            .in2(_gnd_net_),
            .in3(N__8305),
            .lcout(\c0.rx.r_Clock_Count_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\c0.rx.un1_r_Clock_Count_5_cry_4 ),
            .carryout(\c0.rx.un1_r_Clock_Count_5_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_6_LC_7_19_6 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count_RNO_0_6_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_6_LC_7_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_6_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__8422),
            .in2(_gnd_net_),
            .in3(N__8296),
            .lcout(\c0.rx.r_Clock_Count_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\c0.rx.un1_r_Clock_Count_5_cry_5 ),
            .carryout(\c0.rx.un1_r_Clock_Count_5_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_7_LC_7_19_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_0_7_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_7_LC_7_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_7_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__8409),
            .in2(_gnd_net_),
            .in3(N__8293),
            .lcout(\c0.rx.r_Clock_Count_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNIL4RQ_0_LC_7_20_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNIL4RQ_0_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNIL4RQ_0_LC_7_20_0 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNIL4RQ_0_LC_7_20_0  (
            .in0(N__8433),
            .in1(N__8283),
            .in2(_gnd_net_),
            .in3(N__8271),
            .lcout(\c0.rx.N_320 ),
            .ltout(\c0.rx.N_320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNITSB13_3_LC_7_20_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNITSB13_3_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNITSB13_3_LC_7_20_1 .LUT_INIT=16'b0011001111110110;
    LogicCell40 \c0.rx.r_Clock_Count_RNITSB13_3_LC_7_20_1  (
            .in0(N__8734),
            .in1(N__8943),
            .in2(N__8473),
            .in3(N__8351),
            .lcout(\c0.rx.r_Clock_Count_8_f0_0_o2_0_2 ),
            .ltout(\c0.rx.r_Clock_Count_8_f0_0_o2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNINFV94_0_4_LC_7_20_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNINFV94_0_4_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNINFV94_0_4_LC_7_20_2 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \c0.rx.r_SM_Main_RNINFV94_0_4_LC_7_20_2  (
            .in0(N__8944),
            .in1(N__8579),
            .in2(N__8470),
            .in3(N__8625),
            .lcout(\c0.rx.un1_r_Clock_Count_2_sqmuxa_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNICMJ72_3_LC_7_20_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNICMJ72_3_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNICMJ72_3_LC_7_20_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \c0.rx.r_Clock_Count_RNICMJ72_3_LC_7_20_3  (
            .in0(N__8735),
            .in1(N__8364),
            .in2(_gnd_net_),
            .in3(N__8352),
            .lcout(\c0.rx.N_386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNINFV94_4_LC_7_20_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNINFV94_4_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNINFV94_4_LC_7_20_4 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \c0.rx.r_SM_Main_RNINFV94_4_LC_7_20_4  (
            .in0(N__8945),
            .in1(N__8580),
            .in2(N__8452),
            .in3(N__8626),
            .lcout(\c0.rx.N_332 ),
            .ltout(\c0.rx.N_332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_2_LC_7_20_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_2_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_2_LC_7_20_5 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \c0.rx.r_Clock_Count_2_LC_7_20_5  (
            .in0(N__8443),
            .in1(N__8912),
            .in2(N__8437),
            .in3(N__8833),
            .lcout(\c0.rx.r_Clock_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19589),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_7_20_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_7_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_7_20_6  (
            .in0(N__8421),
            .in1(N__8376),
            .in2(N__8410),
            .in3(N__8394),
            .lcout(\c0.rx.N_317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_5_LC_7_20_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_5_LC_7_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_5_LC_7_20_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.rx.r_Clock_Count_5_LC_7_20_7  (
            .in0(N__8383),
            .in1(N__8881),
            .in2(N__8786),
            .in3(N__8834),
            .lcout(\c0.rx.r_Clock_CountZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19589),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNICMJ72_0_3_LC_7_21_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNICMJ72_0_3_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNICMJ72_0_3_LC_7_21_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.rx.r_Clock_Count_RNICMJ72_0_3_LC_7_21_0  (
            .in0(N__8365),
            .in1(N__8736),
            .in2(_gnd_net_),
            .in3(N__8353),
            .lcout(\c0.rx.N_383 ),
            .ltout(\c0.rx.N_383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_1_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_1_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_1_LC_7_21_1 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.rx.r_SM_Main_1_LC_7_21_1  (
            .in0(N__8644),
            .in1(N__8338),
            .in2(N__8332),
            .in3(N__8524),
            .lcout(\c0.rx.r_SM_Main_dup_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19596),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.N_98_ip_RNO_1_LC_7_21_2 .C_ON=1'b0;
    defparam \c0.rx.N_98_ip_RNO_1_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.N_98_ip_RNO_1_LC_7_21_2 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \c0.rx.N_98_ip_RNO_1_LC_7_21_2  (
            .in0(N__9140),
            .in1(N__8512),
            .in2(_gnd_net_),
            .in3(N__9093),
            .lcout(\c0.rx.r_SM_Main_illegal_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNO_0_0_LC_7_21_3 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNO_0_0_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNO_0_0_LC_7_21_3 .LUT_INIT=16'b0000010100001111;
    LogicCell40 \c0.rx.r_SM_Main_RNO_0_0_LC_7_21_3  (
            .in0(N__8969),
            .in1(_gnd_net_),
            .in2(N__8526),
            .in3(N__9142),
            .lcout(),
            .ltout(\c0.rx.N_138r_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_0_LC_7_21_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_0_LC_7_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_0_LC_7_21_4 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \c0.rx.r_SM_Main_0_LC_7_21_4  (
            .in0(N__9061),
            .in1(N__8570),
            .in2(N__8533),
            .in3(N__8645),
            .lcout(\c0.rx.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19596),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.N_98_ip_RNO_0_LC_7_21_5 .C_ON=1'b0;
    defparam \c0.rx.N_98_ip_RNO_0_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.N_98_ip_RNO_0_LC_7_21_5 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \c0.rx.N_98_ip_RNO_0_LC_7_21_5  (
            .in0(N__9091),
            .in1(_gnd_net_),
            .in2(N__8525),
            .in3(N__9141),
            .lcout(),
            .ltout(\c0.rx.N_91_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.N_98_ip_LC_7_21_6 .C_ON=1'b0;
    defparam \c0.rx.N_98_ip_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.N_98_ip_LC_7_21_6 .LUT_INIT=16'b1001111011111111;
    LogicCell40 \c0.rx.N_98_ip_LC_7_21_6  (
            .in0(N__8673),
            .in1(N__8569),
            .in2(N__8485),
            .in3(N__8482),
            .lcout(\c0.rx.N_98_dup ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNIH6OP_3_LC_7_21_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNIH6OP_3_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNIH6OP_3_LC_7_21_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.r_SM_Main_RNIH6OP_3_LC_7_21_7  (
            .in0(N__9092),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8672),
            .lcout(\c0.rx.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2_LC_7_22_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2_LC_7_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_2_LC_7_22_0 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \c0.rx.r_SM_Main_2_LC_7_22_0  (
            .in0(N__9067),
            .in1(N__8970),
            .in2(N__9154),
            .in3(N__8634),
            .lcout(\c0.rx.r_SM_Main_dup_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNO_0_3_LC_7_22_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNO_0_3_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNO_0_3_LC_7_22_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.r_SM_Main_RNO_0_3_LC_7_22_1  (
            .in0(N__14184),
            .in1(N__14125),
            .in2(N__14251),
            .in3(N__9096),
            .lcout(),
            .ltout(\c0.rx.r_SM_Main_ns_0_i_a2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_3_LC_7_22_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_3_LC_7_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_3_LC_7_22_2 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \c0.rx.r_SM_Main_3_LC_7_22_2  (
            .in0(N__8676),
            .in1(N__8707),
            .in2(N__8476),
            .in3(N__8635),
            .lcout(\c0.rx.r_SM_Main_dup_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNO_1_2_LC_7_22_3 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNO_1_2_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNO_1_2_LC_7_22_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.rx.r_SM_Main_RNO_1_2_LC_7_22_3  (
            .in0(N__9144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9060),
            .lcout(\c0.rx.r_SM_Main_ns_0_i_a2_1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNIHKFL1_1_LC_7_22_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNIHKFL1_1_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNIHKFL1_1_LC_7_22_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \c0.rx.r_SM_Main_RNIHKFL1_1_LC_7_22_4  (
            .in0(N__8946),
            .in1(N__9143),
            .in2(N__8650),
            .in3(N__8567),
            .lcout(\c0.rx.N_361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_RNO_1_LC_7_22_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_RNO_1_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_DV_RNO_1_LC_7_22_5 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \c0.rx.r_Rx_DV_RNO_1_LC_7_22_5  (
            .in0(N__8566),
            .in1(N__8674),
            .in2(_gnd_net_),
            .in3(N__9094),
            .lcout(),
            .ltout(\c0.rx.un1_r_Rx_DV7_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_RNO_0_LC_7_22_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_RNO_0_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_DV_RNO_0_LC_7_22_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \c0.rx.r_Rx_DV_RNO_0_LC_7_22_6  (
            .in0(N__8675),
            .in1(N__8705),
            .in2(N__9118),
            .in3(N__8633),
            .lcout(\c0.rx.r_Rx_DV_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNO_0_2_LC_7_22_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNO_0_2_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNO_0_2_LC_7_22_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \c0.rx.r_SM_Main_RNO_0_2_LC_7_22_7  (
            .in0(N__8706),
            .in1(N__14049),
            .in2(_gnd_net_),
            .in3(N__9095),
            .lcout(\c0.rx.r_SM_Main_ns_0_i_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNI7GPF_4_LC_7_23_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNI7GPF_4_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNI7GPF_4_LC_7_23_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.rx.r_SM_Main_RNI7GPF_4_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__9053),
            .in2(_gnd_net_),
            .in3(N__8568),
            .lcout(),
            .ltout(\c0.rx.r_Clock_Count_8_f0_0_a2_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.N_98_ip_RNIJK4J3_LC_7_23_1 .C_ON=1'b0;
    defparam \c0.rx.N_98_ip_RNIJK4J3_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.N_98_ip_RNIJK4J3_LC_7_23_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \c0.rx.N_98_ip_RNIJK4J3_LC_7_23_1  (
            .in0(N__8971),
            .in1(N__8950),
            .in2(N__8923),
            .in3(N__8646),
            .lcout(\c0.rx.N_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_3_LC_7_23_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_3_LC_7_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_3_LC_7_23_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.rx.r_Clock_Count_3_LC_7_23_3  (
            .in0(N__8890),
            .in1(N__8854),
            .in2(N__8775),
            .in3(N__8746),
            .lcout(\c0.rx.r_Clock_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19608),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_4_LC_7_23_5 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_4_LC_7_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_4_LC_7_23_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.rx.r_SM_Main_4_LC_7_23_5  (
            .in0(N__8708),
            .in1(N__8677),
            .in2(_gnd_net_),
            .in3(N__8647),
            .lcout(\c0.rx.r_SM_Main_dup_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19608),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__3_LC_7_25_5 .C_ON=1'b0;
    defparam \c0.data_out_2__3_LC_7_25_5 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__3_LC_7_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__3_LC_7_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17075),
            .lcout(\c0.d_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19621),
            .ce(),
            .sr(N__16881));
    defparam \c0.data_out_0__5_LC_7_25_6 .C_ON=1'b0;
    defparam \c0.data_out_0__5_LC_7_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__5_LC_7_25_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_0__5_LC_7_25_6  (
            .in0(N__17074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19621),
            .ce(),
            .sr(N__16881));
    defparam \c0.data_out_1__1_LC_7_26_7 .C_ON=1'b0;
    defparam \c0.data_out_1__1_LC_7_26_7 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__1_LC_7_26_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_1__1_LC_7_26_7  (
            .in0(N__17060),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19631),
            .ce(),
            .sr(N__16880));
    defparam \c0.data_out_7__7_LC_9_16_7 .C_ON=1'b0;
    defparam \c0.data_out_7__7_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__7_LC_9_16_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_7__7_LC_9_16_7  (
            .in0(N__14875),
            .in1(N__14503),
            .in2(N__9385),
            .in3(N__10090),
            .lcout(\c0.data_out_7_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19590),
            .ce(N__16838),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_7_c_RNO_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNO_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNO_LC_9_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_RNO_LC_9_18_0  (
            .in0(N__11336),
            .in1(N__11048),
            .in2(N__13965),
            .in3(N__12347),
            .lcout(\c0.i12_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__5_LC_9_18_2 .C_ON=1'b0;
    defparam \c0.data_in_3__5_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__5_LC_9_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__5_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11170),
            .lcout(\c0.data_in_3_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19591),
            .ce(N__17716),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__6_LC_9_18_3 .C_ON=1'b0;
    defparam \c0.data_in_3__6_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__6_LC_9_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__6_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16102),
            .lcout(\c0.data_in_3_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19591),
            .ce(N__17716),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__6_LC_9_18_5 .C_ON=1'b0;
    defparam \c0.data_in_2__6_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__6_LC_9_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__6_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11337),
            .lcout(\c0.data_in_2_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19591),
            .ce(N__17716),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__6_LC_9_18_6 .C_ON=1'b0;
    defparam \c0.data_in_1__6_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__6_LC_9_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__6_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13613),
            .lcout(\c0.data_in_1_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19591),
            .ce(N__17716),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_0_c_LC_9_19_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_0_c_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_0_c_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_0_c_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__9160),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\c0.i12_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_1_c_LC_9_19_1 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_1_c_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_1_c_LC_9_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_1_c_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__9307),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_0 ),
            .carryout(\c0.i12_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_2_c_LC_9_19_2 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_2_c_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_2_c_LC_9_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_2_c_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__9676),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_1 ),
            .carryout(\c0.i12_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_3_c_LC_9_19_3 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_3_c_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_3_c_LC_9_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_3_c_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__9640),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_2 ),
            .carryout(\c0.i12_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_4_c_LC_9_19_4 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_4_c_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_4_c_LC_9_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_4_c_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__9721),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_3 ),
            .carryout(\c0.i12_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_5_c_LC_9_19_5 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_5_c_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_5_c_LC_9_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_5_c_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__9688),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_4 ),
            .carryout(\c0.i12_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_6_c_LC_9_19_6 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_6_c_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_6_c_LC_9_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_6_c_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__9682),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_5 ),
            .carryout(\c0.i12_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_7_c_LC_9_19_7 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_7_c_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_LC_9_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9172),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_6 ),
            .carryout(\c0.i12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_THRU_LUT4_0_LC_9_20_0 .C_ON=1'b0;
    defparam \c0.i12_THRU_LUT4_0_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_THRU_LUT4_0_LC_9_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.i12_THRU_LUT4_0_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9163),
            .lcout(\c0.i12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_0_c_RNO_LC_9_20_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_0_c_RNO_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_0_c_RNO_LC_9_20_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_0_c_RNO_LC_9_20_1  (
            .in0(N__10254),
            .in1(N__12711),
            .in2(N__13506),
            .in3(N__16113),
            .lcout(\c0.i12_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_1_c_RNO_LC_9_20_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_1_c_RNO_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_1_c_RNO_LC_9_20_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_1_c_RNO_LC_9_20_3  (
            .in0(N__15869),
            .in1(N__10241),
            .in2(N__11127),
            .in3(N__10968),
            .lcout(\c0.i12_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED_obuf_RNO_1_LC_9_21_1.C_ON=1'b0;
    defparam LED_obuf_RNO_1_LC_9_21_1.SEQ_MODE=4'b0000;
    defparam LED_obuf_RNO_1_LC_9_21_1.LUT_INIT=16'b1010100010001010;
    LogicCell40 LED_obuf_RNO_1_LC_9_21_1 (
            .in0(N__9301),
            .in1(N__9283),
            .in2(N__9262),
            .in3(N__9231),
            .lcout(N_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED_obuf_RNO_0_LC_9_21_2.C_ON=1'b0;
    defparam LED_obuf_RNO_0_LC_9_21_2.SEQ_MODE=4'b0000;
    defparam LED_obuf_RNO_0_LC_9_21_2.LUT_INIT=16'b0010001000100010;
    LogicCell40 LED_obuf_RNO_0_LC_9_21_2 (
            .in0(N__9282),
            .in1(N__9258),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(N_8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED_obuf_RNO_LC_9_21_3.C_ON=1'b0;
    defparam LED_obuf_RNO_LC_9_21_3.SEQ_MODE=4'b0000;
    defparam LED_obuf_RNO_LC_9_21_3.LUT_INIT=16'b0100000101010101;
    LogicCell40 LED_obuf_RNO_LC_9_21_3 (
            .in0(N__9238),
            .in1(N__9232),
            .in2(N__9211),
            .in3(N__9208),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__1_LC_9_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0__1_LC_9_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__1_LC_9_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__1_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15870),
            .lcout(\c0.data_in_0_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19609),
            .ce(N__17723),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__3_LC_9_21_5 .C_ON=1'b0;
    defparam \c0.data_in_0__3_LC_9_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__3_LC_9_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__3_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11123),
            .lcout(\c0.data_in_0_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19609),
            .ce(N__17723),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__4_LC_9_21_6 .C_ON=1'b0;
    defparam \c0.data_in_0__4_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__4_LC_9_21_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_0__4_LC_9_21_6  (
            .in0(N__13773),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_0_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19609),
            .ce(N__17723),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__6_LC_9_21_7 .C_ON=1'b0;
    defparam \c0.data_in_0__6_LC_9_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__6_LC_9_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__6_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13716),
            .lcout(\c0.data_in_0_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19609),
            .ce(N__17723),
            .sr(_gnd_net_));
    defparam \c0.tx.N_90_ip_RNO_1_LC_9_22_0 .C_ON=1'b0;
    defparam \c0.tx.N_90_ip_RNO_1_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.N_90_ip_RNO_1_LC_9_22_0 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \c0.tx.N_90_ip_RNO_1_LC_9_22_0  (
            .in0(N__10650),
            .in1(N__10529),
            .in2(_gnd_net_),
            .in3(N__9852),
            .lcout(\c0.tx.r_SM_Main_illegal_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.N_90_ip_RNIVJLQ_LC_9_22_1 .C_ON=1'b0;
    defparam \c0.tx.N_90_ip_RNIVJLQ_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.N_90_ip_RNIVJLQ_LC_9_22_1 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.tx.N_90_ip_RNIVJLQ_LC_9_22_1  (
            .in0(N__9855),
            .in1(N__9940),
            .in2(_gnd_net_),
            .in3(N__9817),
            .lcout(\c0.tx.N_90_ip_RNIVJLQZ0 ),
            .ltout(\c0.tx.N_90_ip_RNIVJLQZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.N_90_ip_RNIVJLQ_0_LC_9_22_2 .C_ON=1'b0;
    defparam \c0.tx.N_90_ip_RNIVJLQ_0_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.N_90_ip_RNIVJLQ_0_LC_9_22_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \c0.tx.N_90_ip_RNIVJLQ_0_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9370),
            .in3(_gnd_net_),
            .lcout(\c0.tx.N_398_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.N_90_ip_LC_9_22_3 .C_ON=1'b0;
    defparam \c0.tx.N_90_ip_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.N_90_ip_LC_9_22_3 .LUT_INIT=16'b1011011111111011;
    LogicCell40 \c0.tx.N_90_ip_LC_9_22_3  (
            .in0(N__10316),
            .in1(N__9367),
            .in2(N__9984),
            .in3(N__9358),
            .lcout(\c0.tx.N_90_dup ),
            .ltout(\c0.tx.N_90_dup_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNI1GI71_4_LC_9_22_4 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNI1GI71_4_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNI1GI71_4_LC_9_22_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.tx.r_SM_Main_RNI1GI71_4_LC_9_22_4  (
            .in0(N__9980),
            .in1(N__9854),
            .in2(N__9361),
            .in3(N__9770),
            .lcout(\c0.tx.r_Clock_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_3_LC_9_22_5 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_3_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_3_LC_9_22_5 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.tx.r_SM_Main_3_LC_9_22_5  (
            .in0(N__10317),
            .in1(N__9904),
            .in2(N__10618),
            .in3(N__9818),
            .lcout(\c0.tx.r_SM_Main_dup_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19616),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.N_90_ip_RNO_0_LC_9_22_6 .C_ON=1'b0;
    defparam \c0.tx.N_90_ip_RNO_0_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.N_90_ip_RNO_0_LC_9_22_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.tx.N_90_ip_RNO_0_LC_9_22_6  (
            .in0(N__10651),
            .in1(N__10530),
            .in2(_gnd_net_),
            .in3(N__9853),
            .lcout(\c0.tx.N_83_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_0_LC_9_22_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_0_LC_9_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_0_LC_9_22_7 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \c0.tx.r_SM_Main_0_LC_9_22_7  (
            .in0(N__9979),
            .in1(N__9819),
            .in2(N__9913),
            .in3(N__10652),
            .lcout(\c0.tx.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19616),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNO_0_0_LC_9_23_0 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count_RNO_0_0_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNO_0_0_LC_9_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx.r_Clock_Count_RNO_0_0_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__9427),
            .in2(N__9351),
            .in3(N__9352),
            .lcout(\c0.tx.r_Clock_Count_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\c0.tx.un1_r_Clock_Count_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNO_0_1_LC_9_23_1 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count_RNO_0_1_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNO_0_1_LC_9_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx.r_Clock_Count_RNO_0_1_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__9471),
            .in2(_gnd_net_),
            .in3(N__9310),
            .lcout(\c0.tx.r_Clock_Count_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\c0.tx.un1_r_Clock_Count_cry_0 ),
            .carryout(\c0.tx.un1_r_Clock_Count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNO_0_2_LC_9_23_2 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count_RNO_0_2_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNO_0_2_LC_9_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx.r_Clock_Count_RNO_0_2_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__9493),
            .in2(_gnd_net_),
            .in3(N__9508),
            .lcout(\c0.tx.r_Clock_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\c0.tx.un1_r_Clock_Count_cry_1 ),
            .carryout(\c0.tx.un1_r_Clock_Count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNO_0_3_LC_9_23_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_RNO_0_3_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNO_0_3_LC_9_23_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.tx.r_Clock_Count_RNO_0_3_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__9450),
            .in2(_gnd_net_),
            .in3(N__9505),
            .lcout(\c0.tx.r_Clock_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNI522E_4_LC_9_23_4 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNI522E_4_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNI522E_4_LC_9_23_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.r_SM_Main_RNI522E_4_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__9985),
            .in2(_gnd_net_),
            .in3(N__9820),
            .lcout(\c0.tx.r_SM_Main_RNI522EZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNI636A_3_LC_9_23_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_RNI636A_3_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNI636A_3_LC_9_23_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.r_Clock_Count_RNI636A_3_LC_9_23_6  (
            .in0(N__9492),
            .in1(N__9472),
            .in2(N__9451),
            .in3(N__9426),
            .lcout(\c0.tx.N_171_0 ),
            .ltout(\c0.tx.N_171_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_1_LC_9_23_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_1_LC_9_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_1_LC_9_23_7 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.tx.r_SM_Main_1_LC_9_23_7  (
            .in0(N__9821),
            .in1(N__9409),
            .in2(N__9397),
            .in3(N__9863),
            .lcout(\c0.tx.r_SM_Main_dup_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_0_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_0_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_0_LC_9_24_0 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_1_0_LC_9_24_0  (
            .in0(N__9391),
            .in1(N__15529),
            .in2(N__10063),
            .in3(N__15379),
            .lcout(\c0.tx_data_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_0_LC_9_24_1 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_0_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_0_LC_9_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__RNO_0_0_LC_9_24_1  (
            .in0(N__13013),
            .in1(N__14470),
            .in2(_gnd_net_),
            .in3(N__11778),
            .lcout(),
            .ltout(\c0.nextCRC16_3_0_a2_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__0_LC_9_24_2 .C_ON=1'b0;
    defparam \c0.data_out_6__0_LC_9_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__0_LC_9_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__0_LC_9_24_2  (
            .in0(N__14498),
            .in1(N__11517),
            .in2(N__9394),
            .in3(N__10023),
            .lcout(\c0.data_out_6_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19632),
            .ce(N__16837),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_7_LC_9_24_6 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_7_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_7_LC_9_24_6 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.data_out_7__RNO_0_7_LC_9_24_6  (
            .in0(N__10896),
            .in1(N__13329),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__5_LC_9_25_0 .C_ON=1'b0;
    defparam \c0.data_out_5__5_LC_9_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__5_LC_9_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__5_LC_9_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9610),
            .lcout(\c0.d_2_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19638),
            .ce(N__16836),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__1_LC_9_25_2 .C_ON=1'b0;
    defparam \c0.data_out_4__1_LC_9_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__1_LC_9_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__1_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9571),
            .lcout(\c0.d_2_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19638),
            .ce(N__16836),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__3_LC_9_25_6 .C_ON=1'b0;
    defparam \c0.data_out_5__3_LC_9_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__3_LC_9_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__3_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9631),
            .lcout(\c0.d_2_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19638),
            .ce(N__16836),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__1_LC_9_26_3 .C_ON=1'b0;
    defparam \c0.data_out_5__1_LC_9_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__1_LC_9_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__1_LC_9_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9532),
            .lcout(\c0.d_2_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19646),
            .ce(N__16834),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__7_LC_9_26_4 .C_ON=1'b0;
    defparam \c0.data_out_5__7_LC_9_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__7_LC_9_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__7_LC_9_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9589),
            .lcout(\c0.d_2_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19646),
            .ce(N__16834),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__5_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.data_out_4__5_LC_9_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__5_LC_9_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__5_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9664),
            .lcout(\c0.d_2_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19646),
            .ce(N__16834),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__2_LC_9_26_7 .C_ON=1'b0;
    defparam \c0.data_out_4__2_LC_9_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__2_LC_9_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__2_LC_9_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9553),
            .lcout(\c0.d_2_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19646),
            .ce(N__16834),
            .sr(_gnd_net_));
    defparam \c0.data_0_LC_9_27_0 .C_ON=1'b1;
    defparam \c0.data_0_LC_9_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_0_LC_9_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_0_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__10185),
            .in2(_gnd_net_),
            .in3(N__9535),
            .lcout(\c0.dataZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\c0.data_cry_0 ),
            .clk(N__19652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_1_LC_9_27_1 .C_ON=1'b1;
    defparam \c0.data_1_LC_9_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_1_LC_9_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_1_LC_9_27_1  (
            .in0(_gnd_net_),
            .in1(N__9531),
            .in2(_gnd_net_),
            .in3(N__9520),
            .lcout(\c0.dataZ0Z_1 ),
            .ltout(),
            .carryin(\c0.data_cry_0 ),
            .carryout(\c0.data_cry_1 ),
            .clk(N__19652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_2_LC_9_27_2 .C_ON=1'b1;
    defparam \c0.data_2_LC_9_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_2_LC_9_27_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_2_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(N__10149),
            .in2(_gnd_net_),
            .in3(N__9634),
            .lcout(\c0.dataZ0Z_2 ),
            .ltout(),
            .carryin(\c0.data_cry_1 ),
            .carryout(\c0.data_cry_2 ),
            .clk(N__19652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_3_LC_9_27_3 .C_ON=1'b1;
    defparam \c0.data_3_LC_9_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_3_LC_9_27_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_3_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__9627),
            .in2(_gnd_net_),
            .in3(N__9616),
            .lcout(\c0.dataZ0Z_3 ),
            .ltout(),
            .carryin(\c0.data_cry_2 ),
            .carryout(\c0.data_cry_3 ),
            .clk(N__19652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_4_LC_9_27_4 .C_ON=1'b1;
    defparam \c0.data_4_LC_9_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_4_LC_9_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_4_LC_9_27_4  (
            .in0(_gnd_net_),
            .in1(N__10125),
            .in2(_gnd_net_),
            .in3(N__9613),
            .lcout(\c0.dataZ0Z_4 ),
            .ltout(),
            .carryin(\c0.data_cry_3 ),
            .carryout(\c0.data_cry_4 ),
            .clk(N__19652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_5_LC_9_27_5 .C_ON=1'b1;
    defparam \c0.data_5_LC_9_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_5_LC_9_27_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_5_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(N__9606),
            .in2(_gnd_net_),
            .in3(N__9595),
            .lcout(\c0.dataZ0Z_5 ),
            .ltout(),
            .carryin(\c0.data_cry_4 ),
            .carryout(\c0.data_cry_5 ),
            .clk(N__19652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_6_LC_9_27_6 .C_ON=1'b1;
    defparam \c0.data_6_LC_9_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_6_LC_9_27_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_6_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(N__10740),
            .in2(_gnd_net_),
            .in3(N__9592),
            .lcout(\c0.dataZ0Z_6 ),
            .ltout(),
            .carryin(\c0.data_cry_5 ),
            .carryout(\c0.data_cry_6 ),
            .clk(N__19652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_7_LC_9_27_7 .C_ON=1'b1;
    defparam \c0.data_7_LC_9_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_7_LC_9_27_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_7_LC_9_27_7  (
            .in0(_gnd_net_),
            .in1(N__9588),
            .in2(_gnd_net_),
            .in3(N__9577),
            .lcout(\c0.dataZ0Z_7 ),
            .ltout(),
            .carryin(\c0.data_cry_6 ),
            .carryout(\c0.data_cry_7 ),
            .clk(N__19652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_8_LC_9_28_0 .C_ON=1'b1;
    defparam \c0.data_8_LC_9_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_8_LC_9_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_8_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__10113),
            .in2(_gnd_net_),
            .in3(N__9574),
            .lcout(\c0.dataZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_28_0_),
            .carryout(\c0.data_cry_8 ),
            .clk(N__19661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_9_LC_9_28_1 .C_ON=1'b1;
    defparam \c0.data_9_LC_9_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_9_LC_9_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_9_LC_9_28_1  (
            .in0(_gnd_net_),
            .in1(N__9567),
            .in2(_gnd_net_),
            .in3(N__9556),
            .lcout(\c0.dataZ0Z_9 ),
            .ltout(),
            .carryin(\c0.data_cry_8 ),
            .carryout(\c0.data_cry_9 ),
            .clk(N__19661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_10_LC_9_28_2 .C_ON=1'b1;
    defparam \c0.data_10_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_10_LC_9_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_10_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(N__9549),
            .in2(_gnd_net_),
            .in3(N__9538),
            .lcout(\c0.dataZ0Z_10 ),
            .ltout(),
            .carryin(\c0.data_cry_9 ),
            .carryout(\c0.data_cry_10 ),
            .clk(N__19661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_11_LC_9_28_3 .C_ON=1'b1;
    defparam \c0.data_11_LC_9_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_11_LC_9_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_11_LC_9_28_3  (
            .in0(_gnd_net_),
            .in1(N__10161),
            .in2(_gnd_net_),
            .in3(N__9670),
            .lcout(\c0.dataZ0Z_11 ),
            .ltout(),
            .carryin(\c0.data_cry_10 ),
            .carryout(\c0.data_cry_11 ),
            .clk(N__19661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_12_LC_9_28_4 .C_ON=1'b1;
    defparam \c0.data_12_LC_9_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_12_LC_9_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_12_LC_9_28_4  (
            .in0(_gnd_net_),
            .in1(N__10038),
            .in2(_gnd_net_),
            .in3(N__9667),
            .lcout(\c0.dataZ0Z_12 ),
            .ltout(),
            .carryin(\c0.data_cry_11 ),
            .carryout(\c0.data_cry_12 ),
            .clk(N__19661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_13_LC_9_28_5 .C_ON=1'b1;
    defparam \c0.data_13_LC_9_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_13_LC_9_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_13_LC_9_28_5  (
            .in0(_gnd_net_),
            .in1(N__9660),
            .in2(_gnd_net_),
            .in3(N__9649),
            .lcout(\c0.dataZ0Z_13 ),
            .ltout(),
            .carryin(\c0.data_cry_12 ),
            .carryout(\c0.data_cry_13 ),
            .clk(N__19661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_14_LC_9_28_6 .C_ON=1'b1;
    defparam \c0.data_14_LC_9_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_14_LC_9_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_14_LC_9_28_6  (
            .in0(_gnd_net_),
            .in1(N__10173),
            .in2(_gnd_net_),
            .in3(N__9646),
            .lcout(\c0.dataZ0Z_14 ),
            .ltout(),
            .carryin(\c0.data_cry_13 ),
            .carryout(\c0.data_cry_14 ),
            .clk(N__19661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_15_LC_9_28_7 .C_ON=1'b0;
    defparam \c0.data_15_LC_9_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_15_LC_9_28_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_15_LC_9_28_7  (
            .in0(_gnd_net_),
            .in1(N__10137),
            .in2(_gnd_net_),
            .in3(N__9643),
            .lcout(\c0.dataZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__4_LC_10_17_2 .C_ON=1'b0;
    defparam \c0.data_in_3__4_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__4_LC_10_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__4_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13663),
            .lcout(\c0.data_in_3_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19586),
            .ce(N__17715),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__0_LC_10_17_4 .C_ON=1'b0;
    defparam \c0.data_in_3__0_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__0_LC_10_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__0_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14409),
            .lcout(\c0.data_in_3_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19586),
            .ce(N__17715),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__7_LC_10_17_5 .C_ON=1'b0;
    defparam \c0.data_in_3__7_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__7_LC_10_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__7_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11241),
            .lcout(\c0.data_in_3_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19586),
            .ce(N__17715),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__0_LC_10_17_6 .C_ON=1'b0;
    defparam \c0.data_in_4__0_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__0_LC_10_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__0_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12270),
            .lcout(\c0.data_in_4_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19586),
            .ce(N__17715),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_0  (
            .in0(N__11012),
            .in1(N__10991),
            .in2(N__10956),
            .in3(N__12674),
            .lcout(\c0.i12_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__2_LC_10_18_1 .C_ON=1'b0;
    defparam \c0.data_in_2__2_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__2_LC_10_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__2_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12306),
            .lcout(\c0.data_in_2_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19593),
            .ce(N__17718),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__5_LC_10_18_3 .C_ON=1'b0;
    defparam \c0.data_in_2__5_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__5_LC_10_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__5_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11049),
            .lcout(\c0.data_in_2_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19593),
            .ce(N__17718),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__7_LC_10_18_4 .C_ON=1'b0;
    defparam \c0.data_in_2__7_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__7_LC_10_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__7_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13964),
            .lcout(\c0.data_in_2_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19593),
            .ce(N__17718),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__2_LC_10_18_5 .C_ON=1'b0;
    defparam \c0.data_in_1__2_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__2_LC_10_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_1__2_LC_10_18_5  (
            .in0(N__12675),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_1_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19593),
            .ce(N__17718),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__2_LC_10_18_6 .C_ON=1'b0;
    defparam \c0.data_in_3__2_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__2_LC_10_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__2_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11181),
            .lcout(\c0.data_in_3_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19593),
            .ce(N__17718),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_18_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_18_7  (
            .in0(N__11072),
            .in1(N__12305),
            .in2(N__12388),
            .in3(N__15842),
            .lcout(\c0.i12_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_2_c_RNO_LC_10_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_2_c_RNO_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_2_c_RNO_LC_10_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_2_c_RNO_LC_10_19_0  (
            .in0(N__11099),
            .in1(N__12323),
            .in2(N__12504),
            .in3(N__13766),
            .lcout(\c0.i12_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__4_LC_10_19_1 .C_ON=1'b0;
    defparam \c0.data_in_1__4_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__4_LC_10_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_1__4_LC_10_19_1  (
            .in0(N__11196),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_1_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19598),
            .ce(N__17719),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__5_LC_10_19_2 .C_ON=1'b0;
    defparam \c0.data_in_1__5_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__5_LC_10_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__5_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11013),
            .lcout(\c0.data_in_1_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19598),
            .ce(N__17719),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__7_LC_10_19_3 .C_ON=1'b0;
    defparam \c0.data_in_1__7_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__7_LC_10_19_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_1__7_LC_10_19_3  (
            .in0(N__10952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_1_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19598),
            .ce(N__17719),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__0_LC_10_19_4 .C_ON=1'b0;
    defparam \c0.data_in_2__0_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__0_LC_10_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__0_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11079),
            .lcout(\c0.data_in_2_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19598),
            .ce(N__17719),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__5_LC_10_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0__5_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__5_LC_10_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_0__5_LC_10_19_5  (
            .in0(N__12324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_0_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19598),
            .ce(N__17719),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__4_LC_10_19_6 .C_ON=1'b0;
    defparam \c0.data_in_2__4_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__4_LC_10_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__4_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12357),
            .lcout(\c0.data_in_2_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19598),
            .ce(N__17719),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_5_c_RNO_LC_10_19_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_5_c_RNO_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_5_c_RNO_LC_10_19_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.FRAME_MATCHER_i12_5_c_RNO_LC_10_19_7  (
            .in0(N__11195),
            .in1(N__11360),
            .in2(N__13617),
            .in3(N__13709),
            .lcout(\c0.i12_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__7_LC_10_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0__7_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__7_LC_10_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__7_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11100),
            .lcout(\c0.data_in_0_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19603),
            .ce(N__17721),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__0_LC_10_20_2 .C_ON=1'b0;
    defparam \c0.data_in_1__0_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__0_LC_10_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__0_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12500),
            .lcout(\c0.data_in_1_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19603),
            .ce(N__17721),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__1_LC_10_20_3 .C_ON=1'b0;
    defparam \c0.data_in_1__1_LC_10_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__1_LC_10_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__1_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11361),
            .lcout(\c0.data_in_1_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19603),
            .ce(N__17721),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__3_LC_10_20_4 .C_ON=1'b0;
    defparam \c0.data_in_1__3_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__3_LC_10_20_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_1__3_LC_10_20_4  (
            .in0(N__10996),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_1_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19603),
            .ce(N__17721),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__0_LC_10_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0__0_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__0_LC_10_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__0_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10242),
            .lcout(\c0.data_in_0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19603),
            .ce(N__17721),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_20_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_20_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_20_6  (
            .in0(N__12693),
            .in1(N__14430),
            .in2(N__15933),
            .in3(N__11142),
            .lcout(\c0.i12_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__2_LC_10_20_7 .C_ON=1'b0;
    defparam \c0.data_in_0__2_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__2_LC_10_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__2_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15929),
            .lcout(\c0.data_in_0_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19603),
            .ce(N__17721),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_RNO_0_2_LC_10_21_0 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_RNO_0_2_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_RNO_0_2_LC_10_21_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.tx.r_Bit_Index_RNO_0_2_LC_10_21_0  (
            .in0(N__10486),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9734),
            .lcout(),
            .ltout(\c0.tx.r_Bit_Index_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_2_LC_10_21_1 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_2_LC_10_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_2_LC_10_21_1 .LUT_INIT=16'b1000010010001000;
    LogicCell40 \c0.tx.r_Bit_Index_2_LC_10_21_1  (
            .in0(N__10570),
            .in1(N__10398),
            .in2(N__9715),
            .in3(N__10606),
            .lcout(\c0.tx.r_Bit_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_RNO_0_LC_10_21_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_RNO_0_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Tx_Active_RNO_0_LC_10_21_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.tx.r_Tx_Active_RNO_0_LC_10_21_2  (
            .in0(N__10319),
            .in1(N__9822),
            .in2(_gnd_net_),
            .in3(N__9778),
            .lcout(),
            .ltout(\c0.tx.r_Tx_Active_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_LC_10_21_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_LC_10_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_LC_10_21_3 .LUT_INIT=16'b0000101011111111;
    LogicCell40 \c0.tx.r_Tx_Active_LC_10_21_3  (
            .in0(N__9703),
            .in1(_gnd_net_),
            .in2(N__9712),
            .in3(N__9709),
            .lcout(\c0.tx_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_RNI6GJO_LC_10_21_4 .C_ON=1'b0;
    defparam \c0.tx_active_RNI6GJO_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_active_RNI6GJO_LC_10_21_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \c0.tx_active_RNI6GJO_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__9936),
            .in2(_gnd_net_),
            .in3(N__9701),
            .lcout(\c0.byte_transmit_counter15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_LC_10_21_5 .C_ON=1'b0;
    defparam \c0.tx_transmit_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_LC_10_21_5 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \c0.tx_transmit_LC_10_21_5  (
            .in0(N__9702),
            .in1(_gnd_net_),
            .in2(N__9947),
            .in3(_gnd_net_),
            .lcout(\c0.tx_transmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.N_90_ip_RNI1U1E_LC_10_22_0 .C_ON=1'b0;
    defparam \c0.tx.N_90_ip_RNI1U1E_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.N_90_ip_RNI1U1E_LC_10_22_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.tx.N_90_ip_RNI1U1E_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__9814),
            .in2(_gnd_net_),
            .in3(N__9856),
            .lcout(\c0.tx.N_90_ip_RNI1U1EZ0 ),
            .ltout(\c0.tx.N_90_ip_RNI1U1EZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0_LC_10_22_1 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0_LC_10_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_0_LC_10_22_1 .LUT_INIT=16'b1100000000110000;
    LogicCell40 \c0.tx.r_Bit_Index_0_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__10494),
            .in2(N__9691),
            .in3(N__9735),
            .lcout(\c0.tx.r_Bit_IndexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_4_LC_10_22_2 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_4_LC_10_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_4_LC_10_22_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.tx.r_SM_Main_4_LC_10_22_2  (
            .in0(N__10323),
            .in1(N__9902),
            .in2(_gnd_net_),
            .in3(N__9815),
            .lcout(\c0.tx.r_SM_Main_dup_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNO_0_0_LC_10_22_3 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNO_0_0_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNO_0_0_LC_10_22_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.tx.r_SM_Main_RNO_0_0_LC_10_22_3  (
            .in0(N__10318),
            .in1(N__10648),
            .in2(N__9957),
            .in3(N__10537),
            .lcout(\c0.tx.r_SM_Main_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_1_LC_10_22_4 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_1_LC_10_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_1_LC_10_22_4 .LUT_INIT=16'b1001110000000000;
    LogicCell40 \c0.tx.r_Bit_Index_1_LC_10_22_4  (
            .in0(N__9736),
            .in1(N__10605),
            .in2(N__10503),
            .in3(N__10399),
            .lcout(\c0.tx.r_Bit_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNO_0_2_LC_10_22_5 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNO_0_2_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNO_0_2_LC_10_22_5 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \c0.tx.r_SM_Main_RNO_0_2_LC_10_22_5  (
            .in0(N__9901),
            .in1(N__10649),
            .in2(_gnd_net_),
            .in3(N__10538),
            .lcout(),
            .ltout(\c0.tx.r_SM_Main_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_2_LC_10_22_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_2_LC_10_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_2_LC_10_22_6 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \c0.tx.r_SM_Main_2_LC_10_22_6  (
            .in0(N__10468),
            .in1(N__9903),
            .in2(N__9886),
            .in3(N__9816),
            .lcout(\c0.tx.r_SM_Main_dup_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNIVDI71_2_LC_10_22_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNIVDI71_2_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNIVDI71_2_LC_10_22_7 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \c0.tx.r_SM_Main_RNIVDI71_2_LC_10_22_7  (
            .in0(N__9857),
            .in1(N__10647),
            .in2(N__9823),
            .in3(N__9771),
            .lcout(\c0.tx.r_SM_Main_RNIVDI71Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__7_LC_10_23_1 .C_ON=1'b0;
    defparam \c0.data_out_0__7_LC_10_23_1 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__7_LC_10_23_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_0__7_LC_10_23_1  (
            .in0(N__16958),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19624),
            .ce(),
            .sr(N__16879));
    defparam \c0.data_out_2__4_LC_10_23_2 .C_ON=1'b0;
    defparam \c0.data_out_2__4_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__4_LC_10_23_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_out_2__4_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__16960),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19624),
            .ce(),
            .sr(N__16879));
    defparam \c0.data_out_1__7_LC_10_23_3 .C_ON=1'b0;
    defparam \c0.data_out_1__7_LC_10_23_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__7_LC_10_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_1__7_LC_10_23_3  (
            .in0(N__16959),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19624),
            .ce(),
            .sr(N__16879));
    defparam \c0.data_out_0__0_LC_10_23_4 .C_ON=1'b0;
    defparam \c0.data_out_0__0_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__0_LC_10_23_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_out_0__0_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__16955),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19624),
            .ce(),
            .sr(N__16879));
    defparam \c0.data_out_0__1_LC_10_23_5 .C_ON=1'b0;
    defparam \c0.data_out_0__1_LC_10_23_5 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__1_LC_10_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_0__1_LC_10_23_5  (
            .in0(N__16956),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19624),
            .ce(),
            .sr(N__16879));
    defparam \c0.data_out_0__4_LC_10_23_6 .C_ON=1'b0;
    defparam \c0.data_out_0__4_LC_10_23_6 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__4_LC_10_23_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_out_0__4_LC_10_23_6  (
            .in0(_gnd_net_),
            .in1(N__16957),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19624),
            .ce(),
            .sr(N__16879));
    defparam \c0.data_out_2__7_LC_10_23_7 .C_ON=1'b0;
    defparam \c0.data_out_2__7_LC_10_23_7 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__7_LC_10_23_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_2__7_LC_10_23_7  (
            .in0(N__16961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19624),
            .ce(),
            .sr(N__16879));
    defparam CONSTANT_ONE_LUT4_LC_10_24_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_24_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_24_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_2_LC_10_24_2 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_2_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_2_LC_10_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__RNO_0_2_LC_10_24_2  (
            .in0(N__14466),
            .in1(N__12086),
            .in2(_gnd_net_),
            .in3(N__13328),
            .lcout(\c0.nextCRC16_3_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNINVK01_8_LC_10_24_3 .C_ON=1'b0;
    defparam \c0.d_2_RNINVK01_8_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNINVK01_8_LC_10_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNINVK01_8_LC_10_24_3  (
            .in0(N__12637),
            .in1(N__13009),
            .in2(_gnd_net_),
            .in3(N__11862),
            .lcout(\c0.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIIQK01_7_LC_10_24_6 .C_ON=1'b0;
    defparam \c0.d_2_RNIIQK01_7_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIIQK01_7_LC_10_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNIIQK01_7_LC_10_24_6  (
            .in0(N__10895),
            .in1(N__11427),
            .in2(_gnd_net_),
            .in3(N__13327),
            .lcout(\c0.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIQ3DA1_20_LC_10_24_7 .C_ON=1'b0;
    defparam \c0.d_2_RNIQ3DA1_20_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIQ3DA1_20_LC_10_24_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIQ3DA1_20_LC_10_24_7  (
            .in0(N__11513),
            .in1(N__14465),
            .in2(N__12090),
            .in3(N__14497),
            .lcout(\c0.nextCRC16_3_0_a2_6_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__1_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.data_out_7__1_LC_10_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__1_LC_10_25_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__1_LC_10_25_0  (
            .in0(N__10674),
            .in1(N__10789),
            .in2(N__12850),
            .in3(N__10071),
            .lcout(\c0.data_out_7_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19639),
            .ce(N__16832),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNI9INJ_33_LC_10_25_1 .C_ON=1'b0;
    defparam \c0.d_2_RNI9INJ_33_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNI9INJ_33_LC_10_25_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.d_2_RNI9INJ_33_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(N__11762),
            .in2(_gnd_net_),
            .in3(N__11790),
            .lcout(\c0.N_24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNID5VK2_21_LC_10_25_2 .C_ON=1'b0;
    defparam \c0.d_2_RNID5VK2_21_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNID5VK2_21_LC_10_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNID5VK2_21_LC_10_25_2  (
            .in0(N__9998),
            .in1(N__11992),
            .in2(N__14873),
            .in3(N__10022),
            .lcout(),
            .ltout(\c0.nextCRC16_3_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIKDAK6_20_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.d_2_RNIKDAK6_20_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIKDAK6_20_LC_10_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIKDAK6_20_LC_10_25_3  (
            .in0(N__10102),
            .in1(N__12013),
            .in2(N__10096),
            .in3(N__10083),
            .lcout(\c0.N_106 ),
            .ltout(\c0.N_106_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__7_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.data_out_6__7_LC_10_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__7_LC_10_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_6__7_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(N__10822),
            .in2(N__10093),
            .in3(N__10788),
            .lcout(\c0.data_out_6_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19639),
            .ce(N__16832),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNITDBK1_19_LC_10_25_5 .C_ON=1'b0;
    defparam \c0.d_2_RNITDBK1_19_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNITDBK1_19_LC_10_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNITDBK1_19_LC_10_25_5  (
            .in0(N__10440),
            .in1(N__12803),
            .in2(N__13361),
            .in3(N__11588),
            .lcout(\c0.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__0_LC_10_25_6 .C_ON=1'b0;
    defparam \c0.data_out_7__0_LC_10_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__0_LC_10_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__0_LC_10_25_6  (
            .in0(N__10675),
            .in1(N__10717),
            .in2(N__10909),
            .in3(N__10072),
            .lcout(\c0.data_out_7_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19639),
            .ce(N__16832),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__2_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.data_out_6__2_LC_10_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__2_LC_10_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__2_LC_10_26_0  (
            .in0(N__13399),
            .in1(N__13485),
            .in2(N__10054),
            .in3(N__10005),
            .lcout(\c0.data_out_6_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19647),
            .ce(N__16829),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__4_LC_10_26_5 .C_ON=1'b0;
    defparam \c0.data_out_4__4_LC_10_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__4_LC_10_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__4_LC_10_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10042),
            .lcout(\c0.d_2_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19647),
            .ce(N__16829),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__1_LC_10_27_0 .C_ON=1'b0;
    defparam \c0.data_out_6__1_LC_10_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__1_LC_10_27_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__1_LC_10_27_0  (
            .in0(N__14874),
            .in1(N__10027),
            .in2(N__11998),
            .in3(N__10006),
            .lcout(\c0.data_out_6_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19653),
            .ce(N__16827),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__0_LC_10_27_1 .C_ON=1'b0;
    defparam \c0.data_out_5__0_LC_10_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__0_LC_10_27_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_out_5__0_LC_10_27_1  (
            .in0(_gnd_net_),
            .in1(N__10186),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19653),
            .ce(N__16827),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__6_LC_10_27_2 .C_ON=1'b0;
    defparam \c0.data_out_4__6_LC_10_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__6_LC_10_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__6_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10174),
            .lcout(\c0.d_2_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19653),
            .ce(N__16827),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__3_LC_10_27_3 .C_ON=1'b0;
    defparam \c0.data_out_4__3_LC_10_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__3_LC_10_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__3_LC_10_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10162),
            .lcout(\c0.d_2_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19653),
            .ce(N__16827),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__2_LC_10_27_4 .C_ON=1'b0;
    defparam \c0.data_out_5__2_LC_10_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__2_LC_10_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__2_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10150),
            .lcout(\c0.d_2_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19653),
            .ce(N__16827),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__7_LC_10_27_6 .C_ON=1'b0;
    defparam \c0.data_out_4__7_LC_10_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__7_LC_10_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__7_LC_10_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10138),
            .lcout(\c0.d_2_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19653),
            .ce(N__16827),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__4_LC_10_27_7 .C_ON=1'b0;
    defparam \c0.data_out_5__4_LC_10_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__4_LC_10_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__4_LC_10_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10126),
            .lcout(\c0.d_2_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19653),
            .ce(N__16827),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__0_LC_10_28_4 .C_ON=1'b0;
    defparam \c0.data_out_4__0_LC_10_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__0_LC_10_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__0_LC_10_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10114),
            .lcout(\c0.d_2_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19662),
            .ce(N__16825),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__0_LC_11_17_1 .C_ON=1'b0;
    defparam \c0.data_in_5__0_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__0_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__0_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10931),
            .lcout(\c0.data_in_5_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19592),
            .ce(N__17717),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__7_LC_11_17_2 .C_ON=1'b0;
    defparam \c0.data_in_4__7_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__7_LC_11_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__7_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12150),
            .lcout(\c0.data_in_4_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19592),
            .ce(N__17717),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__3_LC_11_17_4 .C_ON=1'b0;
    defparam \c0.data_in_4__3_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__3_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__3_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11230),
            .lcout(\c0.data_in_4_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19592),
            .ce(N__17717),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__7_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.data_in_5__7_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__7_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__7_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13584),
            .lcout(\c0.data_in_5_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19592),
            .ce(N__17717),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__2_LC_11_17_6 .C_ON=1'b0;
    defparam \c0.data_in_5__2_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__2_LC_11_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__2_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17761),
            .lcout(\c0.data_in_5_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19592),
            .ce(N__17717),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__0_LC_11_17_7 .C_ON=1'b0;
    defparam \c0.data_in_6__0_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__0_LC_11_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__0_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17369),
            .lcout(\c0.data_in_6_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19592),
            .ce(N__17717),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__1_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.data_in_5__1_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__1_LC_11_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__1_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13640),
            .lcout(\c0.data_in_5_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19599),
            .ce(N__17720),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__1_LC_11_18_1 .C_ON=1'b0;
    defparam \c0.data_in_4__1_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__1_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__1_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12288),
            .lcout(\c0.data_in_4_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19599),
            .ce(N__17720),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__1_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.data_in_6__1_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__1_LC_11_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__1_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17337),
            .lcout(\c0.data_in_6_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19599),
            .ce(N__17720),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__3_LC_11_18_3 .C_ON=1'b0;
    defparam \c0.data_in_2__3_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__3_LC_11_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__3_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12386),
            .lcout(\c0.data_in_2_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19599),
            .ce(N__17720),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__3_LC_11_18_4 .C_ON=1'b0;
    defparam \c0.data_in_6__3_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__3_LC_11_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__3_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11386),
            .lcout(\c0.data_in_6_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19599),
            .ce(N__17720),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__2_LC_11_18_5 .C_ON=1'b0;
    defparam \c0.data_in_4__2_LC_11_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__2_LC_11_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__2_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12519),
            .lcout(\c0.data_in_4_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19599),
            .ce(N__17720),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__1_LC_11_18_6 .C_ON=1'b0;
    defparam \c0.data_in_3__1_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__1_LC_11_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__1_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11031),
            .lcout(\c0.data_in_3_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19599),
            .ce(N__17720),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__4_LC_11_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__4_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__4_LC_11_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__4_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10261),
            .lcout(\c0.d_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19604),
            .ce(N__17185),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__3_LC_11_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__3_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__3_LC_11_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__3_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11381),
            .lcout(\c0.data_in_frame_7_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19604),
            .ce(N__17185),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__0_LC_11_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__0_LC_11_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__0_LC_11_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__0_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10243),
            .lcout(\c0.d_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19604),
            .ce(N__17185),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__1_LC_11_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__1_LC_11_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__1_LC_11_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__1_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13641),
            .lcout(\c0.data_in_frame_6_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19604),
            .ce(N__17185),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__1_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.data_in_2__1_LC_11_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__1_LC_11_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__1_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15849),
            .lcout(\c0.data_in_2_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19612),
            .ce(N__17724),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__3_LC_11_20_1 .C_ON=1'b0;
    defparam \c0.data_in_3__3_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__3_LC_11_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__3_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12139),
            .lcout(\c0.data_in_3_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19612),
            .ce(N__17724),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__3_LC_11_20_3 .C_ON=1'b0;
    defparam \c0.data_in_7__3_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__3_LC_11_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__3_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10225),
            .lcout(\c0.data_in_7_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19612),
            .ce(N__17724),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__7_LC_11_20_4 .C_ON=1'b0;
    defparam \c0.data_in_6__7_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__7_LC_11_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__7_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13552),
            .lcout(\c0.data_in_6_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19612),
            .ce(N__17724),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__1_LC_11_20_5 .C_ON=1'b0;
    defparam \c0.data_in_7__1_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__1_LC_11_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__1_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10207),
            .lcout(\c0.data_in_7_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19612),
            .ce(N__17724),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__0_LC_11_20_6 .C_ON=1'b0;
    defparam \c0.data_in_7__0_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__0_LC_11_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__0_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10420),
            .lcout(\c0.data_in_7_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19612),
            .ce(N__17724),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__3_LC_11_20_7 .C_ON=1'b0;
    defparam \c0.data_in_5__3_LC_11_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__3_LC_11_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__3_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11310),
            .lcout(\c0.data_in_5_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19612),
            .ce(N__17724),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_5_LC_11_21_4 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_5_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_5_LC_11_21_4 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_5_LC_11_21_4  (
            .in0(N__13174),
            .in1(N__10566),
            .in2(N__11398),
            .in3(N__10599),
            .lcout(),
            .ltout(\c0.tx.o_Tx_Serial_2_3_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_3_LC_11_21_5 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_3_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_3_LC_11_21_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_3_LC_11_21_5  (
            .in0(N__10600),
            .in1(N__14299),
            .in2(N__10402),
            .in3(N__13156),
            .lcout(\c0.tx.o_Tx_Serial_RNO_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_0_LC_11_21_6 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_0_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_0_LC_11_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_0_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10397),
            .lcout(\c0.tx.N_390_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_4_LC_11_22_0 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_4_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_4_LC_11_22_0 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_4_LC_11_22_0  (
            .in0(N__10567),
            .in1(N__13096),
            .in2(N__11608),
            .in3(N__10601),
            .lcout(),
            .ltout(\c0.tx.o_Tx_Serial_2_6_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_2_LC_11_22_1 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_2_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_2_LC_11_22_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_2_LC_11_22_1  (
            .in0(N__10602),
            .in1(N__11404),
            .in2(N__10381),
            .in3(N__11440),
            .lcout(),
            .ltout(\c0.tx.o_Tx_Serial_RNO_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_1_LC_11_22_2 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_1_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_1_LC_11_22_2 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_1_LC_11_22_2  (
            .in0(N__10498),
            .in1(N__10378),
            .in2(N__10372),
            .in3(N__10654),
            .lcout(),
            .ltout(\c0.tx.o_Tx_Serial_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_LC_11_22_3 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_LC_11_22_3 .SEQ_MODE=4'b1001;
    defparam \c0.tx.o_Tx_Serial_LC_11_22_3 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \c0.tx.o_Tx_Serial_LC_11_22_3  (
            .in0(N__10272),
            .in1(N__10356),
            .in2(N__10327),
            .in3(N__10324),
            .lcout(PIN_1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19625),
            .ce(),
            .sr(N__10666));
    defparam \c0.tx.r_SM_Main_RNO_0_3_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNO_0_3_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNO_0_3_LC_11_22_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.r_SM_Main_RNO_0_3_LC_11_22_6  (
            .in0(N__10568),
            .in1(N__10603),
            .in2(N__10504),
            .in3(N__10653),
            .lcout(\c0.tx.r_SM_Main_recr_i_0_a2_0_2_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNO_1_2_LC_11_22_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNO_1_2_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNO_1_2_LC_11_22_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.tx.r_SM_Main_RNO_1_2_LC_11_22_7  (
            .in0(N__10604),
            .in1(N__10569),
            .in2(N__10546),
            .in3(N__10502),
            .lcout(\c0.tx.r_SM_Main_recr_i_i_a2_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__5_LC_11_23_0 .C_ON=1'b0;
    defparam \c0.data_out_7__5_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__5_LC_11_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__5_LC_11_23_0  (
            .in0(N__10834),
            .in1(N__10765),
            .in2(N__10450),
            .in3(N__11598),
            .lcout(\c0.data_out_7_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19633),
            .ce(N__16835),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_5_LC_11_23_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_5_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_5_LC_11_23_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx_data_RNO_1_5_LC_11_23_1  (
            .in0(N__15373),
            .in1(N__10459),
            .in2(N__15568),
            .in3(N__10846),
            .lcout(\c0.tx_data_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_3_LC_11_23_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_3_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_3_LC_11_23_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_3_3_LC_11_23_2  (
            .in0(N__10780),
            .in1(N__15558),
            .in2(N__14830),
            .in3(N__15371),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_3_LC_11_23_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_3_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_3_LC_11_23_3 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_3_LC_11_23_3  (
            .in0(N__15197),
            .in1(N__15652),
            .in2(N__10453),
            .in3(N__10426),
            .lcout(\c0.tx_data_1_0_i_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_3_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_3_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_3_LC_11_23_4 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_4_3_LC_11_23_4  (
            .in0(N__10446),
            .in1(N__15557),
            .in2(N__10711),
            .in3(N__15370),
            .lcout(\c0.tx_data_RNO_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_3_LC_11_23_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_3_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_3_LC_11_23_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx_data_RNO_0_3_LC_11_23_5  (
            .in0(N__15372),
            .in1(N__11711),
            .in2(N__15567),
            .in3(N__10900),
            .lcout(\c0.tx_data_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_2_0_LC_11_23_7 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_2_0_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_2_0_LC_11_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_7__RNO_2_0_LC_11_23_7  (
            .in0(N__11824),
            .in1(N__11710),
            .in2(_gnd_net_),
            .in3(N__11741),
            .lcout(\c0.nextCRC16_3_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_2_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_2_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_2_LC_11_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_0_2_LC_11_24_0  (
            .in0(N__11831),
            .in1(N__12832),
            .in2(N__12942),
            .in3(N__11649),
            .lcout(),
            .ltout(\c0.nextCRC16_3_0_a2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__2_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.data_out_7__2_LC_11_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__2_LC_11_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__2_LC_11_24_1  (
            .in0(N__10803),
            .in1(N__15030),
            .in2(N__10750),
            .in3(N__11671),
            .lcout(\c0.data_out_7_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19640),
            .ce(N__16833),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__6_LC_11_24_2 .C_ON=1'b0;
    defparam \c0.data_out_5__6_LC_11_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__6_LC_11_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__6_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10747),
            .lcout(\c0.d_2_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19640),
            .ce(N__16833),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIFMJ01_45_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.d_2_RNIFMJ01_45_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIFMJ01_45_LC_11_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNIFMJ01_45_LC_11_24_3  (
            .in0(N__12984),
            .in1(N__14934),
            .in2(_gnd_net_),
            .in3(N__12864),
            .lcout(\c0.N_99 ),
            .ltout(\c0.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_3_0_LC_11_24_4 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_3_0_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_3_0_LC_11_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_3_0_LC_11_24_4  (
            .in0(N__14993),
            .in1(N__13039),
            .in2(N__10729),
            .in3(N__10802),
            .lcout(),
            .ltout(\c0.nextCRC16_3_0_a2_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_1_0_LC_11_24_5 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_1_0_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_1_0_LC_11_24_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_1_0_LC_11_24_5  (
            .in0(N__10726),
            .in1(N__12775),
            .in2(N__10720),
            .in3(N__14793),
            .lcout(\c0.nextCRC16_3_0_a2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIDLMJ_16_LC_11_24_6 .C_ON=1'b0;
    defparam \c0.d_2_RNIDLMJ_16_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIDLMJ_16_LC_11_24_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.d_2_RNIDLMJ_16_LC_11_24_6  (
            .in0(N__14959),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12602),
            .lcout(\c0.N_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIM3JT_12_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.d_2_RNIM3JT_12_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIM3JT_12_LC_11_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNIM3JT_12_LC_11_25_2  (
            .in0(N__12035),
            .in1(N__14894),
            .in2(_gnd_net_),
            .in3(N__11947),
            .lcout(\c0.N_81 ),
            .ltout(\c0.N_81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNII92R1_27_LC_11_25_3 .C_ON=1'b0;
    defparam \c0.d_2_RNII92R1_27_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNII92R1_27_LC_11_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNII92R1_27_LC_11_25_3  (
            .in0(N__10710),
            .in1(N__13136),
            .in2(N__10678),
            .in3(N__14819),
            .lcout(\c0.N_105 ),
            .ltout(\c0.N_105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__5_LC_11_25_4 .C_ON=1'b0;
    defparam \c0.data_out_6__5_LC_11_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__5_LC_11_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_6__5_LC_11_25_4  (
            .in0(_gnd_net_),
            .in1(N__12933),
            .in2(N__10849),
            .in3(N__13404),
            .lcout(\c0.data_out_6_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19648),
            .ce(N__16830),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_1_7_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_1_7_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_1_7_LC_11_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__RNO_1_7_LC_11_25_5  (
            .in0(N__11740),
            .in1(N__11835),
            .in2(N__12941),
            .in3(N__14789),
            .lcout(),
            .ltout(\c0.nextCRC16_3_0_a2_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_7_LC_11_25_6 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_7_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_7_LC_11_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__RNO_0_7_LC_11_25_6  (
            .in0(N__10816),
            .in1(N__11666),
            .in2(N__10837),
            .in3(N__10833),
            .lcout(\c0.nextCRC16_3_0_a2_5_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_2_7_LC_11_25_7 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_2_7_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_2_7_LC_11_25_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__RNO_2_7_LC_11_25_7  (
            .in0(N__14895),
            .in1(N__13135),
            .in2(N__11955),
            .in3(N__14818),
            .lcout(\c0.nextCRC16_3_0_a2_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIJ2812_44_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.d_2_RNIJ2812_44_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIJ2812_44_LC_11_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIJ2812_44_LC_11_26_0  (
            .in0(N__14747),
            .in1(N__13293),
            .in2(N__13448),
            .in3(N__10761),
            .lcout(\c0.N_95 ),
            .ltout(\c0.N_95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIJDOU2_14_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.d_2_RNIJDOU2_14_LC_11_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIJDOU2_14_LC_11_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.d_2_RNIJDOU2_14_LC_11_26_1  (
            .in0(_gnd_net_),
            .in1(N__15031),
            .in2(N__10810),
            .in3(N__10807),
            .lcout(\c0.nextCRC16_3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__7_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.data_out_3__7_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__7_LC_11_26_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_3__7_LC_11_26_2  (
            .in0(N__17020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19654),
            .ce(),
            .sr(N__16877));
    defparam \c0.data_out_0__3_LC_11_26_3 .C_ON=1'b0;
    defparam \c0.data_out_0__3_LC_11_26_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__3_LC_11_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__3_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17019),
            .lcout(\c0.d_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19654),
            .ce(),
            .sr(N__16877));
    defparam \c0.d_2_RNI6EK01_3_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.d_2_RNI6EK01_3_LC_11_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNI6EK01_3_LC_11_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNI6EK01_3_LC_11_26_4  (
            .in0(N__12114),
            .in1(N__11638),
            .in2(_gnd_net_),
            .in3(N__10776),
            .lcout(\c0.N_75 ),
            .ltout(\c0.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_0_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_0_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_0_LC_11_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_7__RNO_0_0_LC_11_26_5  (
            .in0(_gnd_net_),
            .in1(N__13441),
            .in2(N__10912),
            .in3(N__14748),
            .lcout(\c0.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__2_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.data_out_0__2_LC_11_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__2_LC_11_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__2_LC_11_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17018),
            .lcout(\c0.d_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19654),
            .ce(),
            .sr(N__16877));
    defparam \c0.data_out_6__RNO_0_4_LC_11_27_0 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_4_LC_11_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_4_LC_11_27_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_6__RNO_0_4_LC_11_27_0  (
            .in0(_gnd_net_),
            .in1(N__11940),
            .in2(_gnd_net_),
            .in3(N__13395),
            .lcout(\c0.nextCRC16_3_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_6_LC_11_27_1 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_6_LC_11_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_6_LC_11_27_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_7__RNO_0_6_LC_11_27_1  (
            .in0(_gnd_net_),
            .in1(N__12113),
            .in2(_gnd_net_),
            .in3(N__10894),
            .lcout(\c0.un144_newcrc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__1_LC_11_28_4 .C_ON=1'b0;
    defparam \c0.data_out_3__1_LC_11_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__1_LC_11_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__1_LC_11_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.d_2_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19668),
            .ce(),
            .sr(N__16873));
    defparam \c0.data_out_3__0_LC_11_28_7 .C_ON=1'b0;
    defparam \c0.data_out_3__0_LC_11_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__0_LC_11_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__0_LC_11_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.d_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19668),
            .ce(),
            .sr(N__16873));
    defparam \c0.data_in_7__7_LC_12_16_5 .C_ON=1'b0;
    defparam \c0.data_in_7__7_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__7_LC_12_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__7_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10870),
            .lcout(\c0.data_in_7_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19605),
            .ce(N__17722),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__5_LC_12_16_7 .C_ON=1'b0;
    defparam \c0.data_in_4__5_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__5_LC_12_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__5_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11877),
            .lcout(\c0.data_in_4_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19605),
            .ce(N__17722),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__5_LC_12_17_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__5_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__5_LC_12_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__5_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11878),
            .lcout(\c0.d_4_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19597),
            .ce(N__17177),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__6_LC_12_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__6_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__6_LC_12_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__6_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16087),
            .lcout(\c0.d_4_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19597),
            .ce(N__17177),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__0_LC_12_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__0_LC_12_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__0_LC_12_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__0_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10932),
            .lcout(\c0.data_in_frame_6_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19597),
            .ce(N__17177),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__5_LC_12_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__5_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__5_LC_12_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__5_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11020),
            .lcout(\c0.d_4_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19597),
            .ce(N__17177),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__2_LC_12_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__2_LC_12_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__2_LC_12_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__2_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17757),
            .lcout(\c0.data_in_frame_6_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19597),
            .ce(N__17177),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__3_LC_12_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__3_LC_12_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__3_LC_12_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__3_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10992),
            .lcout(\c0.d_4_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19597),
            .ce(N__17177),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__2_LC_12_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__2_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__2_LC_12_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__2_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17775),
            .lcout(\c0.data_in_frame_7_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19597),
            .ce(N__17177),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNINGK21_21_LC_12_18_0 .C_ON=1'b0;
    defparam \c0.d_4_RNINGK21_21_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNINGK21_21_LC_12_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNINGK21_21_LC_12_18_0  (
            .in0(N__17582),
            .in1(N__18869),
            .in2(N__14394),
            .in3(N__13688),
            .lcout(\c0.N_126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__7_LC_12_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__7_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__7_LC_12_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__7_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10975),
            .lcout(\c0.d_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19606),
            .ce(N__17181),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__7_LC_12_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__7_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__7_LC_12_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__7_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10957),
            .lcout(\c0.d_4_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19606),
            .ce(N__17181),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIT2KP_20_LC_12_18_3 .C_ON=1'b0;
    defparam \c0.d_4_RNIT2KP_20_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIT2KP_20_LC_12_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIT2KP_20_LC_12_18_3  (
            .in0(N__13689),
            .in1(N__12193),
            .in2(N__10933),
            .in3(N__17960),
            .lcout(\c0.un1_data_in_6__0_0_a2_5_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__4_LC_12_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__4_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__4_LC_12_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__4_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11203),
            .lcout(\c0.d_4_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19606),
            .ce(N__17181),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__2_LC_12_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__2_LC_12_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__2_LC_12_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_frame_4__2_LC_12_18_5  (
            .in0(N__11182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19606),
            .ce(N__17181),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIQ7PC_23_LC_12_18_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIQ7PC_23_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIQ7PC_23_LC_12_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIQ7PC_23_LC_12_18_6  (
            .in0(N__14390),
            .in1(N__16437),
            .in2(N__17649),
            .in3(N__11303),
            .lcout(\c0.un1_data_in_6__3_0_a2_5_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__5_LC_12_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__5_LC_12_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__5_LC_12_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__5_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11166),
            .lcout(\c0.d_4_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19606),
            .ce(N__17181),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__0_LC_12_19_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__0_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__0_LC_12_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__0_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11149),
            .lcout(\c0.d_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19613),
            .ce(N__17182),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__3_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__3_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__3_LC_12_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__3_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11131),
            .lcout(\c0.d_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19613),
            .ce(N__17182),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__7_LC_12_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__7_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__7_LC_12_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__7_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11104),
            .lcout(\c0.d_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19613),
            .ce(N__17182),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__0_LC_12_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__0_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__0_LC_12_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__0_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11083),
            .lcout(\c0.d_4_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19613),
            .ce(N__17182),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__5_LC_12_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__5_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__5_LC_12_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__5_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11056),
            .lcout(\c0.d_4_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19613),
            .ce(N__17182),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__1_LC_12_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__1_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__1_LC_12_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__1_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11032),
            .lcout(\c0.d_4_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19613),
            .ce(N__17182),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__7_LC_12_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__7_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__7_LC_12_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__7_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11245),
            .lcout(\c0.d_4_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19613),
            .ce(N__17182),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__3_LC_12_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__3_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__3_LC_12_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__3_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11226),
            .lcout(\c0.d_4_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19613),
            .ce(N__17182),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI5L571_45_LC_12_20_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI5L571_45_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI5L571_45_LC_12_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI5L571_45_LC_12_20_0  (
            .in0(N__17676),
            .in1(N__12738),
            .in2(N__11284),
            .in3(N__14612),
            .lcout(\c0.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIH9JJ_4_LC_12_20_1 .C_ON=1'b0;
    defparam \c0.d_4_RNIH9JJ_4_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIH9JJ_4_LC_12_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNIH9JJ_4_LC_12_20_1  (
            .in0(N__12198),
            .in1(N__18054),
            .in2(_gnd_net_),
            .in3(N__12472),
            .lcout(\c0.N_108 ),
            .ltout(\c0.N_108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNICGS41_17_LC_12_20_2 .C_ON=1'b0;
    defparam \c0.d_4_RNICGS41_17_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNICGS41_17_LC_12_20_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.d_4_RNICGS41_17_LC_12_20_2  (
            .in0(N__11281),
            .in1(_gnd_net_),
            .in2(N__11215),
            .in3(N__14613),
            .lcout(),
            .ltout(\c0.N_122_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIJUS53_16_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.d_4_RNIJUS53_16_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIJUS53_16_LC_12_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIJUS53_16_LC_12_20_3  (
            .in0(N__16545),
            .in1(N__12259),
            .in2(N__11212),
            .in3(N__12550),
            .lcout(\c0.un1_data_in_7__1_0_a2_24_a2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIVCPC_26_LC_12_20_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIVCPC_26_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIVCPC_26_LC_12_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIVCPC_26_LC_12_20_4  (
            .in0(N__13927),
            .in1(N__17606),
            .in2(N__13583),
            .in3(N__16046),
            .lcout(),
            .ltout(\c0.un1_data_in_6__7_0_a2_17_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIIAP41_26_LC_12_20_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIIAP41_26_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIIAP41_26_LC_12_20_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.d_4_RNIIAP41_26_LC_12_20_5  (
            .in0(N__16301),
            .in1(_gnd_net_),
            .in2(N__11209),
            .in3(N__13801),
            .lcout(),
            .ltout(\c0.un1_data_in_6__7_0_a2_17_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIP5RG3_15_LC_12_20_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIP5RG3_15_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIP5RG3_15_LC_12_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIP5RG3_15_LC_12_20_6  (
            .in0(N__16501),
            .in1(N__16546),
            .in2(N__11206),
            .in3(N__16157),
            .lcout(\c0.un1_data_in_6__7_0_a2_17_a2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIN7VG_47_LC_12_21_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIN7VG_47_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIN7VG_47_LC_12_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIN7VG_47_LC_12_21_0  (
            .in0(N__11282),
            .in1(N__18095),
            .in2(N__11385),
            .in3(N__17514),
            .lcout(\c0.un1_data_in_7__3_0_a2_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__1_LC_12_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__1_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__1_LC_12_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__1_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11362),
            .lcout(\c0.d_4_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19626),
            .ce(N__17187),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__6_LC_12_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__6_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__6_LC_12_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__6_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11344),
            .lcout(\c0.d_4_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19626),
            .ce(N__17187),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_3_LC_12_21_4 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_3_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_3_LC_12_21_4 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx2_data_RNO_1_3_LC_12_21_4  (
            .in0(N__18361),
            .in1(N__11290),
            .in2(N__11323),
            .in3(N__18571),
            .lcout(\c0.tx2_data_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__3_LC_12_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__3_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__3_LC_12_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__3_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11311),
            .lcout(\c0.data_in_frame_6_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19626),
            .ce(N__17187),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_1_LC_12_21_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_1_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_1_LC_12_21_6 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \c0.tx2_data_RNO_4_1_LC_12_21_6  (
            .in0(N__11283),
            .in1(N__18572),
            .in2(N__18374),
            .in3(N__15826),
            .lcout(\c0.tx2_data_RNO_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_1_LC_12_22_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_1_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_1_LC_12_22_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \c0.tx2_data_RNO_2_1_LC_12_22_2  (
            .in0(N__16633),
            .in1(N__18715),
            .in2(N__11263),
            .in3(N__18799),
            .lcout(),
            .ltout(\c0.m161_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_1_LC_12_22_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_1_LC_12_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_1_LC_12_22_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx2.r_Tx_Data_1_LC_12_22_3  (
            .in0(N__18716),
            .in1(N__16597),
            .in2(N__11254),
            .in3(N__11251),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19634),
            .ce(N__19978),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_1_LC_12_22_4 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_1_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_1_LC_12_22_4 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \c0.tx2_data_RNO_0_1_LC_12_22_4  (
            .in0(N__15985),
            .in1(N__18578),
            .in2(N__18376),
            .in3(N__12479),
            .lcout(\c0.tx2_data_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_2_LC_12_22_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_2_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_2_LC_12_22_5 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \c0.tx2_data_RNO_0_2_LC_12_22_5  (
            .in0(N__16336),
            .in1(N__18370),
            .in2(N__18594),
            .in3(N__12199),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_2_LC_12_22_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_2_LC_12_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_2_LC_12_22_6 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \c0.tx2.r_Tx_Data_2_LC_12_22_6  (
            .in0(N__11458),
            .in1(N__14335),
            .in2(N__11485),
            .in3(N__18717),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19634),
            .ce(N__19978),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_2_LC_12_22_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_2_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_2_LC_12_22_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx2_data_RNO_1_2_LC_12_22_7  (
            .in0(N__18577),
            .in1(N__11482),
            .in2(N__11470),
            .in3(N__18369),
            .lcout(\c0.tx2_data_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_7_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_7_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_7_LC_12_23_0 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \c0.tx_data_RNO_4_7_LC_12_23_0  (
            .in0(N__11650),
            .in1(N__15565),
            .in2(N__11997),
            .in3(N__15374),
            .lcout(\c0.tx_data_RNO_4Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_3_LC_12_23_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_3_LC_12_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_3_LC_12_23_1 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \c0.tx.r_Tx_Data_3_LC_12_23_1  (
            .in0(N__11452),
            .in1(N__13216),
            .in2(N__15212),
            .in3(N__11446),
            .lcout(\c0.tx.r_Tx_DataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19641),
            .ce(N__14279),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_7_LC_12_23_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_7_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_7_LC_12_23_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_3_7_LC_12_23_2  (
            .in0(N__11431),
            .in1(N__15566),
            .in2(N__11749),
            .in3(N__15375),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_7_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_7_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_7_LC_12_23_3 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_7_LC_12_23_3  (
            .in0(N__15198),
            .in1(N__15658),
            .in2(N__11416),
            .in3(N__11413),
            .lcout(),
            .ltout(\c0.tx_data_1_0_i_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_7_LC_12_23_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_7_LC_12_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_7_LC_12_23_4 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \c0.tx.r_Tx_Data_7_LC_12_23_4  (
            .in0(N__13339),
            .in1(N__15199),
            .in2(N__11407),
            .in3(N__12559),
            .lcout(\c0.tx.r_Tx_DataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19641),
            .ce(N__14279),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_4_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_4_LC_12_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_4_LC_12_23_5 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \c0.tx.r_Tx_Data_4_LC_12_23_5  (
            .in0(N__13282),
            .in1(N__11890),
            .in2(N__15213),
            .in3(N__11536),
            .lcout(\c0.tx.r_Tx_DataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19641),
            .ce(N__14279),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_5_LC_12_23_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_5_LC_12_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_5_LC_12_23_6 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \c0.tx.r_Tx_Data_5_LC_12_23_6  (
            .in0(N__12961),
            .in1(N__11614),
            .in2(N__15214),
            .in3(N__12751),
            .lcout(\c0.tx.r_Tx_DataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19641),
            .ce(N__14279),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_1_6_LC_12_24_0 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_1_6_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_1_6_LC_12_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_1_6_LC_12_24_0  (
            .in0(N__12811),
            .in1(N__12879),
            .in2(N__11530),
            .in3(N__11599),
            .lcout(),
            .ltout(\c0.un144_newcrc_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__6_LC_12_24_1 .C_ON=1'b0;
    defparam \c0.data_out_7__6_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__6_LC_12_24_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_7__6_LC_12_24_1  (
            .in0(N__11572),
            .in1(N__14749),
            .in2(N__11563),
            .in3(N__12606),
            .lcout(\c0.data_out_7_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19649),
            .ce(N__16831),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_6_LC_12_24_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_6_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_6_LC_12_24_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx_data_RNO_1_6_LC_12_24_2  (
            .in0(N__15346),
            .in1(N__11545),
            .in2(N__11560),
            .in3(N__15531),
            .lcout(\c0.tx_data_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__6_LC_12_24_3 .C_ON=1'b0;
    defparam \c0.data_out_6__6_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__6_LC_12_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__6_LC_12_24_3  (
            .in0(N__12886),
            .in1(N__11551),
            .in2(_gnd_net_),
            .in3(N__11712),
            .lcout(\c0.data_out_6_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19649),
            .ce(N__16831),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_4_LC_12_24_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_4_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_4_LC_12_24_4 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx_data_RNO_3_4_LC_12_24_4  (
            .in0(N__15345),
            .in1(N__12878),
            .in2(N__14902),
            .in3(N__15532),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_4_LC_12_24_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_4_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_4_LC_12_24_5 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_4_LC_12_24_5  (
            .in0(N__15166),
            .in1(N__15657),
            .in2(N__11539),
            .in3(N__11497),
            .lcout(\c0.tx_data_1_0_i_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_4_LC_12_24_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_4_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_4_LC_12_24_6 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \c0.tx_data_RNO_4_4_LC_12_24_6  (
            .in0(N__15344),
            .in1(N__12828),
            .in2(N__11529),
            .in3(N__15530),
            .lcout(\c0.tx_data_RNO_4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__4_LC_12_25_0 .C_ON=1'b0;
    defparam \c0.data_out_7__4_LC_12_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__4_LC_12_25_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_7__4_LC_12_25_0  (
            .in0(N__11491),
            .in1(N__14958),
            .in2(N__15001),
            .in3(N__11797),
            .lcout(\c0.data_out_7_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19655),
            .ce(N__16828),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_0_LC_12_25_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_0_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_0_LC_12_25_1 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \c0.tx_data_RNO_3_0_LC_12_25_1  (
            .in0(N__11866),
            .in1(N__15511),
            .in2(N__11842),
            .in3(N__15341),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_0_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_0_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_0_LC_12_25_2 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_0_LC_12_25_2  (
            .in0(N__15186),
            .in1(N__15656),
            .in2(N__11806),
            .in3(N__11803),
            .lcout(\c0.tx_data_1_0_i_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_0_LC_12_25_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_0_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_0_LC_12_25_3 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_4_0_LC_12_25_3  (
            .in0(N__14957),
            .in1(N__15510),
            .in2(N__12091),
            .in3(N__15340),
            .lcout(\c0.tx_data_RNO_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_1_LC_12_25_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_1_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_1_LC_12_25_4 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx_data_RNO_0_1_LC_12_25_4  (
            .in0(N__15342),
            .in1(N__12036),
            .in2(N__15540),
            .in3(N__11796),
            .lcout(\c0.tx_data_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_2_LC_12_25_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_2_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_2_LC_12_25_5 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \c0.tx_data_RNO_0_2_LC_12_25_5  (
            .in0(N__12934),
            .in1(N__15515),
            .in2(N__11779),
            .in3(N__15343),
            .lcout(\c0.tx_data_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_3_LC_12_26_0 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_3_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_3_LC_12_26_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_7__RNO_0_3_LC_12_26_0  (
            .in0(_gnd_net_),
            .in1(N__13452),
            .in2(_gnd_net_),
            .in3(N__11748),
            .lcout(),
            .ltout(\c0.un105_newcrc_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__3_LC_12_26_1 .C_ON=1'b0;
    defparam \c0.data_out_7__3_LC_12_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__3_LC_12_26_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_7__3_LC_12_26_1  (
            .in0(N__11620),
            .in1(N__11713),
            .in2(N__11674),
            .in3(N__11667),
            .lcout(\c0.data_out_7_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19663),
            .ce(N__16826),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNI9GJ01_29_LC_12_26_2 .C_ON=1'b0;
    defparam \c0.d_2_RNI9GJ01_29_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNI9GJ01_29_LC_12_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNI9GJ01_29_LC_12_26_2  (
            .in0(N__14997),
            .in1(N__16905),
            .in2(_gnd_net_),
            .in3(N__13049),
            .lcout(\c0.N_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_1_3_LC_12_26_3 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_1_3_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_1_3_LC_12_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_1_3_LC_12_26_3  (
            .in0(N__13365),
            .in1(N__12121),
            .in2(N__14938),
            .in3(N__11645),
            .lcout(\c0.un105_newcrc_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_0_LC_12_26_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_0_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_0_LC_12_26_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_0_0_LC_12_26_6  (
            .in0(N__12120),
            .in1(N__15516),
            .in2(N__11959),
            .in3(N__15332),
            .lcout(\c0.tx_data_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_1_4_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_1_4_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_1_4_LC_12_27_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__RNO_1_4_LC_12_27_0  (
            .in0(N__14829),
            .in1(N__15706),
            .in2(N__12082),
            .in3(N__12641),
            .lcout(),
            .ltout(\c0.nextCRC16_3_4_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__4_LC_12_27_1 .C_ON=1'b0;
    defparam \c0.data_out_6__4_LC_12_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__4_LC_12_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__4_LC_12_27_1  (
            .in0(N__14794),
            .in1(N__12049),
            .in2(N__12043),
            .in3(N__12040),
            .lcout(\c0.data_out_6_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19669),
            .ce(N__16824),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIGMI01_10_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.d_2_RNIGMI01_10_LC_12_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIGMI01_10_LC_12_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNIGMI01_10_LC_12_27_4  (
            .in0(N__13400),
            .in1(N__15705),
            .in2(_gnd_net_),
            .in3(N__13489),
            .lcout(\c0.N_94 ),
            .ltout(\c0.N_94_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__3_LC_12_27_5 .C_ON=1'b0;
    defparam \c0.data_out_6__3_LC_12_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__3_LC_12_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__3_LC_12_27_5  (
            .in0(N__12642),
            .in1(N__11917),
            .in2(N__12001),
            .in3(N__13020),
            .lcout(\c0.data_out_6_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19669),
            .ce(N__16824),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_3_LC_12_27_6 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_3_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_3_LC_12_27_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__RNO_0_3_LC_12_27_6  (
            .in0(N__11996),
            .in1(N__13140),
            .in2(_gnd_net_),
            .in3(N__11954),
            .lcout(\c0.nextCRC16_3_0_a2_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_4_LC_12_27_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_4_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_4_LC_12_27_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_1_4_LC_12_27_7  (
            .in0(N__15471),
            .in1(N__11911),
            .in2(N__11905),
            .in3(N__15334),
            .lcout(\c0.tx_data_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__5_LC_13_16_0 .C_ON=1'b0;
    defparam \c0.data_in_5__5_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__5_LC_13_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__5_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17299),
            .lcout(\c0.data_in_5_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19614),
            .ce(N__17725),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__4_LC_13_16_1 .C_ON=1'b0;
    defparam \c0.data_in_7__4_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__4_LC_13_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__4_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12238),
            .lcout(\c0.data_in_7_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19614),
            .ce(N__17725),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__2_LC_13_16_2 .C_ON=1'b0;
    defparam \c0.data_in_7__2_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__2_LC_13_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__2_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12217),
            .lcout(\c0.data_in_7_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19614),
            .ce(N__17725),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__4_LC_13_16_4 .C_ON=1'b0;
    defparam \c0.data_in_4__4_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__4_LC_13_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__4_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12537),
            .lcout(\c0.data_in_4_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19614),
            .ce(N__17725),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__4_LC_13_16_7 .C_ON=1'b0;
    defparam \c0.data_in_5__4_LC_13_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__4_LC_13_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__4_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16015),
            .lcout(\c0.data_in_5_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19614),
            .ce(N__17725),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIJLQL_19_LC_13_17_1 .C_ON=1'b0;
    defparam \c0.d_4_RNIJLQL_19_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIJLQL_19_LC_13_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIJLQL_19_LC_13_17_1  (
            .in0(N__14628),
            .in1(N__14700),
            .in2(N__13750),
            .in3(N__17504),
            .lcout(\c0.N_125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI6FQT_21_LC_13_17_2 .C_ON=1'b0;
    defparam \c0.d_4_RNI6FQT_21_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI6FQT_21_LC_13_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI6FQT_21_LC_13_17_2  (
            .in0(N__17904),
            .in1(N__13903),
            .in2(N__13541),
            .in3(N__17583),
            .lcout(),
            .ltout(\c0.un1_data_in_7__7_0_a2_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI675O1_33_LC_13_17_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI675O1_33_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI675O1_33_LC_13_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI675O1_33_LC_13_17_3  (
            .in0(N__12194),
            .in1(N__12480),
            .in2(N__12169),
            .in3(N__12426),
            .lcout(),
            .ltout(\c0.un1_data_in_7__7_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI8SR93_20_LC_13_17_4 .C_ON=1'b0;
    defparam \c0.d_4_RNI8SR93_20_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI8SR93_20_LC_13_17_4 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \c0.d_4_RNI8SR93_20_LC_13_17_4  (
            .in0(N__12166),
            .in1(N__13732),
            .in2(N__12157),
            .in3(N__16403),
            .lcout(\c0.m163_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__7_LC_13_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__7_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__7_LC_13_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__7_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12154),
            .lcout(\c0.d_4_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19602),
            .ce(N__17174),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__3_LC_13_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__3_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__3_LC_13_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__3_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12138),
            .lcout(\c0.d_4_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19602),
            .ce(N__17174),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIO7RC_40_LC_13_18_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIO7RC_40_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIO7RC_40_LC_13_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIO7RC_40_LC_13_18_0  (
            .in0(N__16183),
            .in1(N__17984),
            .in2(N__17221),
            .in3(N__18174),
            .lcout(),
            .ltout(\c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI240O_40_LC_13_18_1 .C_ON=1'b0;
    defparam \c0.d_4_RNI240O_40_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI240O_40_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.d_4_RNI240O_40_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__12251),
            .in2(N__12361),
            .in3(N__13797),
            .lcout(\c0.un1_data_in_6__6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__4_LC_13_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__4_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__4_LC_13_18_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_frame_3__4_LC_13_18_2  (
            .in0(N__12358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19615),
            .ce(N__17178),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI1VL6_13_LC_13_18_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI1VL6_13_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI1VL6_13_LC_13_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNI1VL6_13_LC_13_18_3  (
            .in0(N__17922),
            .in1(N__16039),
            .in2(_gnd_net_),
            .in3(N__15962),
            .lcout(\c0.N_132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__5_LC_13_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__5_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__5_LC_13_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__5_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12331),
            .lcout(\c0.d_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19615),
            .ce(N__17178),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__2_LC_13_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__2_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__2_LC_13_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__2_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12310),
            .lcout(\c0.d_4_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19615),
            .ce(N__17178),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__1_LC_13_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__1_LC_13_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__1_LC_13_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__1_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12292),
            .lcout(\c0.d_4_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19615),
            .ce(N__17178),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__0_LC_13_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__0_LC_13_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__0_LC_13_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__0_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12277),
            .lcout(\c0.d_4_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19615),
            .ce(N__17178),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI1LAI2_12_LC_13_19_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI1LAI2_12_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI1LAI2_12_LC_13_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI1LAI2_12_LC_13_19_0  (
            .in0(N__16302),
            .in1(N__12258),
            .in2(N__12400),
            .in3(N__16161),
            .lcout(),
            .ltout(\c0.un1_data_in_7__0_0_a2_1_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI20TA7_15_LC_13_19_1 .C_ON=1'b0;
    defparam \c0.d_4_RNI20TA7_15_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI20TA7_15_LC_13_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI20TA7_15_LC_13_19_1  (
            .in0(N__16505),
            .in1(N__16544),
            .in2(N__12433),
            .in3(N__12409),
            .lcout(\c0.un1_data_in_7__0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIJ66B_11_LC_13_19_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIJ66B_11_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIJ66B_11_LC_13_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIJ66B_11_LC_13_19_2  (
            .in0(N__18818),
            .in1(N__14579),
            .in2(N__16438),
            .in3(N__13883),
            .lcout(\c0.N_121 ),
            .ltout(\c0.N_121_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNITCL32_11_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.d_4_RNITCL32_11_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNITCL32_11_LC_13_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.d_4_RNITCL32_11_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__13833),
            .in2(N__12430),
            .in3(N__12427),
            .lcout(),
            .ltout(\c0.un1_data_in_6__7_0_a2_17_a2_4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIV4MJ3_10_LC_13_19_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIV4MJ3_10_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIV4MJ3_10_LC_13_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIV4MJ3_10_LC_13_19_4  (
            .in0(N__15892),
            .in1(N__12445),
            .in2(N__12412),
            .in3(N__16404),
            .lcout(\c0.N_136 ),
            .ltout(\c0.N_136_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIK2SL3_14_LC_13_19_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIK2SL3_14_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIK2SL3_14_LC_13_19_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.d_4_RNIK2SL3_14_LC_13_19_5  (
            .in0(N__16272),
            .in1(_gnd_net_),
            .in2(N__12403),
            .in3(_gnd_net_),
            .lcout(\c0.un1_data_in_7__1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIG6H4_39_LC_13_19_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIG6H4_39_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIG6H4_39_LC_13_19_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.d_4_RNIG6H4_39_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__17465),
            .in2(_gnd_net_),
            .in3(N__18173),
            .lcout(\c0.N_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIH0UG_12_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIH0UG_12_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIH0UG_12_LC_13_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIH0UG_12_LC_13_20_0  (
            .in0(N__14667),
            .in1(N__16184),
            .in2(N__17370),
            .in3(N__18036),
            .lcout(\c0.un1_data_in_7__0_0_a2_1_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__3_LC_13_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__3_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__3_LC_13_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__3_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12387),
            .lcout(\c0.d_4_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19627),
            .ce(N__17183),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIQ3V8_12_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIQ3V8_12_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIQ3V8_12_LC_13_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIQ3V8_12_LC_13_20_2  (
            .in0(N__14666),
            .in1(N__16328),
            .in2(N__13934),
            .in3(N__18035),
            .lcout(),
            .ltout(\c0.un1_data_in_7__1_0_a2_24_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIQ7KN_16_LC_13_20_3 .C_ON=1'b0;
    defparam \c0.d_4_RNIQ7KN_16_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIQ7KN_16_LC_13_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIQ7KN_16_LC_13_20_3  (
            .in0(N__17993),
            .in1(N__17333),
            .in2(N__12553),
            .in3(N__18849),
            .lcout(\c0.un1_data_in_7__1_0_a2_24_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__4_LC_13_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__4_LC_13_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__4_LC_13_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__4_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12544),
            .lcout(\c0.d_4_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19627),
            .ce(N__17183),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__2_LC_13_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__2_LC_13_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__2_LC_13_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__2_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12526),
            .lcout(\c0.d_4_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19627),
            .ce(N__17183),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__0_LC_13_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__0_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__0_LC_13_20_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_frame_2__0_LC_13_20_6  (
            .in0(N__12508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19627),
            .ce(N__17183),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIA0HJ_0_LC_13_20_7 .C_ON=1'b0;
    defparam \c0.d_4_RNIA0HJ_0_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIA0HJ_0_LC_13_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNIA0HJ_0_LC_13_20_7  (
            .in0(N__18094),
            .in1(N__18894),
            .in2(_gnd_net_),
            .in3(N__18848),
            .lcout(\c0.N_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI34PL_16_LC_13_21_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI34PL_16_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI34PL_16_LC_13_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI34PL_16_LC_13_21_0  (
            .in0(N__18096),
            .in1(N__18847),
            .in2(N__12481),
            .in3(N__14611),
            .lcout(),
            .ltout(\c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI6DG41_18_LC_13_21_1 .C_ON=1'b0;
    defparam \c0.d_4_RNI6DG41_18_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI6DG41_18_LC_13_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI6DG41_18_LC_13_21_1  (
            .in0(N__12657),
            .in1(N__15750),
            .in2(N__12448),
            .in3(N__13935),
            .lcout(\c0.un1_data_in_7__4_0_a2_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIABPL_18_LC_13_21_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIABPL_18_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIABPL_18_LC_13_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIABPL_18_LC_13_21_2  (
            .in0(N__17964),
            .in1(N__12656),
            .in2(N__16371),
            .in3(N__17900),
            .lcout(\c0.N_124 ),
            .ltout(\c0.N_124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__RNIBJH41_6_LC_13_21_3 .C_ON=1'b0;
    defparam \c0.data_in_7__RNIBJH41_6_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_7__RNIBJH41_6_LC_13_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_7__RNIBJH41_6_LC_13_21_3  (
            .in0(N__17251),
            .in1(N__18401),
            .in2(N__12436),
            .in3(N__14709),
            .lcout(),
            .ltout(\c0.un1_data_in_7__6_0_a2_5_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIDD8G3_18_LC_13_21_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIDD8G3_18_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIDD8G3_18_LC_13_21_4 .LUT_INIT=16'b0001001001001000;
    LogicCell40 \c0.d_4_RNIDD8G3_18_LC_13_21_4  (
            .in0(N__12745),
            .in1(N__13942),
            .in2(N__12727),
            .in3(N__12724),
            .lcout(\c0.m163_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__3_LC_13_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__3_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__3_LC_13_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__3_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12718),
            .lcout(\c0.d_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19635),
            .ce(N__17186),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__5_LC_13_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__5_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__5_LC_13_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__5_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12700),
            .lcout(\c0.d_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19635),
            .ce(N__17186),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_7_LC_13_22_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_7_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_7_LC_13_22_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \c0.tx2_data_RNO_2_7_LC_13_22_0  (
            .in0(N__13675),
            .in1(N__18714),
            .in2(N__14374),
            .in3(N__18797),
            .lcout(\c0.m60_0_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_2_LC_13_22_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_2_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_2_LC_13_22_1 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx2_data_RNO_4_2_LC_13_22_1  (
            .in0(N__18576),
            .in1(N__16050),
            .in2(N__12661),
            .in3(N__18354),
            .lcout(\c0.tx2_data_RNO_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__2_LC_13_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__2_LC_13_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__2_LC_13_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__2_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12682),
            .lcout(\c0.d_4_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19642),
            .ce(N__17188),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_6_LC_13_23_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_6_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_6_LC_13_23_1 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx_data_RNO_4_6_LC_13_23_1  (
            .in0(N__15533),
            .in1(N__14983),
            .in2(N__14464),
            .in3(N__15365),
            .lcout(\c0.tx_data_RNO_4Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_6_LC_13_23_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_6_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_6_LC_13_23_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx_data_RNO_0_6_LC_13_23_2  (
            .in0(N__15368),
            .in1(N__12643),
            .in2(N__12613),
            .in3(N__15537),
            .lcout(\c0.tx_data_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_7_LC_13_23_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_7_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_7_LC_13_23_3 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_1_7_LC_13_23_3  (
            .in0(N__15536),
            .in1(N__12586),
            .in2(N__12574),
            .in3(N__15369),
            .lcout(\c0.tx_data_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_5_LC_13_23_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_5_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_5_LC_13_23_4 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \c0.tx_data_RNO_0_5_LC_13_23_4  (
            .in0(N__15367),
            .in1(N__15535),
            .in2(N__13021),
            .in3(N__12985),
            .lcout(\c0.tx_data_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_6_LC_13_23_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_6_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_6_LC_13_23_6 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx_data_RNO_3_6_LC_13_23_6  (
            .in0(N__15366),
            .in1(N__14502),
            .in2(N__15026),
            .in3(N__15534),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_6_LC_13_23_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_6_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_6_LC_13_23_7 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_6_LC_13_23_7  (
            .in0(N__15165),
            .in1(N__15651),
            .in2(N__12955),
            .in3(N__12952),
            .lcout(\c0.tx_data_1_0_i_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIK3C71_13_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.d_2_RNIK3C71_13_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIK3C71_13_LC_13_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIK3C71_13_LC_13_24_0  (
            .in0(N__14775),
            .in1(N__12827),
            .in2(N__12946),
            .in3(N__12767),
            .lcout(\c0.nextCRC16_3_3_1 ),
            .ltout(\c0.nextCRC16_3_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_1_LC_13_24_1 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_1_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_1_LC_13_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_0_1_LC_13_24_1  (
            .in0(N__12880),
            .in1(N__13054),
            .in2(N__12853),
            .in3(N__14926),
            .lcout(\c0.nextCRC16_3_0_a2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__5_LC_13_24_2 .C_ON=1'b0;
    defparam \c0.data_out_1__5_LC_13_24_2 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__5_LC_13_24_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_out_1__5_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__17006),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19656),
            .ce(),
            .sr(N__16878));
    defparam \c0.data_out_3__4_LC_13_24_3 .C_ON=1'b0;
    defparam \c0.data_out_3__4_LC_13_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__4_LC_13_24_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_3__4_LC_13_24_3  (
            .in0(N__17007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19656),
            .ce(),
            .sr(N__16878));
    defparam \c0.tx_data_RNO_3_5_LC_13_24_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_5_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_5_LC_13_24_5 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_3_5_LC_13_24_5  (
            .in0(N__12810),
            .in1(N__15556),
            .in2(N__12774),
            .in3(N__15339),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_5_LC_13_24_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_5_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_5_LC_13_24_6 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_5_LC_13_24_6  (
            .in0(N__15163),
            .in1(N__15640),
            .in2(N__12754),
            .in3(N__13204),
            .lcout(\c0.tx_data_1_0_i_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_5_LC_13_24_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_5_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_5_LC_13_24_7 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \c0.tx_data_RNO_4_5_LC_13_24_7  (
            .in0(N__16909),
            .in1(N__15555),
            .in2(N__14866),
            .in3(N__15338),
            .lcout(\c0.tx_data_RNO_4Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_0_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_0_LC_13_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_0_LC_13_25_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \c0.tx.r_Tx_Data_0_LC_13_25_0  (
            .in0(N__13198),
            .in1(N__13186),
            .in2(N__15209),
            .in3(N__13180),
            .lcout(\c0.tx.r_Tx_DataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19664),
            .ce(N__14283),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_2_LC_13_25_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_2_LC_13_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_2_LC_13_25_2 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \c0.tx.r_Tx_Data_2_LC_13_25_2  (
            .in0(N__13060),
            .in1(N__13162),
            .in2(N__15210),
            .in3(N__13414),
            .lcout(\c0.tx.r_Tx_DataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19664),
            .ce(N__14283),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_1_LC_13_25_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_1_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_1_LC_13_25_4 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_4_1_LC_13_25_4  (
            .in0(N__14933),
            .in1(N__15517),
            .in2(N__13144),
            .in3(N__15364),
            .lcout(),
            .ltout(\c0.tx_data_RNO_4Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_1_LC_13_25_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_1_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_1_LC_13_25_5 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \c0.tx_data_RNO_2_1_LC_13_25_5  (
            .in0(N__15650),
            .in1(N__15187),
            .in2(N__13108),
            .in3(N__13459),
            .lcout(),
            .ltout(\c0.tx_data_1_0_i_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_1_LC_13_25_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_1_LC_13_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_1_LC_13_25_6 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \c0.tx.r_Tx_Data_1_LC_13_25_6  (
            .in0(N__13105),
            .in1(N__15164),
            .in2(N__13099),
            .in3(N__13246),
            .lcout(\c0.tx.r_Tx_DataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19664),
            .ce(N__14283),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_2_LC_13_26_0 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_2_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_2_LC_13_26_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx_data_RNO_1_2_LC_13_26_0  (
            .in0(N__15289),
            .in1(N__13084),
            .in2(N__15539),
            .in3(N__13072),
            .lcout(\c0.tx_data_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_2_LC_13_26_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_2_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_2_LC_13_26_1 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \c0.tx_data_RNO_4_2_LC_13_26_1  (
            .in0(N__14776),
            .in1(N__15500),
            .in2(N__14743),
            .in3(N__15284),
            .lcout(\c0.tx_data_RNO_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_1_LC_13_26_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_1_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_1_LC_13_26_2 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \c0.tx_data_RNO_3_1_LC_13_26_2  (
            .in0(N__15286),
            .in1(N__13050),
            .in2(N__15538),
            .in3(N__13484),
            .lcout(\c0.tx_data_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_2_LC_13_26_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_2_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_2_LC_13_26_3 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \c0.tx_data_RNO_3_2_LC_13_26_3  (
            .in0(N__15704),
            .in1(N__15503),
            .in2(N__13453),
            .in3(N__15285),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_2_LC_13_26_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_2_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_2_LC_13_26_4 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_2_LC_13_26_4  (
            .in0(N__15167),
            .in1(N__15631),
            .in2(N__13423),
            .in3(N__13420),
            .lcout(\c0.tx_data_1_0_i_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_7_LC_13_26_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_7_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_7_LC_13_26_5 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_0_7_LC_13_26_5  (
            .in0(N__13408),
            .in1(N__15502),
            .in2(N__13366),
            .in3(N__15288),
            .lcout(\c0.tx_data_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_4_LC_13_26_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_4_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_4_LC_13_26_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_0_4_LC_13_26_7  (
            .in0(N__13330),
            .in1(N__15501),
            .in2(N__13303),
            .in3(N__15287),
            .lcout(\c0.tx_data_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_1_LC_13_27_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_1_LC_13_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_1_LC_13_27_3 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_1_1_LC_13_27_3  (
            .in0(N__15473),
            .in1(N__13270),
            .in2(N__13261),
            .in3(N__15333),
            .lcout(\c0.tx_data_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNI7Q6P_6_LC_13_27_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNI7Q6P_6_LC_13_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNI7Q6P_6_LC_13_27_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \c0.byte_transmit_counter_RNI7Q6P_6_LC_13_27_4  (
            .in0(_gnd_net_),
            .in1(N__15676),
            .in2(_gnd_net_),
            .in3(N__15682),
            .lcout(),
            .ltout(\c0.m2_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNIQP0V1_3_LC_13_27_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNIQP0V1_3_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNIQP0V1_3_LC_13_27_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.byte_transmit_counter_RNIQP0V1_3_LC_13_27_5  (
            .in0(N__13594),
            .in1(N__15664),
            .in2(N__13237),
            .in3(N__15670),
            .lcout(\c0.N_132_mux ),
            .ltout(\c0.N_132_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_3_LC_13_27_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_3_LC_13_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_3_LC_13_27_6 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \c0.tx_data_RNO_1_3_LC_13_27_6  (
            .in0(N__13234),
            .in1(N__13228),
            .in2(N__13219),
            .in3(N__15472),
            .lcout(\c0.tx_data_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5_LC_13_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5_LC_13_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_5_LC_13_28_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_5_LC_13_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19676),
            .ce(N__15075),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0_LC_13_28_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0_LC_13_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_0_LC_13_28_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.byte_transmit_counter_0_LC_13_28_5  (
            .in0(_gnd_net_),
            .in1(N__15474),
            .in2(_gnd_net_),
            .in3(N__15335),
            .lcout(\c0.byte_transmit_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19676),
            .ce(N__15075),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_2_LC_13_28_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_2_LC_13_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_2_LC_13_28_6 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \c0.byte_transmit_counter_2_LC_13_28_6  (
            .in0(N__15336),
            .in1(N__15133),
            .in2(N__15528),
            .in3(N__15633),
            .lcout(\c0.byte_transmit_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19676),
            .ce(N__15075),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__4_LC_14_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__4_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__4_LC_14_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__4_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15746),
            .lcout(\c0.data_in_frame_7_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19619),
            .ce(N__17172),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_7_LC_14_17_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_7_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_7_LC_14_17_0 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.tx2_data_RNO_1_7_LC_14_17_0  (
            .in0(N__13558),
            .in1(N__18347),
            .in2(N__13522),
            .in3(N__18590),
            .lcout(\c0.tx2_data_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__7_LC_14_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__7_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__7_LC_14_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__7_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13588),
            .lcout(\c0.data_in_frame_6_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19610),
            .ce(N__17173),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__7_LC_14_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__7_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__7_LC_14_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__7_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13548),
            .lcout(\c0.data_in_frame_7_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19610),
            .ce(N__17173),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_6_LC_14_17_3 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_6_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_6_LC_14_17_3 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \c0.tx2_data_RNO_3_6_LC_14_17_3  (
            .in0(N__18591),
            .in1(N__16268),
            .in2(N__18372),
            .in3(N__13749),
            .lcout(\c0.tx2_data_RNO_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__6_LC_14_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__6_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__6_LC_14_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__6_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13513),
            .lcout(\c0.d_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19610),
            .ce(N__17173),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIUBBH_6_LC_14_17_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIUBBH_6_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIUBBH_6_LC_14_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.d_4_RNIUBBH_6_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__13748),
            .in2(_gnd_net_),
            .in3(N__14704),
            .lcout(\c0.N_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__6_LC_14_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__6_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__6_LC_14_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__6_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13723),
            .lcout(\c0.d_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19610),
            .ce(N__17173),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_7_LC_14_17_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_7_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_7_LC_14_17_7 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \c0.tx2_data_RNO_3_7_LC_14_17_7  (
            .in0(N__18589),
            .in1(N__16516),
            .in2(N__18371),
            .in3(N__13696),
            .lcout(\c0.tx2_data_RNO_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__4_LC_14_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__4_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__4_LC_14_18_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_in_frame_4__4_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__13659),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19620),
            .ce(N__17175),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIJ8G4_36_LC_14_18_1 .C_ON=1'b0;
    defparam \c0.d_4_RNIJ8G4_36_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIJ8G4_36_LC_14_18_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.d_4_RNIJ8G4_36_LC_14_18_1  (
            .in0(N__13901),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17648),
            .lcout(),
            .ltout(\c0.N_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__RNIKD2F_1_LC_14_18_2 .C_ON=1'b0;
    defparam \c0.data_in_6__RNIKD2F_1_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_6__RNIKD2F_1_LC_14_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_6__RNIKD2F_1_LC_14_18_2  (
            .in0(N__13642),
            .in1(N__16435),
            .in2(N__13621),
            .in3(N__14705),
            .lcout(\c0.un1_data_in_6__1_0_a2_4_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI76N6_22_LC_14_18_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI76N6_22_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI76N6_22_LC_14_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNI76N6_22_LC_14_18_3  (
            .in0(N__13900),
            .in1(N__17647),
            .in2(_gnd_net_),
            .in3(N__18117),
            .lcout(\c0.N_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__6_LC_14_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__6_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__6_LC_14_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__6_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13618),
            .lcout(\c0.d_4_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19620),
            .ce(N__17175),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__6_LC_14_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__6_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__6_LC_14_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__6_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16098),
            .lcout(\c0.d_4_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19620),
            .ce(N__17175),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_4_LC_14_18_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_4_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_4_LC_14_18_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \c0.tx2_data_RNO_0_4_LC_14_18_6  (
            .in0(N__18588),
            .in1(N__13936),
            .in2(N__18375),
            .in3(N__13902),
            .lcout(\c0.tx2_data_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_6_LC_14_18_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_6_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_6_LC_14_18_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx2_data_RNO_0_6_LC_14_18_7  (
            .in0(N__16436),
            .in1(N__18587),
            .in2(N__16372),
            .in3(N__18365),
            .lcout(\c0.tx2_data_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI23VN_11_LC_14_19_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI23VN_11_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI23VN_11_LC_14_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI23VN_11_LC_14_19_0  (
            .in0(N__13793),
            .in1(N__14586),
            .in2(N__13810),
            .in3(N__13884),
            .lcout(),
            .ltout(\c0.un1_data_in_6__5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNITNPS1_11_LC_14_19_1 .C_ON=1'b0;
    defparam \c0.d_4_RNITNPS1_11_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNITNPS1_11_LC_14_19_1 .LUT_INIT=16'b0000011000001001;
    LogicCell40 \c0.d_4_RNITNPS1_11_LC_14_19_1  (
            .in0(N__13885),
            .in1(N__13870),
            .in2(N__13858),
            .in3(N__15891),
            .lcout(),
            .ltout(\c0.m163_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__RNIAQG64_1_LC_14_19_2 .C_ON=1'b0;
    defparam \c0.data_in_6__RNIAQG64_1_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_6__RNIAQG64_1_LC_14_19_2 .LUT_INIT=16'b0100000000010000;
    LogicCell40 \c0.data_in_6__RNIAQG64_1_LC_14_19_2  (
            .in0(N__13855),
            .in1(N__13849),
            .in2(N__13843),
            .in3(N__13840),
            .lcout(),
            .ltout(\c0.m163_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIFGESA_24_LC_14_19_3 .C_ON=1'b0;
    defparam \c0.d_4_RNIFGESA_24_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIFGESA_24_LC_14_19_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.d_4_RNIFGESA_24_LC_14_19_3  (
            .in0(N__16282),
            .in1(N__16381),
            .in2(N__13822),
            .in3(N__13819),
            .lcout(\c0.m163_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIN4PC_25_LC_14_19_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIN4PC_25_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIN4PC_25_LC_14_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIN4PC_25_LC_14_19_4  (
            .in0(N__17291),
            .in1(N__14665),
            .in2(N__15980),
            .in3(N__15818),
            .lcout(\c0.un1_data_in_6__5_0_a2_5_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI9TE4_12_LC_14_19_5 .C_ON=1'b0;
    defparam \c0.d_4_RNI9TE4_12_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI9TE4_12_LC_14_19_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.d_4_RNI9TE4_12_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__16327),
            .in2(_gnd_net_),
            .in3(N__18034),
            .lcout(\c0.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__4_LC_14_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__4_LC_14_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__4_LC_14_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__4_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13777),
            .lcout(\c0.d_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19628),
            .ce(N__17179),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIC7M21_1_LC_14_20_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIC7M21_1_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIC7M21_1_LC_14_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIC7M21_1_LC_14_20_0  (
            .in0(N__18402),
            .in1(N__16245),
            .in2(N__16675),
            .in3(N__14365),
            .lcout(\c0.N_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_7_c_RNIGB9N4_LC_14_20_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNIGB9N4_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNIGB9N4_LC_14_20_1 .LUT_INIT=16'b1000010000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_RNIGB9N4_LC_14_20_1  (
            .in0(N__14032),
            .in1(N__14026),
            .in2(N__15946),
            .in3(N__19287),
            .lcout(),
            .ltout(\c0.m163_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIGIT3F_14_LC_14_20_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIGIT3F_14_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIGIT3F_14_LC_14_20_2 .LUT_INIT=16'b0111111111101111;
    LogicCell40 \c0.d_4_RNIGIT3F_14_LC_14_20_2  (
            .in0(N__14020),
            .in1(N__14011),
            .in2(N__14002),
            .in3(N__13999),
            .lcout(),
            .ltout(\c0.m163_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI7JOT41_15_LC_14_20_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI7JOT41_15_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI7JOT41_15_LC_14_20_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.d_4_RNI7JOT41_15_LC_14_20_3  (
            .in0(N__13993),
            .in1(N__16132),
            .in2(N__13987),
            .in3(N__13984),
            .lcout(\c0.N_164_0 ),
            .ltout(\c0.N_164_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_RNIG45P61_LC_14_20_4 .C_ON=1'b0;
    defparam \c0.tx2_transmit_RNIG45P61_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_transmit_RNIG45P61_LC_14_20_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.tx2_transmit_RNIG45P61_LC_14_20_4  (
            .in0(N__19339),
            .in1(N__20013),
            .in2(N__13978),
            .in3(N__17809),
            .lcout(\c0.N_173_0 ),
            .ltout(\c0.N_173_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_active_RNIABU671_LC_14_20_5 .C_ON=1'b0;
    defparam \c0.tx2_active_RNIABU671_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_active_RNIABU671_LC_14_20_5 .LUT_INIT=16'b0011000000110000;
    LogicCell40 \c0.tx2_active_RNIABU671_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__19721),
            .in2(N__13975),
            .in3(_gnd_net_),
            .lcout(\c0.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIM5UG_19_LC_14_21_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIM5UG_19_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIM5UG_19_LC_14_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIM5UG_19_LC_14_21_0  (
            .in0(N__18400),
            .in1(N__16243),
            .in2(N__17275),
            .in3(N__14640),
            .lcout(\c0.un1_data_in_7__5_0_a2_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__7_LC_14_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__7_LC_14_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__7_LC_14_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__7_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13972),
            .lcout(\c0.d_4_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19643),
            .ce(N__17184),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIB3JJ_2_LC_14_21_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIB3JJ_2_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIB3JJ_2_LC_14_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNIB3JJ_2_LC_14_21_2  (
            .in0(N__18399),
            .in1(N__16242),
            .in2(_gnd_net_),
            .in3(N__14360),
            .lcout(\c0.d_4_RNIB3JJZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__2_LC_14_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__2_LC_14_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__2_LC_14_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__2_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14437),
            .lcout(\c0.d_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19643),
            .ce(N__17184),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__0_LC_14_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__0_LC_14_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__0_LC_14_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__0_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14419),
            .lcout(\c0.d_4_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19643),
            .ce(N__17184),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_7_LC_14_21_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_7_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_7_LC_14_21_5 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \c0.tx2_data_RNO_4_7_LC_14_21_5  (
            .in0(N__16244),
            .in1(N__18305),
            .in2(N__18570),
            .in3(N__14398),
            .lcout(\c0.tx2_data_RNO_4Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_2_LC_14_21_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_2_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_2_LC_14_21_6 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \c0.tx2_data_RNO_3_2_LC_14_21_6  (
            .in0(N__15910),
            .in1(N__18514),
            .in2(N__18353),
            .in3(N__14361),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_2_LC_14_21_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_2_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_2_LC_14_21_7 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \c0.tx2_data_RNO_2_2_LC_14_21_7  (
            .in0(N__18657),
            .in1(N__14347),
            .in2(N__14338),
            .in3(N__18784),
            .lcout(\c0.m131_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_6_LC_14_22_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_6_LC_14_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_6_LC_14_22_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \c0.tx.r_Tx_Data_6_LC_14_22_0  (
            .in0(N__14323),
            .in1(N__14311),
            .in2(N__15211),
            .in3(N__14305),
            .lcout(\c0.tx.r_Tx_DataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19650),
            .ce(N__14287),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNIC9J951_LC_14_22_2 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNIC9J951_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNIC9J951_LC_14_22_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.wait_for_transmission_RNIC9J951_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(N__19342),
            .in2(_gnd_net_),
            .in3(N__18142),
            .lcout(\c0.tx2_transmit_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_RNIRD3K_1_LC_14_22_5 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_RNIRD3K_1_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Bit_Index_RNIRD3K_1_LC_14_22_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \c0.rx.r_Bit_Index_RNIRD3K_1_LC_14_22_5  (
            .in0(N__14247),
            .in1(N__14185),
            .in2(_gnd_net_),
            .in3(N__14124),
            .lcout(\c0.rx.N_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_3_LC_14_23_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_3_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_3_LC_14_23_0 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \c0.tx2_data_RNO_0_3_LC_14_23_0  (
            .in0(N__16198),
            .in1(N__18357),
            .in2(N__18595),
            .in3(N__14713),
            .lcout(\c0.tx2_data_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_3_LC_14_23_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_3_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_3_LC_14_23_1 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \c0.tx2_data_RNO_4_3_LC_14_23_1  (
            .in0(N__18355),
            .in1(N__14674),
            .in2(N__14647),
            .in3(N__18582),
            .lcout(\c0.tx2_data_RNO_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_3_LC_14_23_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_3_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_3_LC_14_23_2 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx2_data_RNO_3_3_LC_14_23_2  (
            .in0(N__18586),
            .in1(N__14617),
            .in2(N__14593),
            .in3(N__18356),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_3_LC_14_23_3 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_3_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_3_LC_14_23_3 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \c0.tx2_data_RNO_2_3_LC_14_23_3  (
            .in0(N__18798),
            .in1(N__14566),
            .in2(N__14560),
            .in3(N__18719),
            .lcout(),
            .ltout(\c0.m105_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_3_LC_14_23_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_3_LC_14_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_3_LC_14_23_4 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \c0.tx2.r_Tx_Data_3_LC_14_23_4  (
            .in0(N__14557),
            .in1(N__18721),
            .in2(N__14551),
            .in3(N__14548),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19657),
            .ce(N__19973),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_3_LC_14_23_5 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_3_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_3_LC_14_23_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_3_LC_14_23_5  (
            .in0(N__14509),
            .in1(N__14536),
            .in2(_gnd_net_),
            .in3(N__19822),
            .lcout(\c0.tx2.o_Tx_Serial_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_7_LC_14_23_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_7_LC_14_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_7_LC_14_23_6 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \c0.tx2.r_Tx_Data_7_LC_14_23_6  (
            .in0(N__18720),
            .in1(N__17452),
            .in2(N__14530),
            .in3(N__14515),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19657),
            .ce(N__19973),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__6_LC_14_24_1 .C_ON=1'b0;
    defparam \c0.data_out_0__6_LC_14_24_1 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__6_LC_14_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__6_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17008),
            .lcout(\c0.d_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19665),
            .ce(),
            .sr(N__16875));
    defparam \c0.data_out_2__6_LC_14_24_5 .C_ON=1'b0;
    defparam \c0.data_out_2__6_LC_14_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__6_LC_14_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__6_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17010),
            .lcout(\c0.d_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19665),
            .ce(),
            .sr(N__16875));
    defparam \c0.data_out_1__6_LC_14_24_6 .C_ON=1'b0;
    defparam \c0.data_out_1__6_LC_14_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__6_LC_14_24_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_1__6_LC_14_24_6  (
            .in0(N__17009),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19665),
            .ce(),
            .sr(N__16875));
    defparam \c0.data_out_3__6_LC_14_24_7 .C_ON=1'b0;
    defparam \c0.data_out_3__6_LC_14_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__6_LC_14_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__6_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17011),
            .lcout(\c0.d_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19665),
            .ce(),
            .sr(N__16875));
    defparam \c0.data_out_2__0_LC_14_25_0 .C_ON=1'b0;
    defparam \c0.data_out_2__0_LC_14_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__0_LC_14_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__0_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17087),
            .lcout(\c0.d_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19670),
            .ce(),
            .sr(N__16874));
    defparam \c0.data_out_2__1_LC_14_25_1 .C_ON=1'b0;
    defparam \c0.data_out_2__1_LC_14_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__1_LC_14_25_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_2__1_LC_14_25_1  (
            .in0(N__17088),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19670),
            .ce(),
            .sr(N__16874));
    defparam \c0.data_out_1__4_LC_14_25_2 .C_ON=1'b0;
    defparam \c0.data_out_1__4_LC_14_25_2 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__4_LC_14_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_1__4_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17086),
            .lcout(\c0.d_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19670),
            .ce(),
            .sr(N__16874));
    defparam \c0.data_out_2__5_LC_14_25_3 .C_ON=1'b0;
    defparam \c0.data_out_2__5_LC_14_25_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__5_LC_14_25_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_2__5_LC_14_25_3  (
            .in0(N__17090),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19670),
            .ce(),
            .sr(N__16874));
    defparam \c0.data_out_1__3_LC_14_25_4 .C_ON=1'b0;
    defparam \c0.data_out_1__3_LC_14_25_4 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__3_LC_14_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_1__3_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17085),
            .lcout(\c0.d_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19670),
            .ce(),
            .sr(N__16874));
    defparam \c0.data_out_3__2_LC_14_25_5 .C_ON=1'b0;
    defparam \c0.data_out_3__2_LC_14_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__2_LC_14_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__2_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.d_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19670),
            .ce(),
            .sr(N__16874));
    defparam \c0.data_out_2__2_LC_14_25_6 .C_ON=1'b0;
    defparam \c0.data_out_2__2_LC_14_25_6 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__2_LC_14_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__2_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17089),
            .lcout(\c0.d_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19670),
            .ce(),
            .sr(N__16874));
    defparam \c0.data_out_1__2_LC_14_26_1 .C_ON=1'b0;
    defparam \c0.data_out_1__2_LC_14_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__2_LC_14_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_1__2_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17091),
            .lcout(\c0.d_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19673),
            .ce(),
            .sr(N__16872));
    defparam \c0.byte_transmit_counter_1_LC_14_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1_LC_14_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1_LC_14_27_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \c0.byte_transmit_counter_1_LC_14_27_0  (
            .in0(N__15632),
            .in1(N__15478),
            .in2(_gnd_net_),
            .in3(N__15337),
            .lcout(\c0.byte_transmit_counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19677),
            .ce(N__15079),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_6_LC_14_27_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_6_LC_14_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_6_LC_14_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_6_LC_14_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19677),
            .ce(N__15079),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_7_LC_14_27_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_7_LC_14_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_7_LC_14_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_7_LC_14_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19677),
            .ce(N__15079),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_3_LC_14_27_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_3_LC_14_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_3_LC_14_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_3_LC_14_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19677),
            .ce(N__15079),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4_LC_14_27_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4_LC_14_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_4_LC_14_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_4_LC_14_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19677),
            .ce(N__15079),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNIL77O2_1_LC_14_28_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNIL77O2_1_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNIL77O2_1_LC_14_28_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \c0.byte_transmit_counter_RNIL77O2_1_LC_14_28_2  (
            .in0(N__15610),
            .in1(N__15429),
            .in2(_gnd_net_),
            .in3(N__15282),
            .lcout(),
            .ltout(\c0.N_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNI4QES5_2_LC_14_28_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNI4QES5_2_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNI4QES5_2_LC_14_28_3 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \c0.byte_transmit_counter_RNI4QES5_2_LC_14_28_3  (
            .in0(N__15283),
            .in1(N__15110),
            .in2(N__15082),
            .in3(N__15063),
            .lcout(\c0.data_out_0__1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__4_LC_15_16_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__4_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__4_LC_15_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__4_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16011),
            .lcout(\c0.data_in_frame_6_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19629),
            .ce(N__17170),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_4_LC_15_17_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_4_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_4_LC_15_17_0 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \c0.tx2_data_RNO_1_4_LC_15_17_0  (
            .in0(N__15802),
            .in1(N__18348),
            .in2(N__18593),
            .in3(N__15796),
            .lcout(\c0.tx2_data_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_4_LC_15_17_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_4_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_4_LC_15_17_2 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \c0.tx2_data_RNO_2_4_LC_15_17_2  (
            .in0(N__18709),
            .in1(N__17941),
            .in2(N__18016),
            .in3(N__18795),
            .lcout(),
            .ltout(\c0.m120_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_4_LC_15_17_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_4_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_4_LC_15_17_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \c0.tx2.r_Tx_Data_4_LC_15_17_3  (
            .in0(N__15790),
            .in1(N__15784),
            .in2(N__15778),
            .in3(N__18711),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19617),
            .ce(N__19977),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_6_LC_15_17_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_6_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_6_LC_15_17_5 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \c0.tx2_data_RNO_2_6_LC_15_17_5  (
            .in0(N__18796),
            .in1(N__15775),
            .in2(N__18073),
            .in3(N__18710),
            .lcout(),
            .ltout(\c0.m90_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_6_LC_15_17_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_6_LC_15_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_6_LC_15_17_6 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \c0.tx2.r_Tx_Data_6_LC_15_17_6  (
            .in0(N__15769),
            .in1(N__18718),
            .in2(N__15763),
            .in3(N__15760),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19617),
            .ce(N__19977),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_6_LC_15_17_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_6_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_6_LC_15_17_7 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \c0.tx2_data_RNO_1_6_LC_15_17_7  (
            .in0(N__18592),
            .in1(N__17227),
            .in2(N__18373),
            .in3(N__17197),
            .lcout(\c0.tx2_data_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__4_LC_15_18_1 .C_ON=1'b0;
    defparam \c0.data_in_6__4_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__4_LC_15_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__4_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15754),
            .lcout(\c0.data_in_6_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19630),
            .ce(N__17726),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__5_LC_15_18_2 .C_ON=1'b0;
    defparam \c0.data_in_6__5_LC_15_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__5_LC_15_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__5_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17270),
            .lcout(\c0.data_in_6_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19630),
            .ce(N__17726),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__5_LC_15_18_3 .C_ON=1'b0;
    defparam \c0.data_in_7__5_LC_15_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__5_LC_15_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__5_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15727),
            .lcout(\c0.data_in_7_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19630),
            .ce(N__17726),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__6_LC_15_18_4 .C_ON=1'b0;
    defparam \c0.data_in_4__6_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__6_LC_15_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__6_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16080),
            .lcout(\c0.data_in_4_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19630),
            .ce(N__17726),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__6_LC_15_18_5 .C_ON=1'b0;
    defparam \c0.data_in_5__6_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__6_LC_15_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__6_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17216),
            .lcout(\c0.data_in_5_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19630),
            .ce(N__17726),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__6_LC_15_18_6 .C_ON=1'b0;
    defparam \c0.data_in_6__6_LC_15_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__6_LC_15_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__6_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17246),
            .lcout(\c0.data_in_6_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19630),
            .ce(N__17726),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__6_LC_15_18_7 .C_ON=1'b0;
    defparam \c0.data_in_7__6_LC_15_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__6_LC_15_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__6_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16069),
            .lcout(\c0.data_in_7_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19630),
            .ce(N__17726),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIFRNC_10_LC_15_19_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIFRNC_10_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIFRNC_10_LC_15_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIFRNC_10_LC_15_19_0  (
            .in0(N__15906),
            .in1(N__16051),
            .in2(N__16010),
            .in3(N__15981),
            .lcout(\c0.un1_data_in_6__4_0_a2_5_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__2_LC_15_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__2_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__2_LC_15_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__2_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15937),
            .lcout(\c0.d_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19636),
            .ce(N__17176),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIH6GJ_10_LC_15_19_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIH6GJ_10_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIH6GJ_10_LC_15_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNIH6GJ_10_LC_15_19_2  (
            .in0(N__15905),
            .in1(N__16646),
            .in2(_gnd_net_),
            .in3(N__15819),
            .lcout(\c0.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__1_LC_15_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__1_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__1_LC_15_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__1_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15877),
            .lcout(\c0.d_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19636),
            .ce(N__17176),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__1_LC_15_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__1_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__1_LC_15_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__1_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15853),
            .lcout(\c0.d_4_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19636),
            .ce(N__17176),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNISRG61_39_LC_15_19_5 .C_ON=1'b0;
    defparam \c0.d_4_RNISRG61_39_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNISRG61_39_LC_15_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNISRG61_39_LC_15_19_5  (
            .in0(N__16647),
            .in1(N__18876),
            .in2(N__17484),
            .in3(N__17745),
            .lcout(),
            .ltout(\c0.un1_data_in_6__2_0_a2_6_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIK7NH1_24_LC_15_19_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIK7NH1_24_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIK7NH1_24_LC_15_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIK7NH1_24_LC_15_19_6  (
            .in0(N__16434),
            .in1(N__16405),
            .in2(N__16384),
            .in3(N__18819),
            .lcout(\c0.un1_data_in_6__2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI5G09_46_LC_15_20_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI5G09_46_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI5G09_46_LC_15_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI5G09_46_LC_15_20_0  (
            .in0(N__17619),
            .in1(N__16367),
            .in2(N__18004),
            .in3(N__16335),
            .lcout(),
            .ltout(\c0.un1_data_in_7__2_0_a2_0_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI9IAQ1_14_LC_15_20_1 .C_ON=1'b0;
    defparam \c0.d_4_RNI9IAQ1_14_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI9IAQ1_14_LC_15_20_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.d_4_RNI9IAQ1_14_LC_15_20_1  (
            .in0(N__16306),
            .in1(_gnd_net_),
            .in2(N__16285),
            .in3(N__16222),
            .lcout(\c0.un1_data_in_7__2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIQ1PT_14_LC_15_20_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIQ1PT_14_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIQ1PT_14_LC_15_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIQ1PT_14_LC_15_20_2  (
            .in0(N__16273),
            .in1(N__16670),
            .in2(N__17791),
            .in3(N__16246),
            .lcout(\c0.un1_data_in_7__2_0_a2_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI9FFL_29_LC_15_20_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI9FFL_29_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI9FFL_29_LC_15_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNI9FFL_29_LC_15_20_3  (
            .in0(N__16213),
            .in1(N__16197),
            .in2(_gnd_net_),
            .in3(N__17620),
            .lcout(),
            .ltout(\c0.un1_data_in_7__3_0_a2_0_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI6GFI3_15_LC_15_20_4 .C_ON=1'b0;
    defparam \c0.d_4_RNI6GFI3_15_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI6GFI3_15_LC_15_20_4 .LUT_INIT=16'b0010100000010100;
    LogicCell40 \c0.d_4_RNI6GFI3_15_LC_15_20_4  (
            .in0(N__16162),
            .in1(N__16480),
            .in2(N__16141),
            .in3(N__16138),
            .lcout(\c0.m163_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__1_LC_15_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__1_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__1_LC_15_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__1_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16123),
            .lcout(\c0.d_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19644),
            .ce(N__17180),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI26S41_15_LC_15_20_7 .C_ON=1'b0;
    defparam \c0.d_4_RNI26S41_15_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI26S41_15_LC_15_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.d_4_RNI26S41_15_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(N__16532),
            .in2(_gnd_net_),
            .in3(N__16515),
            .lcout(\c0.N_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0_LC_15_21_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_0_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_0_LC_15_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.byte_transmit_counter2_0_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__18531),
            .in2(N__16474),
            .in3(N__16473),
            .lcout(\c0.byte_transmit_counter2Z0Z_0 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\c0.un1_byte_transmit_counter2_1_cry_0 ),
            .clk(N__19651),
            .ce(),
            .sr(N__19365));
    defparam \c0.byte_transmit_counter2_1_LC_15_21_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_1_LC_15_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_1_LC_15_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.byte_transmit_counter2_1_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__18764),
            .in2(_gnd_net_),
            .in3(N__16459),
            .lcout(\c0.byte_transmit_counter2Z0Z_1 ),
            .ltout(),
            .carryin(\c0.un1_byte_transmit_counter2_1_cry_0 ),
            .carryout(\c0.un1_byte_transmit_counter2_1_cry_1 ),
            .clk(N__19651),
            .ce(),
            .sr(N__19365));
    defparam \c0.byte_transmit_counter2_2_LC_15_21_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2_LC_15_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2_LC_15_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.byte_transmit_counter2_2_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__18708),
            .in2(_gnd_net_),
            .in3(N__16456),
            .lcout(\c0.byte_transmit_counter2Z0Z_2 ),
            .ltout(),
            .carryin(\c0.un1_byte_transmit_counter2_1_cry_1 ),
            .carryout(\c0.un1_byte_transmit_counter2_1_cry_2 ),
            .clk(N__19651),
            .ce(),
            .sr(N__19365));
    defparam \c0.byte_transmit_counter2_3_LC_15_21_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_3_LC_15_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_3_LC_15_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.byte_transmit_counter2_3_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__17863),
            .in2(_gnd_net_),
            .in3(N__16453),
            .lcout(\c0.byte_transmit_counter2Z0Z_3 ),
            .ltout(),
            .carryin(\c0.un1_byte_transmit_counter2_1_cry_2 ),
            .carryout(\c0.un1_byte_transmit_counter2_1_cry_3 ),
            .clk(N__19651),
            .ce(),
            .sr(N__19365));
    defparam \c0.byte_transmit_counter2_4_LC_15_21_4 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_4_LC_15_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_4_LC_15_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.byte_transmit_counter2_4_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__17824),
            .in2(_gnd_net_),
            .in3(N__16450),
            .lcout(\c0.byte_transmit_counter2Z0Z_4 ),
            .ltout(),
            .carryin(\c0.un1_byte_transmit_counter2_1_cry_3 ),
            .carryout(\c0.un1_byte_transmit_counter2_1_cry_4 ),
            .clk(N__19651),
            .ce(),
            .sr(N__19365));
    defparam \c0.byte_transmit_counter2_5_LC_15_21_5 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_5_LC_15_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_5_LC_15_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.byte_transmit_counter2_5_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__17839),
            .in2(_gnd_net_),
            .in3(N__16447),
            .lcout(\c0.byte_transmit_counter2Z0Z_5 ),
            .ltout(),
            .carryin(\c0.un1_byte_transmit_counter2_1_cry_4 ),
            .carryout(\c0.un1_byte_transmit_counter2_1_cry_5 ),
            .clk(N__19651),
            .ce(),
            .sr(N__19365));
    defparam \c0.byte_transmit_counter2_6_LC_15_21_6 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_6_LC_15_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_6_LC_15_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.byte_transmit_counter2_6_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__17851),
            .in2(_gnd_net_),
            .in3(N__16444),
            .lcout(\c0.byte_transmit_counter2Z0Z_6 ),
            .ltout(),
            .carryin(\c0.un1_byte_transmit_counter2_1_cry_5 ),
            .carryout(\c0.un1_byte_transmit_counter2_1_cry_6 ),
            .clk(N__19651),
            .ce(),
            .sr(N__19365));
    defparam \c0.byte_transmit_counter2_7_LC_15_21_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_7_LC_15_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_7_LC_15_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.byte_transmit_counter2_7_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__17875),
            .in2(_gnd_net_),
            .in3(N__16441),
            .lcout(\c0.byte_transmit_counter2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19651),
            .ce(),
            .sr(N__19365));
    defparam \c0.tx2_data_RNO_3_1_LC_15_22_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_1_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_1_LC_15_22_1 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \c0.tx2_data_RNO_3_1_LC_15_22_1  (
            .in0(N__16674),
            .in1(N__18526),
            .in2(N__18333),
            .in3(N__16651),
            .lcout(\c0.tx2_data_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_2_LC_15_22_2 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_2_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_2_LC_15_22_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_2_LC_15_22_2  (
            .in0(N__19818),
            .in1(N__17554),
            .in2(_gnd_net_),
            .in3(N__16624),
            .lcout(\c0.tx2.o_Tx_Serial_RNOZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_1_LC_15_22_3 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_1_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_1_LC_15_22_3 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \c0.tx2_data_RNO_1_1_LC_15_22_3  (
            .in0(N__18282),
            .in1(N__18527),
            .in2(N__16615),
            .in3(N__17311),
            .lcout(\c0.tx2_data_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_15_22_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_15_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_15_22_4  (
            .in0(N__16570),
            .in1(N__17103),
            .in2(_gnd_net_),
            .in3(N__18968),
            .lcout(\c0.tx2.r_Clock_Count_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_5_LC_15_22_5 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_5_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_5_LC_15_22_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_5_LC_15_22_5  (
            .in0(N__16588),
            .in1(N__18601),
            .in2(_gnd_net_),
            .in3(N__19817),
            .lcout(\c0.tx2.o_Tx_Serial_RNOZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_LC_15_22_7 .C_ON=1'b0;
    defparam \c0.tx2_transmit_LC_15_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_LC_15_22_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx2_transmit_LC_15_22_7  (
            .in0(N__19722),
            .in1(N__19353),
            .in2(_gnd_net_),
            .in3(N__16579),
            .lcout(\c0.tx2_transmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_LC_15_23_0 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_LC_15_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_0_c_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__16569),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\c0.tx2.r_Clock_Count12_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_15_23_1 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_15_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__16558),
            .in2(N__17112),
            .in3(N__19001),
            .lcout(\c0.tx2.r_Clock_Count_i_1 ),
            .ltout(),
            .carryin(\c0.tx2.r_Clock_Count12_cry_0 ),
            .carryout(\c0.tx2.r_Clock_Count12_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_15_23_2 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_15_23_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_15_23_2  (
            .in0(N__19019),
            .in1(N__16552),
            .in2(N__17114),
            .in3(_gnd_net_),
            .lcout(\c0.tx2.r_Clock_Count_i_2 ),
            .ltout(),
            .carryin(\c0.tx2.r_Clock_Count12_cry_1 ),
            .carryout(\c0.tx2.r_Clock_Count12_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_15_23_3 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_15_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__17125),
            .in2(N__17113),
            .in3(N__18983),
            .lcout(\c0.tx2.r_Clock_Count_i_3 ),
            .ltout(),
            .carryin(\c0.tx2.r_Clock_Count12_cry_2 ),
            .carryout(\c0.tx2.r_Clock_Count12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_15_23_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_15_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17119),
            .lcout(\c0.tx2.r_Clock_Count12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__5_LC_15_23_5 .C_ON=1'b0;
    defparam \c0.data_out_3__5_LC_15_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__5_LC_15_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_3__5_LC_15_23_5  (
            .in0(N__17093),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19666),
            .ce(),
            .sr(N__16876));
    defparam \c0.tx2.o_Tx_Serial_RNO_6_LC_15_24_0 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_6_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_6_LC_15_24_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_6_LC_15_24_0  (
            .in0(N__16732),
            .in1(N__16720),
            .in2(_gnd_net_),
            .in3(N__19811),
            .lcout(),
            .ltout(\c0.tx2.o_Tx_Serial_RNOZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_4_LC_15_24_1 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_4_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_4_LC_15_24_1 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_4_LC_15_24_1  (
            .in0(N__19741),
            .in1(N__19191),
            .in2(N__16708),
            .in3(N__16705),
            .lcout(),
            .ltout(\c0.tx2.m195_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_1_LC_15_24_2 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_1_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_1_LC_15_24_2 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_1_LC_15_24_2  (
            .in0(N__16696),
            .in1(N__19193),
            .in2(N__16690),
            .in3(N__16687),
            .lcout(),
            .ltout(\c0.tx2.N_196_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_0_LC_15_24_3 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_0_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_0_LC_15_24_3 .LUT_INIT=16'b0011000000110011;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_0_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__19048),
            .in2(N__16678),
            .in3(N__19138),
            .lcout(\c0.tx2.N_205_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNI7NQN_2_LC_15_24_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNI7NQN_2_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNI7NQN_2_LC_15_24_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \c0.tx2.r_SM_Main_RNI7NQN_2_LC_15_24_4  (
            .in0(N__19870),
            .in1(_gnd_net_),
            .in2(N__19141),
            .in3(_gnd_net_),
            .lcout(\c0.tx2.N_493 ),
            .ltout(\c0.tx2.N_493_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0_LC_15_24_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0_LC_15_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_0_LC_15_24_5 .LUT_INIT=16'b0000000010011100;
    LogicCell40 \c0.tx2.r_Bit_Index_0_LC_15_24_5  (
            .in0(N__19249),
            .in1(N__19192),
            .in2(N__17413),
            .in3(N__19764),
            .lcout(\c0.tx2.r_Bit_IndexZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19671),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_LC_15_24_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_LC_15_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_LC_15_24_6 .LUT_INIT=16'b1111110011011100;
    LogicCell40 \c0.tx2.r_Tx_Active_LC_15_24_6  (
            .in0(N__19078),
            .in1(N__19946),
            .in2(N__19720),
            .in3(N__19248),
            .lcout(\c0.tx2_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19671),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_LC_15_25_0 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_LC_15_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.tx2.o_Tx_Serial_LC_15_25_0 .LUT_INIT=16'b1110000011110001;
    LogicCell40 \c0.tx2.o_Tx_Serial_LC_15_25_0  (
            .in0(N__19222),
            .in1(N__19875),
            .in2(N__17391),
            .in3(N__17410),
            .lcout(PIN_3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19674),
            .ce(),
            .sr(N__19771));
    defparam \c0.data_in_frame_7__0_LC_16_17_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__0_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__0_LC_16_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__0_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17374),
            .lcout(\c0.data_in_frame_7_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19623),
            .ce(N__17171),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__1_LC_16_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__1_LC_16_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__1_LC_16_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__1_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17341),
            .lcout(\c0.data_in_frame_7_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19623),
            .ce(N__17171),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__5_LC_16_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__5_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__5_LC_16_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__5_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17292),
            .lcout(\c0.data_in_frame_6_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19623),
            .ce(N__17171),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__5_LC_16_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__5_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__5_LC_16_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__5_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17271),
            .lcout(\c0.data_in_frame_7_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19623),
            .ce(N__17171),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__6_LC_16_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__6_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__6_LC_16_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__6_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17247),
            .lcout(\c0.data_in_frame_7_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19623),
            .ce(N__17171),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__6_LC_16_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__6_LC_16_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__6_LC_16_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__6_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17217),
            .lcout(\c0.data_in_frame_6_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19623),
            .ce(N__17171),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__2_LC_16_18_4 .C_ON=1'b0;
    defparam \c0.data_in_6__2_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__2_LC_16_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__2_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17790),
            .lcout(\c0.data_in_6_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19637),
            .ce(N__17727),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_5_LC_16_19_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_5_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_5_LC_16_19_0 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx2_data_RNO_0_5_LC_16_19_0  (
            .in0(N__18567),
            .in1(N__17677),
            .in2(N__17656),
            .in3(N__18301),
            .lcout(\c0.tx2_data_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_5_LC_16_19_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_5_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_5_LC_16_19_1 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \c0.tx2_data_RNO_4_5_LC_16_19_1  (
            .in0(N__18569),
            .in1(N__17618),
            .in2(N__18352),
            .in3(N__17590),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_4Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_5_LC_16_19_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_5_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_5_LC_16_19_2 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \c0.tx2_data_RNO_2_5_LC_16_19_2  (
            .in0(N__18712),
            .in1(N__17881),
            .in2(N__17566),
            .in3(N__18791),
            .lcout(),
            .ltout(\c0.m75_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_5_LC_16_19_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_5_LC_16_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_5_LC_16_19_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \c0.tx2.r_Tx_Data_5_LC_16_19_3  (
            .in0(N__18713),
            .in1(N__17563),
            .in2(N__17557),
            .in3(N__17521),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19645),
            .ce(N__19969),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_5_LC_16_19_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_5_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_5_LC_16_19_5 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx2_data_RNO_1_5_LC_16_19_5  (
            .in0(N__18304),
            .in1(N__17542),
            .in2(N__17533),
            .in3(N__18568),
            .lcout(\c0.tx2_data_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_7_LC_16_19_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_7_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_7_LC_16_19_6 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx2_data_RNO_0_7_LC_16_19_6  (
            .in0(N__18565),
            .in1(N__17515),
            .in2(N__17485),
            .in3(N__18302),
            .lcout(\c0.tx2_data_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_0_LC_16_19_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_0_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_0_LC_16_19_7 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx2_data_RNO_1_0_LC_16_19_7  (
            .in0(N__18303),
            .in1(N__17440),
            .in2(N__17425),
            .in3(N__18566),
            .lcout(\c0.tx2_data_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_0_LC_16_20_0 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_0_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_0_LC_16_20_0 .LUT_INIT=16'b1110000011101111;
    LogicCell40 \c0.wait_for_transmission_RNO_0_LC_16_20_0  (
            .in0(N__17805),
            .in1(N__20012),
            .in2(N__19340),
            .in3(N__18141),
            .lcout(\c0.N_170_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_6_LC_16_20_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_6_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_6_LC_16_20_1 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx2_data_RNO_4_6_LC_16_20_1  (
            .in0(N__18519),
            .in1(N__18124),
            .in2(N__18106),
            .in3(N__18278),
            .lcout(\c0.tx2_data_RNO_4Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_4_LC_16_20_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_4_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_4_LC_16_20_2 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \c0.tx2_data_RNO_3_4_LC_16_20_2  (
            .in0(N__18513),
            .in1(N__18061),
            .in2(N__18331),
            .in3(N__18043),
            .lcout(\c0.tx2_data_RNO_3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_4_LC_16_20_4 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_4_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_4_LC_16_20_4 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \c0.tx2_data_RNO_4_4_LC_16_20_4  (
            .in0(N__18003),
            .in1(N__18518),
            .in2(N__18332),
            .in3(N__17968),
            .lcout(\c0.tx2_data_RNO_4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_5_LC_16_20_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_5_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_5_LC_16_20_5 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx2_data_RNO_3_5_LC_16_20_5  (
            .in0(N__18520),
            .in1(N__17929),
            .in2(N__17911),
            .in3(N__18274),
            .lcout(\c0.tx2_data_RNO_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNI8GE8_7_LC_16_21_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNI8GE8_7_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNI8GE8_7_LC_16_21_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \c0.byte_transmit_counter2_RNI8GE8_7_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__17874),
            .in2(_gnd_net_),
            .in3(N__17862),
            .lcout(),
            .ltout(\c0.m45_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNIK84L_4_LC_16_21_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNIK84L_4_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNIK84L_4_LC_16_21_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.byte_transmit_counter2_RNIK84L_4_LC_16_21_1  (
            .in0(N__17850),
            .in1(N__17838),
            .in2(N__17827),
            .in3(N__17823),
            .lcout(\c0.N_204_mux ),
            .ltout(\c0.N_204_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNIKKP11_1_LC_16_21_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNIKKP11_1_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNIKKP11_1_LC_16_21_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \c0.byte_transmit_counter2_RNIKKP11_1_LC_16_21_2  (
            .in0(N__18654),
            .in1(N__18762),
            .in2(N__17812),
            .in3(N__18482),
            .lcout(\c0.N_215_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_0_LC_16_21_3 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_0_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_0_LC_16_21_3 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \c0.tx2_data_RNO_3_0_LC_16_21_3  (
            .in0(N__18483),
            .in1(N__18901),
            .in2(N__18329),
            .in3(N__18883),
            .lcout(\c0.tx2_data_RNO_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_0_LC_16_21_4 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_0_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_0_LC_16_21_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx2_data_RNO_4_0_LC_16_21_4  (
            .in0(N__18532),
            .in1(N__18856),
            .in2(N__18829),
            .in3(N__18267),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_0_LC_16_21_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_0_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_0_LC_16_21_5 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \c0.tx2_data_RNO_2_0_LC_16_21_5  (
            .in0(N__18763),
            .in1(N__18730),
            .in2(N__18724),
            .in3(N__18655),
            .lcout(),
            .ltout(\c0.m146_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_0_LC_16_21_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_0_LC_16_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_0_LC_16_21_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx2.r_Tx_Data_0_LC_16_21_6  (
            .in0(N__18656),
            .in1(N__18613),
            .in2(N__18604),
            .in3(N__18157),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19659),
            .ce(N__19968),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_0_LC_16_21_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_0_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_0_LC_16_21_7 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \c0.tx2_data_RNO_0_0_LC_16_21_7  (
            .in0(N__18484),
            .in1(N__18406),
            .in2(N__18330),
            .in3(N__18181),
            .lcout(\c0.tx2_data_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_0_LC_16_22_0 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count_0_LC_16_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count_0_LC_16_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \c0.tx2.r_Clock_Count_0_LC_16_22_0  (
            .in0(N__18947),
            .in1(N__18970),
            .in2(N__18933),
            .in3(N__18934),
            .lcout(\c0.tx2.r_Clock_CountZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\c0.tx2.un1_r_Clock_Count_cry_0 ),
            .clk(N__19667),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_1_LC_16_22_1 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count_1_LC_16_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count_1_LC_16_22_1 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \c0.tx2.r_Clock_Count_1_LC_16_22_1  (
            .in0(N__18954),
            .in1(_gnd_net_),
            .in2(N__19006),
            .in3(N__18151),
            .lcout(\c0.tx2.r_Clock_CountZ0Z_1 ),
            .ltout(),
            .carryin(\c0.tx2.un1_r_Clock_Count_cry_0 ),
            .carryout(\c0.tx2.un1_r_Clock_Count_cry_1 ),
            .clk(N__19667),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_2_LC_16_22_2 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count_2_LC_16_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count_2_LC_16_22_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \c0.tx2.r_Clock_Count_2_LC_16_22_2  (
            .in0(N__18948),
            .in1(_gnd_net_),
            .in2(N__19024),
            .in3(N__18148),
            .lcout(\c0.tx2.r_Clock_CountZ0Z_2 ),
            .ltout(),
            .carryin(\c0.tx2.un1_r_Clock_Count_cry_1 ),
            .carryout(\c0.tx2.un1_r_Clock_Count_cry_2 ),
            .clk(N__19667),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_3_LC_16_22_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count_3_LC_16_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count_3_LC_16_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \c0.tx2.r_Clock_Count_3_LC_16_22_3  (
            .in0(N__18955),
            .in1(N__18987),
            .in2(_gnd_net_),
            .in3(N__18145),
            .lcout(\c0.tx2.r_Clock_CountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19667),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_RNIE5AU_3_LC_16_22_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count_RNIE5AU_3_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count_RNIE5AU_3_LC_16_22_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx2.r_Clock_Count_RNIE5AU_3_LC_16_22_6  (
            .in0(N__19020),
            .in1(N__19002),
            .in2(N__18988),
            .in3(N__18969),
            .lcout(\c0.tx2.N_171_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNI9USD1_4_LC_16_23_0 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNI9USD1_4_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNI9USD1_4_LC_16_23_0 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \c0.tx2.r_SM_Main_RNI9USD1_4_LC_16_23_0  (
            .in0(N__19246),
            .in1(N__19221),
            .in2(N__19912),
            .in3(N__19857),
            .lcout(\c0.tx2.N_16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNI9USD1_0_4_LC_16_23_1 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNI9USD1_0_4_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNI9USD1_0_4_LC_16_23_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.tx2.r_SM_Main_RNI9USD1_0_4_LC_16_23_1  (
            .in0(N__19856),
            .in1(N__19219),
            .in2(N__19915),
            .in3(N__19245),
            .lcout(\c0.tx2.r_Clock_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_0_LC_16_23_2 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_0_LC_16_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_0_LC_16_23_2 .LUT_INIT=16'b1111111100110010;
    LogicCell40 \c0.tx2.r_SM_Main_0_LC_16_23_2  (
            .in0(N__19220),
            .in1(N__19134),
            .in2(N__19258),
            .in3(N__19858),
            .lcout(\c0.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.N_90_ip_RNO_0_LC_16_23_3 .C_ON=1'b0;
    defparam \c0.tx2.N_90_ip_RNO_0_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.N_90_ip_RNO_0_LC_16_23_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.tx2.N_90_ip_RNO_0_LC_16_23_3  (
            .in0(N__19133),
            .in1(N__19164),
            .in2(_gnd_net_),
            .in3(N__19899),
            .lcout(),
            .ltout(\c0.tx2.N_83_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.N_90_ip_LC_16_23_4 .C_ON=1'b0;
    defparam \c0.tx2.N_90_ip_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.N_90_ip_LC_16_23_4 .LUT_INIT=16'b1001111011111111;
    LogicCell40 \c0.tx2.N_90_ip_LC_16_23_4  (
            .in0(N__19218),
            .in1(N__19045),
            .in2(N__18916),
            .in3(N__18907),
            .lcout(\c0.N_90_dup ),
            .ltout(\c0.N_90_dup_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNO_0_1_LC_16_23_5 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNO_0_1_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNO_0_1_LC_16_23_5 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \c0.tx2.r_SM_Main_RNO_0_1_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(N__19105),
            .in2(N__18913),
            .in3(N__19903),
            .lcout(),
            .ltout(\c0.tx2.i97_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_1_LC_16_23_6 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_1_LC_16_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_1_LC_16_23_6 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \c0.tx2.r_SM_Main_1_LC_16_23_6  (
            .in0(N__19166),
            .in1(N__19952),
            .in2(N__18910),
            .in3(_gnd_net_),
            .lcout(\c0.tx2.r_SM_Main_dup_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.N_90_ip_RNO_1_LC_16_23_7 .C_ON=1'b0;
    defparam \c0.tx2.N_90_ip_RNO_1_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.N_90_ip_RNO_1_LC_16_23_7 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \c0.tx2.N_90_ip_RNO_1_LC_16_23_7  (
            .in0(N__19132),
            .in1(N__19165),
            .in2(_gnd_net_),
            .in3(N__19898),
            .lcout(\c0.tx2.r_SM_Main_illegal_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNO_0_0_LC_16_24_0 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNO_0_0_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNO_0_0_LC_16_24_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.tx2.r_SM_Main_RNO_0_0_LC_16_24_0  (
            .in0(N__19047),
            .in1(N__20011),
            .in2(_gnd_net_),
            .in3(N__19167),
            .lcout(\c0.tx2.N_214_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_RNIPHKF1_0_LC_16_24_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_RNIPHKF1_0_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_RNIPHKF1_0_LC_16_24_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \c0.tx2.r_Bit_Index_RNIPHKF1_0_LC_16_24_1  (
            .in0(N__19861),
            .in1(N__19139),
            .in2(N__19198),
            .in3(N__19247),
            .lcout(\c0.tx2.N_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNI8OQN_3_LC_16_24_2 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNI8OQN_3_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNI8OQN_3_LC_16_24_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx2.r_SM_Main_RNI8OQN_3_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(N__19046),
            .in2(_gnd_net_),
            .in3(N__19859),
            .lcout(\c0.tx2.N_17_0 ),
            .ltout(\c0.tx2.N_17_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_4_LC_16_24_3 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_4_LC_16_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_4_LC_16_24_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.tx2.r_SM_Main_4_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19225),
            .in3(N__19106),
            .lcout(\c0.tx2.r_SM_Main_dup_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_RNIN3O01_1_LC_16_24_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_RNIN3O01_1_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_RNIN3O01_1_LC_16_24_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx2.r_Bit_Index_RNIN3O01_1_LC_16_24_4  (
            .in0(N__19747),
            .in1(N__19194),
            .in2(_gnd_net_),
            .in3(N__19815),
            .lcout(\c0.tx2.N_212_0 ),
            .ltout(\c0.tx2.N_212_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNO_0_2_LC_16_24_5 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNO_0_2_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNO_0_2_LC_16_24_5 .LUT_INIT=16'b0101010100000100;
    LogicCell40 \c0.tx2.r_SM_Main_RNO_0_2_LC_16_24_5  (
            .in0(N__19860),
            .in1(N__19140),
            .in2(N__19171),
            .in3(N__19168),
            .lcout(),
            .ltout(\c0.tx2.N_496_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_2_LC_16_24_6 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_2_LC_16_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_2_LC_16_24_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.tx2.r_SM_Main_2_LC_16_24_6  (
            .in0(N__19056),
            .in1(_gnd_net_),
            .in2(N__19144),
            .in3(N__19107),
            .lcout(\c0.tx2.r_SM_Main_dup_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_3_LC_16_24_7 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_3_LC_16_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_3_LC_16_24_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.tx2.r_SM_Main_3_LC_16_24_7  (
            .in0(N__19108),
            .in1(N__19077),
            .in2(N__19066),
            .in3(N__19057),
            .lcout(\c0.tx2.r_SM_Main_dup_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_RNILRI51_LC_16_25_0 .C_ON=1'b0;
    defparam \c0.tx2_transmit_RNILRI51_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_transmit_RNILRI51_LC_16_25_0 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \c0.tx2_transmit_RNILRI51_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(N__19913),
            .in2(N__19876),
            .in3(N__20014),
            .lcout(\c0.N_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNI5LQN_0_LC_16_25_1 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNI5LQN_0_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNI5LQN_0_LC_16_25_1 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \c0.tx2.r_SM_Main_RNI5LQN_0_LC_16_25_1  (
            .in0(N__19914),
            .in1(N__19871),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.tx2.N_9_1 ),
            .ltout(\c0.tx2.N_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_2_LC_16_25_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_2_LC_16_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_2_LC_16_25_2 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \c0.tx2.r_Bit_Index_2_LC_16_25_2  (
            .in0(N__19746),
            .in1(N__19780),
            .in2(N__19825),
            .in3(N__19816),
            .lcout(\c0.tx2.r_Bit_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_1_LC_16_25_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_1_LC_16_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_1_LC_16_25_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \c0.tx2.r_Bit_Index_1_LC_16_25_6  (
            .in0(N__19745),
            .in1(N__19779),
            .in2(_gnd_net_),
            .in3(N__19763),
            .lcout(\c0.tx2.r_Bit_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_LC_17_20_0 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_LC_17_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.wait_for_transmission_LC_17_20_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.wait_for_transmission_LC_17_20_0  (
            .in0(N__19723),
            .in1(N__19326),
            .in2(_gnd_net_),
            .in3(N__19684),
            .lcout(\c0.wait_for_transmissionZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19660),
            .ce(),
            .sr(N__19369));
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_18_16_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_18_16_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__19341),
            .in2(_gnd_net_),
            .in3(N__19291),
            .lcout(\c0.data_in_frame_0__0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
